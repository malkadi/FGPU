../../../../../VHDL_Files/V3/loc_indcs_generator.vhd