`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
gD7l84kB+WAh1ATog3H36h0/cMgn9QL5jGe9p9PjvP7N+FJAVvGVlrxcgBw6dZaWDNZqNANQuRFv
ZSE8fsSCFg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
YQUcxim/tlzHeVlJ7otHN7u41KO3Yg5DFb1yF4GCsbXGLtUvWNlkFjY+UPIlgYImR4Zo4dTHJQ+j
3BaUNSUOqAVzT9CfyUelv2YD2ZTfAtzIe1Mboyb3+StKnuzxnZmIhVPiZlowdW5lQ1r7BjDPOsge
ztxOfUTbvYcTUE1ABIE=

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
eu4MFD/NMz3pssr62VCh1XDd9mthYydX9VaOq3lWUwHi5/7e5dl2SAWHtYwTnBgGPY+jCcMycJhy
WSlkhQxVj5BsMm2aAItwXFvH2mSbjlPggtI0/+DNGQ4x8LQSFLTDYnnQbBrHlJymsS+/asMkXACD
SJ2tF8LF5tMhAlMPZZ0=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
rNAzbNlIFUMjdhvgzZ2FokzvR4AuFtV+1AHGDKa9QgeBsZ1e0Fom48uKbJ9iakvqUoUcKKAvRzeY
OBkbx9P7Imx0gvIgzFsgiVw23cBYWOhbhSqVb7mef9aKx8yeF8T48n7gKldUkwBHIPeqaayRI9/Q
HCZO+k2+HCjRZE6L/Gzd+IOdEVUFOg3NtWFPk2JFkfZkxs8X7Vg/xxtvH7uvp+/EbVyiMbnwDT/p
NSqOyA+rJwBJYD3xRIPTFDI83XJLCF+1i4E8hyu7Y0F9MtjKugqEHwAG+JK3jde00nzNNaeLVUQ1
OfFMZJpkk0Cg66d2cvJY/G11oPkmvTq/JZ4+5g==

`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
apuTRT8aJu0TR7Ciy6ONiGK4AT7TUEiokS4gFf1g+kDg6PdKk9VRun4HKszIadRtahjPQo0of9uS
yvu3GS4EQo+Y+T116wnAIXnZSa8EQaEsDkziOI+rCvXv8IgaPYN8Cq0aRlASFL7IHOWNI49V0c0A
FIG/+5U7ZyNQFCVwuE4gCgK/pA6apm5kY4FGJft/EdZ5YAbR/nCTzK4P53+XsKHrtGfw+/MthFWz
tI0OtloKqc7laKZWKOVFqWq8Qmq7UL6utFODtxEQqzczH+q+Gw4rkUyOosIY+cbB67hX+GlmXXEF
jMwvUcen9t6c+wiH6rmBDcUIiuUHHz6q+jCwJQ==

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
dfDj35aI8y6zqcW/IHFxmCDw2mpyex25qQAUnsL+tIRxivv/85PqpCOrf3b7NWnwUKMrsxtw+JBY
mtlPsVxQKR1gn6VkaHwbEgwxXXxFe71Z+1nWQhfF8Nt55jGvq1joWKMrurSV7Mo+HkvHMSszXj3v
8ElD0S6sN91oml0nObejOhxzHf0ybK+sGag+CFA7aBr4k4rYglf7AzOYrPl3nNoCkyrFDQFa46/w
SXJm/os7zUHbsDI5GGUH3BU+NktHZV6GK3iyhtHTwrMgDtpGk6vKHMKULM1Gjv9g1/jp9Ao4cUhr
bCVOXM1v2e8A3564rmh3if78zTzCKamPRAB5Ig==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5312)
`protect data_block
KwL5t2oQy0aWVwqsJj4aeW7VHmQ+JCGa+3Bi6mfEboVHQysd8CO8DGYaXDl7J0+3eDimAPPhh9BA
HpAnRupuvBy+QfB8Hw5xnnLG+ZUXuGPlIbrVQ6ot1EYyBLXzEHt5NjSLPUzDZsbptuISGCxiHGDB
uJnWeYkcfo8cdqO/WK1nsqTO1kpZ/h6RfdrKmhCyLBOpXkNUm/4k/YvTAPh9LI5otZgqaGtJt2l5
JUuJdF5XjtPSiY+IjWh7Ts5SEEaTrf6SRjnDhXOJu1aPOM4wNDSAiM9D9mwmyaELBXQsFWPM43H9
A7rzPza1SRt0Z3qyyZ5SD0TP3EJ5mmNo0/jK+b5PpmmzySFQE8B8JixIBXQQIss/9QcEK2dg9MBF
6MtxJup3ZRXuYLcftjSPVz8ccjpU68cnA+ZNXmk7yyoiNoBEh4MJ0jUpnTTyhBXDjaA9fTTFoGgb
lXlZGcpJZJA3CevRCUTz5/xm0VX4AcBVSohsAt60QDXv+9LVYv6Zi6V9w63mvVRLm+Q1KYTis6+S
2o59ijBMvyr9GsntcVnvcipKyyI9L5nc72HBNMZkGvPrlmL3URVjB05Z2X1GAhS5WTOab6elScCV
8FXXQm7zfdsU9OzYdShYaZ2/Frt6HJHF9Y3mo4/mhssj1BVFp7QH1VCjosytOBXUijaLxmFrJbB0
PYVpdz02+Bz4eCqbMR3snV6aAwsrgooMB4ow6I+9LiaC1WyKoLasb6JfL2ViZJrGa7Cay8AA5tup
N94bgGZnOZedq+y+ap7lzjUrd3sCTBBP01DFpLygUBm3KdtkaBbRJalGC9U+0gujGfdYxNfthn9f
JylnoWWI1hp7Aki7kmKDq7G8OPeZeTcqCaPJF2IXZ391eE8suq/qHJmoCUAOITN5JC7T82hB5qnY
tph++2VdvlQ2JNt7/HPFb4VjhMHVsESgBqgtJxFvh0gN/30QvmQWnzqyrZ4h/0ZbAf7pHi9AJbe0
qAZQmKcw8asxWuG9H8cGQi/dpVnslWDtCmIvXFgCE0pM7Kn2DNBR35APnoYgWyG7WC763a2d8NyZ
cC8e6NivQWPMvyd4C2qlC78NLEQLNXZJM2nDkgn/nnJzjvhMzgmBOeccIfmT5HLJmgcwlyAS9lJJ
DJMSNWUYRxusAvXPJ564n3Bu4WJhCg1/cF2eZaA92IZPF1YiA3ZL7KNGlh8AS0NGEQdGHCBPLjiL
9KTBVZysSPyPbPpUBOJaGfmvc4Sar66MU2Qv6F2cDiiHQz4HD+LKRaOUVliwcAMsr2PM5V8qmrOk
tx7VwSXwdOzkKze1rubnmGmfmMHdwTiv3zB8AYAGUae5+a1rvHeBplnC3UbeJRhEBtO8sr5XQL1N
KDhg/LWFDXv499kYGGw0A7iHkrDsyTjmM3FJLljK85oVFM420o6fU3npDUltgN7SdQvhzwpCU1jg
NFP/rB/X7Nps0pOFu702PCgVA3uIYvjigTpCEgtTq4/SKMJgn3znwS8VGJYDAbxa3miEz+xKrKLm
Aq/l6C3mpKpYK6TCcgLDbjsLC5tcwms6mjelc+C5UJyJf54QImFpk4+CefREdNBL9hx0WLuQ/xaA
nxGO1HXRocs/X2r2fg/H/r3y3LCSN4PJEc3yCSHUJbaEPRfngH35XGdWkv9tdGRaRxTwUb9OUYqP
LX2wTXhxrmKFfCv//D78qpjQvj3rGz9Of+Iefh7349hRfQ/bQFXNki6eBEmSngfmHdNlQDCIaRFk
oauUF2aFCem7ytjZ5azzFm9eRwpvoKvnn0WnGFC0SkDjZ3wSs3epmSnmEE8qcqf5H9e+ZpFpW6Xk
Or04CFO6Rp1njKao/FqPA3uH6+wS0ifamDKdZNLJiTbbPev0zekYJpwPIQUQYzASLpgtflT4gS8F
aOT5Wfh1URHsCJljhVKwwVWCCezRFDY/3s/ZkQcGwo2lWcLZvLjOqO9S1CXrt8N9blQeQF9h+D40
R/SBKBZWDGwuapA43qjwRC3cBA8JiOy75AG7mhi8yB75PltDRx7AoFGaU7LPLw2htfzMffWOSp/p
sjAW8GX/aK2ILB1j50PHS/FgeCbiqIgK1fLyP4L2hL0wZbtt9eeG3G0Bng9ZzaQMilOR4nHsNydq
wetKvqG8Ej+YaXT7xKpdYzPr/YzgB9iQ7ha+j7Pjqa3YoPIfyR3lKOVKbKIlrLBvaBSBe/7GKuRT
xVlWclUXwZtQwu127ZbvAKuAaLy9ZMhyENcUVrr2vndTDcx85W51RJ4/Id6wI+QuB/c11mAPwO3n
LXDE6MoNDlNxri27cDt7jhV0c2pv/zbhh7Xuh3t2pMHpWFmPv58jhFGz/gMzdSHHEw9jaQgy9kSH
xoVcOXan2co0GVmxl4uyAjoDHksf99lMGfMDWuLn32NiO9MxO5Y3QmB5it/sGQAC+CjQ22cRbxSA
+iEuAuBsQNB5oZGhM3keHpqbZohAzc1TAA7lQENDpuOhOG3kkimitlCtlNOXwDC85YTvh42lPeIe
dhEVE9Hl7coa+6U0H1U/6FO1gQKGwldSRv+GJjyis0RTFymi8ScuhF4uX1hA7AwONgWAbI857S3R
tUX+iNqkEM9/Guh4fwNCtiVoiJT1TQ9UiHJDBS3aMPZOEtL3Dr+XYTbIvnJDfSKyueJYaXB5x0sA
OyZ/35sbUJjULKzhTJAZN6cAN2XeV6/OhAO8LyF46yfdAWuLSTEfM1Jm+WzvQ54Y2VfYm7+KYa27
+wSbU3H62xoZtPcnShePYFWkdJIiE9amlj4szXbVwkOr0jk5WiniyFRn3/3YULASrIZqWz0uQvCk
66jxv+V0FMiJl+S/B4q9HiqAhMwLmoDPsUx6nm9O4ZNTYFR9Rwlj7n3Rrnj5vaRt9/kvqCeC38s6
XxQ/Q3Lb2f9+fQuKtVNQlzp9QXJilG1lcaZk0faCNPMAkLLr/pcwcN1NSovJrzVLVsR0Hit3Beyh
l3d+GRLvmTTu6dHVAWf+GS8JCSXncVgDGaK7e9QONI9yGKLhISZ5caVL/nLm2usPM+6GUfm3cUIc
WFdxfdXACMItZfC/P3HoMyD/hVmbn1zzwxd2dqL/Q75CQ5DBUIqXdSeOJiI5JdILkrDsKzZfAGg7
lccuF8M/7c0t9C18pB8Emtqg5foLLWVMXmZz/t1Wq3/G9Af/bNHIdqBZz3boV2Tj9oYIKj9DYZUV
sJr+UWVYyEv/LKR8JxDK4E6Uvwz+24VEQgGRRXHZQeGvJGgkcirz98UPzxbfufLV87GdPtlRJh3b
xfx08+fTJh4nN4HJ8N+HSfwhn1jSyq6yJOGEEk2qEZa+i5RxYkFivMy74qu7bmAV3NmZFlrQayHJ
LBMGEpwBHCjrZH5zOG0tywSE96KQ4ay0kyPdsHBYIW+MOwC+cpwZjvdOvHFqaTdoe342OrcDpq4F
WM/v7zOmrBaYpgxkLcSU2I0IVWxWkvPe8+6lmHfpww861kaWkIv2ndg0lf+ulWYTXLcPPMaqvoGW
2JPeiPIj4bJ6BWJam5hfMILEHJEHS2BD0HJS8mPGX6fxEDwXglVCQtvoPt6rtQFnd3YAlDiaLTBQ
PKfKINmW+j4SB5PfPzfAF7g9WXcEkw0/53kEzUqS+xECDBoKDP3EvttVoFX8Zbqlf2UsNj00x/Vt
0yz94KRvn2Jb8m89QZcVw0I2tVjgwg5p51bjdv+p8PUpuCappVck4X6SzjoiQ/4oaweHTotCBABS
TPyramJBVhSdS5co60MQG/tT6JUpALjqCO9rTfCBZmPkP3NlkziHiiAVtRV4Knb57+DBFe0H7iSV
BtbPoikuc02fUYzz+hTR0IgpgGMrxmwM4YeQzeoHKAdvxgIVYZumgxQmCPSUl9eJ+H+zQtwp0mlG
07lt4v8v/g5en+qzwSp2xRnM2JraUJRtfz4AzHCGLNQExpO83JYCraZ2s7QfbnCQCobIHnHOCHKd
0Y4DsNn/9UodrbNf8wq1Wx0s46ALDJhW58J8yQs4briVC4tTo0pJzvcP+L2hMA9F2oqLPoxLsnR6
BxYnUJyoCTzIULSwIWjc254PVGCYraJo/RdpVMv0ST/UC2410VT3SkRKNLd/txTGh1pTnptXwFXA
yTFjU1JUlNNe2MAsGDHGZuuB4qrik+yz6q77HMjZd7mBjKOK8fyxnOodPoNg/mNXHqbkStG5mczC
LPmt7r1PhPH9VMBlVysZprpNxWNinoPe99KDkZlQxNunHn4P7THmLbhy55Yx1iO4RKXxzhuYjEDT
n6SODVISDOBjG9aLoMXMFuuDSAuCoQRu7N7ITeJcyCdfGOBRgGdQRtEQ0BlUlqYFYJ8pnNSApTvA
RLRgYndO8uTiJnwBq6+Mga5tXkssJjaf19ihFuK9xzUwvf33YaZZpVSW5AdjOohwBNSX2qlLjSYi
DubnrcCH/nlgN/eBDtCX9lsHj4OSqPDqS3FACi7kFm9s4Sv2zCFgnsMzfF4P+2uOgF1cu4iRkUB2
byrVfCNCLZy6UPDyehJEZ7UobhJvIwO8BBzgTLTmAjkR1Dtdruc+E2hDS2KRB9PPId7et4ahH8/k
THtBrtTqU11qB+h6EVi+oTVzQxtABlIkDLWZmjdSrYkdbQvhg11VSooRCpeR4DlAE4od3ciVgLFo
dQw+jmlbYcHNtX99HFTdk1xykmx1nUqHRJBLkKB64z+k2X+E1glMlth9LuwxnlXcuXTBOXW5fLR9
wdf+PnnurroXGzrOL+oB0PB71qqkb4Tnp3lEoTArXNpAYM4oxrVD6ZFVxDTtdg9A6m8Tch7R6qfR
VMYYqlaI06RQOZrI9vBDdraKRRjatLWbFZzGVmlzRAs9LwbZR0Ha71U20cZoFmBmc8apDdmFEF/J
IGHmPgV8WkpAOb+BJrpygun+70hzkcAORqprb5+Kse7SMI0YtVSCRSHLqw2jEw5xIpqrsCNs9BSH
ZOt/jpp4XRwcIKxwg+xuMdiRXNxkxXpJY5LMoQXmykfKC1cmA26EqlvDazAO+NsedgawnLsE7XKL
0EE7X/De8Px22DGucCrAHh6b+dOcCeHEB7t1ZliP4wgnRPx8s6H9VdUnPFzg4XxeFMVLSwOFhV/m
btNaCyP4got5FGEl2qZ8WbKgA3DgrczyPVGlq/1S7lqYXHUSxPPSGrfiHBwlt9O3BiYFJLeSuxHF
tPMMP3Do55zw0IQRGRzfsLAG6+NFgbXNFlpBwQ1Eih5sIb4gm1AzHXwOzj7Xg93O9CpSuwYYat/G
kedviA6u7nsapX62suBvVKpZF5OtfeG+6r7VmfUJWdiCqvBgPwzHAhS+zaAogT/n7KlQbQ0Vb9yW
Gx2lAFvWdQ3FIi1jYPKSMQhb9bON8lWxpNhuxv3gm0hAdDpTj1T/eHWqejLChgXUMOiCY8Fh8/rM
znoyF2psvt4zZZm2Iy0vJfRneHHKwT12PvscYZ8MgK2WeHZXMYRcQxOhDE2VSZoMPuIsrPldCNSf
/q6jKOiidRYiZPq9VyHol9+8hbB8XilvCydI4ATPKGjxbsSasNXM3vupYjcYWFYl7NtJZ0Pol0e5
WsvCFFRm4sEzaOXvVlRux+YCXQT+VtsCuQ+0uDJEBiBbIMV86HfswJ4H/cAXrqM9RMtPhplvBfJ3
dqOqPf9THf68721atAdYzswgxOaRzjtFjRML4+g70XjwD/CVVNC2yK3NikofKDygWtDLZfkby01k
0YkwcPzmdYWCc5D7fGlNeVitj+jUyHWIw/YJ0mD6fKiKeuVDTOlQLx5MllXO9ZGXOLtBop/6kUdd
ZWXAPgX/KqFs6yDywZRoTTcwJkS7HqKoS8SqpAkg6Cr+cp0hbvw6s+p6zq5QkU/PHHPRvzXX3hIH
RvSsUG/PxOsPm5c6vfvlFJyOV/9Wsh3O5hEZ8t6DX6K61xcAXp/KwlEzt/zBELLc4KbeIz/QrU/3
Ha+r9YER7pp9Uas9oo4ECVutgHvURREdGeesxHgfCMEfU4J9aD3CyKkOifCfN+yF4veFqKiwG4kS
/2T2z6wCSdktCf9WXs4dINL8WK/ysQHc81UrPcLIwA79QDh0FK4kcU0XEGTSqU2Aqr4pKRcMJhsW
FftNlqEANvnrqXj7YJODjaH4E7q3ap3K5GutL23b6Wy9KM5WpqW6g/18uO6RqUhaYztfbJbY1mm4
K064VinuSlbPxsZ1wxEkW6IZ4MA3i4PagO1wxil9MeZ5hBDbprxSNEDXFNKoQYWVMus8CNNp4v8b
98059loOQIcqs7EPai01MhhKgY8LgmrDKHym3Bim4LCEVFWZoO1Cyowd2aJnT3hSkhAcIZ9DfBbn
j7RG92Yz0GoKsWt7YLdcODlLvRoLgU4DzUNdhukQdcDLToagcQIYczmuNiwRK+wnMrOqNB6s9NNJ
EJv0EW8wgm1c5RkW/KbsCV+TqhkMcEZQr9LBDe8u7nHTvIHJk8WNJndiva8DnV5uWZufLSn8O6M8
hCULhHv2tQZOmxw3w7Qmk6UtDUxmUSGB3CSXQMNBO1F5Pet/ihB2P0z9Jdlfef+9iw9U0AmuO+hQ
WwSXFLKb6ZCHn39QXTxBlWiyFn8TMZpTEv0cYEz/00loYrRTcU2sLFBOcBeAtt8Fj4exKXARXlRx
gDogLRNeEsT0ED+VB9Hly/LV+rKLcmKj4lkmjjy9q7tJ0xY6Tx1pZl5pvScqJydukEbPb0xo1nr4
WL07p93xNfRrK43CK3n5Ly7TEmmEBVCyE2MRnQAwc9mUynGTuF8NH9h3qEixFH2QFCcWEVq7qCUO
EEICTu5bNO+RWMIBnQvBfAs3f3BqTuwzp8nWxODJ6GI2yAqqQxSzGYHndfnls1cqbY2zZuybyLPq
IB7NQG7saz0MgL7Pw7Vfb/ilUkpwN0nE78rlqxuzPXqo2N0IhedHi8jeQ0avDR5+TuXPvqyXNqVg
S9iIZrCJddAETuw/7LK77bwhdZt/MiGtX/MEawamCRmT12kn+wMS9PI7yOAKe3i1gaYPNHscJ1cG
X5/w1p5pax8qREhRyAiTF+L7k4N4GtmRDwfJmflGnCkHAgt8ClAA7mHXMaWDZR1CAyG3yq1wTwkY
80v5tusTwzDChc0=
`protect end_protected
