../../../../../VHDL_Files/V3/mult_add_sub.vhd