`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
VbV3K+no6bnPIa+zTPjJm+Za4h+e+mAdgfsol9fh12i5ry1s/9jFxbKNRkpLXaPaKwPx6tUXx2dM
rz7eLZ9g0Q==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
kTHC1aaUWUk/RMP8ryE9Otenia3ejjUZ515o8MyC5LPe9Q9HU4j6bokGKsgb9UOn6jCH1yruRDSs
b5lYfhLsxwdG5/eDjBvnNCSnM0RpZJbFrI7JmsFggBcbNUey9IsoQpsnxotoGgl++yh2M6dZZxeh
M1HjDezNtQIQF/ZYUx8=

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
snOGGdaAqd0xCCnl9qpy1A393jt9hiIkPmkASlieApKF1LOzirx0ZtNLBlVn/2B/+8mCYjHiacYR
yXR79FQlFUsb7jR6ke5jpzqLDYHrXjsSYlP6XweX9Iba7CTKn3lrruzWWFzPkW4aciBjkat8zMl+
9yQhqwSY0mgGYoE6xIU=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
VQtZeHq0wwSVd11a6wGUrcsL8nkp++GpoEJBF7q/cJp1a5TPQvxpDAKpIvxahkyYavXQtD2H32nS
gwb37S5yvNwWpKhcI75qsKCgrHwPz0e58zT8OT1nTnN4wbF1FEBlXqVhaSTCc+ruoYfFgLOvq8Vv
3UIMxyu4DNPhA3cgj0i5I/Qu4n9bb5ARKmILDDDRdJH79iOGyfSi4jSRGCnPG4R2jh+afwgHnGWt
mNPbEs6smG2ApIULJcWURoCv+u4G6+NuD3qACnBJrJOsa24eMAMLstL4ATkGasikUUNzIj2pEJk9
8hRULYLSgD4dit5Jx+Lh3eUe3LnJ8JB9XVtoZw==

`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
aCN2iFOrSMMrFBC1bx0+qYoAW1mWivPbraxjFsh9goPWGNSJROEmbdaUCrQw+sK5IYVwzj76ptqV
hsAbNcAaqw5xKu9/s0kIvO/tlRqx54JykJuHqpzdnuBilOYKpjmnbgm9GNfp/+2BtOw2C5F+WfKd
t/aWE78rilJxgDDpFvROYhHeArroRiPDpH4FEpMDsabE/eDN1VYxJ197aihMGaAb8fIZX+lksOX8
SFmUPSICS6CVQ6P8licCLIY/CEHAngVTpNVAiFE+py2fimPTacxjGEoMWvWoZ1i6T6AQTrYMMz+R
1X4TRxNWtAN+GlPoa5SiOGwGxNi7ipB7xDxwaw==

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qrTdR5jHfRKLAYgifBWWG6p4Z4xOoCaPlTZeSph/qlRBY+GOLFZqse0DC500mzihUvVh9uqSL0sf
QqIVIKXtc/vmkLTVkrTjVWF//xVSppNyDBiDklq4+hMBQ1FTa5kt+FmZnTAwglWAnFB9je3STA7g
1vEddZZb+4GvMNQLT8fmcEvlxiOCwHGS3w1CmsJDrgnj3mXpIWYgCYJussuOzZYHKflNfTUDZBPe
cnCqgDCFeSfQaV9rV08HR3U+NRSxKPM+ou7WhrHfBIPk4L59Sk5mI6TtkBzh+VX6GcvtZsnUqyUJ
yQju1UjuKFN4rX8QdS8sgdKQohC4pjYIVuoz0A==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 214080)
`protect data_block
nT6bncpOc6t34NIB5RhqMnLjJwmbqEsAwzjZuT0pnSR+SnFrbSaqKu/8i6SJK4qKpb+2nfcZmLqe
1R1vVcKVToo9pEvRyOVQLsZYDH1bIHTLco/zyaLmjBkP6iqoZ0eqUAl3t+9NRa7AF/ueuzrs7FLP
zq233fGdmagypUYylvN9Btg776mYB7x4A7iq4dkY+aap23s542HxL6JaIO1jq/2ffL3pSfX1Zs4N
F2Rz0e8FpCLIwB0IkEuFFZ7zaSx53NeeVFnjyOdVdOQpJ30fU//Mi6e8pB6YTNN3qJF/T/P05poQ
Cls2BWMKzSeTomB34tFBE/INwmH5DCDzidXH257zPEUIrRGznuqRpJPIH9q+fbVGsc5LNYnHqwBD
55JL55hpBg0vK0dDpmOZxDu81nHBgpVCIz62znBD/o0HQ5MuFORqWYGXa0BHUnzwSlfoq4L8TVCV
WLd8OEoB5gv4UEvnlmHNaKKRamfXmCWdx2WRrN9UcXBEFJ2FFVUU/lD4G4vbGgAwVO20pu3T5BVe
/mM6LobR/KJvadZ3wQjCGk+IgFJkOAiUgm1lHEr3is+7I9ZYD4p0JAFU1L/XW9Kq0K0NgK+khPJf
lwvdE3QvVDVJRrha/+yw6y6GK7zCmCj4TfyV//eZWkopSh1WOi507Pp9E7PC12t/Y9y2d3ZSs8o7
Dx9BGcNyuq7pReATrwi6oVPzeSHiwAn0y1Ih5JkWSpOfH+J4kONtx/5DRDbjsI6nicsqdQiwoiKj
nWp75CHupOT0obwIho7k2FFZM9yH/eUGhE104IzMHxZ0202rCh+s9cjZbnp7puPyi3WWlrXX/Hhl
KP3H/mAyHDmUas+fxuREID/sNniF3fcY4B2Crlf5rpZzRg8cCrWwaf1zUsTtBiQZL2Q3I0jxzk3I
5BW0W88LvwTMWi71/XQQVCxH+i+wFQqUYtIUBSd+GgTHFkXVufr945bOUWgxQy2j6E8VfGEYm8Gz
QQJQgGLoBHh6F/SsODJRF5YTnO4hk7dxh6cDChPxcuVAM6NZfi2tIXgLn3Oceu3SIX3Qe7HDFVQz
xMjmuLTHnOfs8TdcIY9nlMJgDFwzvsGnAtGWkVolaqVdFHaNPTLwkk2dhZ9qQvw0NZreN+XDl8Zo
bqBJzCt1A51DoTK4WDQQYUyTWY7RcIqSPgGcHwFXKMNHHjKpf32o7DTvuE7cVlQGJ6hgOS/Q0w2P
8ns1qmCMO/xYjnUSJOj0oKQWCYmJb1ZkE+hjl6I02SfHfTB+WKb3XjPeA14q3+irscrCDF4j7XDm
8c6HWV0m629qa5xT3ERnYoo2/RbesvoMgcE7uL5ODsyEvDa1GqkM27WHdCG2FcogQnb081kT4oqt
l6C1mRgKlZlWZmStQolb7BAjXPyBHArsEbGgbSk9ipt+J22BMvPrB90OGcHaPv/2eP8CCfalG3wL
YDatS/aujfOTfG7ehgFzZWcS8GFcCP+gfcZ9mcIkO2x48/4qpVAVxKvLH79xq5+sZK/IH3CgyVBI
cp3q/BomOzkk339suWcaXtdinYhnj1atoFntA+4lz8NjpyLNX9PrAOCPAsVW7pg1Zrzoj76ESAZg
2RHmPGaPcyEXYd8cx94WMiAo09kyonqjDlR7+pZ6XXrj4ywjKmccz3l2htasS11ebOWadxSZhaoi
Vb869rR63i9kdru3FVv9dpJAQIA1tf1/UyWB4GV2GIhO8JYQHhCzgf22Egp6QATrl4hLAL05OtZd
Qp5m3jlwKUKQ29++yr407aNxTRSyV0bG5IdKCJbpd/EFBkN/fSiUYXPeu/A3lN9cglkylQcyBjOy
hTTYCdwpAdot7D7KJ2a/e2Dlm9FInNJ5b/Ggu3WWTFxCHL2Cugzm7/R4F5X1aUXANpRmmTcCvUwe
QUTZkbOlNGlSB1wj2J4wlx2sf8fWXom+an9iwZ3OsR4PCnxNHb9V6Nyfx7TWBwNV9nMt4d92oEjn
N91q20y9vC6BpEmQZW+jd97j9VILuNBksLK6zu6fAGI8mFQG/xVJE/Wb0H2OCxclqsi9rnH7d4/o
J7IgYVRutyUZ8eRWpIkyEF6iHcp7n/S1HOG6aJMhNCLMzhdmxzFxLOJ5xv/aDoxxyLIACvARsF+H
WzHBBtnvlvPCH9ER50PTs4vmudzmIDDPUwH3EDQT/szu8nbmOxXqpSb5P62G524G9n8A+NDrAr6t
EOVCsdmXAGkS+2JBx5nP4HxTR3dyYz9nlFaivFva9ZGSiOhJZsZYPliyg9xshBBXVOlxxQ5hSwBy
GMz+3NqCcjq6YPoNI1OIAi3LGnXTURCOyeubNk38fMVDHsqvuFULi2wIMW59EqolcNjZht0mh+GX
qOGO3m98IroveNKTYy7tmYKFeyDQdDyow1Zc0O7I0Me5DESkUwSBaK+Sz3I9NGcnYJaQC+k0Ybve
63avOg4dJMpnNp0Kw/A5BW++4PbZzQ5Tg3VDjkDx4IaPoi41jcLR6jek1HcCQgsvzJ99Xup+3vp7
DZ/NViEdEzwAL1RtJp0YM0ZhWb0EU115+AzPjnsiqVoC8LI942QThRKGPCzDh7NeJlLUsFUvFlwW
cP0RpaNb+9O5eIoroVHyWXuHKueD/EhMCzFrt7HXG+yBlCkZ0CLC0VZPgWQ5vOuhsIMg2OkNAgBc
u07pz1pmcvihXCDdBIiXQ/iDsMwD7jNM6RX7BMo/SjxQXC9GWKS3/S1lT+GBE/hVpiXyVLDgU5qk
SJqnja2KM1XcY4cGHlXXpyJkhmzwQLvPKoeQZTV7eB4bQBmf4MQKWqT2nt1RPHkOv0BAWpirOWlj
Y1k6oGURrOSwNzlVxn4C8TcWgY8d+X4jEVKlZSoZNqgkOJMBEsMpUIhshALV2a2+GGxjN3GQql/j
IeIZ31usNJokhevOWZLnxUO2GLm4w3dqNGcNOf8NENOUVswVg9NoGpqM1bq6eRg14O6JrTKtTpz1
a3seI/KYRU2RTIaKx5IwnYj4UBq0oM+YBfY+EGz+wGjXBOUjqYY4Mjkjy1h6t1vix/mNE9/YrXp1
SUnJbiGjcT8P+4EfbeS0/bKUXyVJ0AB99iZj7rIAMfhdJnGguJNBtTJqJxJnz9CAtUiDpohNiPUM
rseEFhObJYiQzEc8Y2+KLvhnEbfds2HMb96+yEB9sDnWvpzUgPcWpjqK8zzf9dWJext32GkmAiMD
1uaT7CijaCb8hdCnffHPyEK4XIxUnux3SC4KlHWjOuxLeGZk7zddMwcEVJbzCBQpw0zvKzWl6B9N
QUd2te4MAezzcW8lci/ykD6F9SjbIu7g+oMdS0dXHv2OfjeMPJviCJ0trQ/eOLOtsSX2mHHlWoLk
vHjRuf8tKFHfqHUFbaAhnczcwFCHt8h70autzrHpnZxisVOhqEhdD6tZqRMeKX+wTsZo/0Dvqi9S
9frCReYR6C1S9lotd+BLtQiCnYjReGNMJ6H2fj8vnkIyOOm0MtSLo+esKkVL1VXo2cfqdr87P3Pb
/whjKvb9OGEqPMpdtqhbN5ehIGZTvBscNeZNAMUAx4pS/azStbmJT3aLBWtFGeywLQitBf7ZQdqG
+sJqf92/rD3Y3AoAxM8DlCol9rc/A7m/IloB5eW0FBP1z3lwWqueJw8J/Fzvj94TyVYKYVSBnVke
1lXZx8M/TPL/SRkXwFfGFZAGbGTkZEORmbUsoe63SDKle6bJYBXMZE1dDaBfw5Eu3F5wEBx4flX4
R7FNb6Md/84Qy7zDrfCpUhSYugcNGM5/W3/Cf+MKENQT7hUKwzlGr216DFM10+ATIz5mPNnIcWUZ
ieHpWB1ZKOTsh6SfCWMVhB3aGDNwKnaTC672IdfqMRcA0iQyAExTj0/MsRT5qOs5LayPtXd3izru
BpklBQn62gwUFSmNXh9QrQAWgJQTcItN1iOcJ3ZnpwKxKwUUOa17AD2liuXQLoBmIfSW2KOxz5sU
uAXPGIr/qD26o4Cyk/RLiyqhMKE8Tm9iAq8cqT5oK5eDHbG7QvRtf5MDdF3Q0KEnQaWD50xhVIOB
0OIErI5qQVkxiRUsnUz2SbwV+uDlVAZB5nwa3YqIOuG/NgGJieJVnibPE7Eo5EtoLwrfJjV6hGI/
KNKk8j7yqv6rKFsNNn6peK9hiX/pEthe0kHQ9TKgkSZ6xheqkTSINhjvzCrBAZANUtNR3vlN/Knq
W7ORtYpYMQp080RlrcqFOjJXFjVUeBHybgsDpdLwdf0RKcZVmvhuSt1zec8sL8Oa/jRFzvrkMaf1
PT/Hs5r9F4Q65J7aXK4YyZaIAqIXqwECEm13bPGKfxUNacfRxrkqWmqxI1+TqdKpb9DdxD6R0mXO
qozjpW1jMDFiW/Qfsrmp+oTnrWZnivDHv5axSs+9jfqgEuof5Zzr/iPk1QurPZPMeeRYxpSrtQHE
IOXJdaQknazhjVKKuZj8FZLqT5hu9PAMYQjz5AVpZUePa84wbcej5dld5s8pWBNM2rMh5uQGzYps
UOLLNQ48tbqyBhVz7hrDUpKAoia6y5sVV/+ovkaJQnCO7esW9r22dfMg3oApLU+HRwiip0F9Hdad
eovtIoQkZvDAgbsnsur68V823BFFbw4kVjTMBXdkVcFukM5jyaX3dluy3XiT7eAQ/ZaLUSARxoaR
gKsxHkMd4HBryL2ynR3/Gv3ICrRmEc+WobdXN7oXt3qUxXZHv0XkKR6W7rE+e8XUjcqIOxiSXcfz
KKtWd+HA/GeW3TNbZmKzr/FkTNpXAHSC8KqppcYs3IWB66R54bse+H38E7mFMtYC/OMOzgqYnjiq
w4FIi+d9QmOhTO1OK9VSB5vwNsDZLEZCARVMwjhmZI7gPGkCOSpdPNT+QTj3LUKPJeXtDPifCD9l
ufbMu29dlUwwmGwGJvXKRt+5zRu4PRwpwarT+RkV9CuqZO7fiIa4P5PDP16lJyTM2VKfN+RvlWd5
+QV/ZPsrK7anKsxPhdM9whDnhysCjUKkfY4NF752IyXWyTwASl+sB+iAUv2l/rtH9zkzi2uc3Kdw
hn3OFbenyi+FNLP5Dstwg5AaDlMWGrAzhHOTcCG8Q0ZEeqKkELYVzUmm7UjQPYAXi/vrZQIzPLX3
kPVpCbFBotZLbHMfXhwBd7YVIW6a9fgpIHQnDD5qJi852yG3AhIT3QHLHztPr7ZPvgy9hWmQ5hfO
OlPbrIr00MXyL+4eIZJyRpg8doNblOWaw5YioCdlO3U+0EYaZ4+GwrNsgz/TKY8X2UaArtYgHxn/
illgH3i8LBLf2r0BHFqEp7ZLDflqoCT4RdBRZS0uxHspiUOKR1xEpXMRavmNBoE23uGwPXnxyej3
rGjDLJXEb0+Ujmya4+WMUnTeS/7CapolFLB9KRyK5VCI7mBrEbqqIk5/AVq5A8GqyuirDQro+VIw
egtqazTsQhZ53k1AdOxZpJWUtPWbxDuSEBKOvIMk83ygKjFif+Xy4103Lw826nT9GwizZv5NEjj9
ME8VXj869bdjJg2ZCAe+Rjto+B2hRAmDInKsQW9EiyDsUEfTBvxETTC4Y4MX+9FYj3FNgnks6jMe
e6P6QhTkHyo6eNKxEIIEGe8Zp3LmhQ438azKT+3WjLGgTfq0cM1I0vHkFmeBQO3JhqCNLjJlgSPH
PleafaU5vwiQ+w/w3eKytl/rY6qC8UqkYW871hNPDWp7YKOL424xQ/YbdruvPWpf27MAhwaGztIC
72j9IaGzqw56BQtwysspkwBAhGhok790s/lMpFssoCdCfIEzfNEMMHe9XXHSEUsOXH/mw6xy8N5n
ipDYqtRfOFOkjVQ0rsLVk1yrnVkNJG403i6kMXeLAAK8Fef67Mbh0EtWnfei5NlYiPf+IRR5cx7l
DlcmC8cLG53WP93A+oyzInulA9X9hY3y8CKWAC3BalF5fHY7mafBxXDREgTSphDBsHoVL1qQND38
24uft/IJTbPspafYwdQ97VzoLq7FoYmy7usXjUU2mj3QS4KPOxIGm0DaYyzP5Rp5o7XYnGZl1gax
f2iNwFKqGGcmrX1P7NYMdENvOqxxtscUPckzQwzx36WTdYS0ol/1vB2pcGncjpRHptYD33Yva2f8
TrHejVPzjrYwbX1Dp3GD6AhTr64UErId6DI0Js87WacMUNL2VLfnu3Z8n5P86WTLpcFX+zLN+X7r
BFGoygd9QYvcWP/TQrTXSGafAUz/EOPmDPpcNe/Jimak7cTbhTy3P19wkFBeL2n/MsT31kkxs3rA
Sso0naj02UAy+cIxwYTqFS0jRoq4lbL6XBWuTOxSBfYMyD1NJuIAM5PhtTmZKV/YPrhWJ625HA1e
SZdPAz0F8Z/HZ0xJSOF4Ew0y7JL6BFUm8LV3mM1hZvc8pjBW/HEhP/r33xryWJALOVGSVMhLKAk4
CmwnBZ+emm0egUH54cZVOhZNNrxxyX3ZJ9jSEgHne3Q1K2YgSM/sK1N2aaoy42XHKSOspfox5n3A
LmVn+YHSu0vKM7yD+NU3UHx8bA6BqLboF29WGoCC5U7d1vStg54lTYhuZbNchUbvH2ylukX+veTw
W7Uq7R7kny9eAS+F7o8RKKEjNb5+cvKaE22QCyEYQOrq8C/ckL3NpI2bURzhG9bFeqSIKH924P8y
SQn1i6N2K1LCM0WPauYTx5fQy5ke2es7aPbsqlr1FnyV19wYg3zcV1AxrN3t9XRZbbHW0YX7ulfM
uDf3X0xP+Fd8JWRXinSqsB8g3k65taS7Tb5ocBC52pwe8IJ3AWY/S1vkSUIc2aagD10MDBYJwWnS
8Lj9pJBkFbQI1m45eIj1qqmlmweRBeFgj9PGsGnqHifAGouE8arCdwKFUZ0yu6P7hONdN+uf8m0i
U/n9kiptSfqOoqlphNLY4/X006JuUtmeaKHcCCYyLZfgFrSVPwxuQuIkEj6w6g/fasg0O/AWZuxf
EDVXPwRbHlAEuUL1oAU5FUtB5b2v0U5l+SeDWCrWLw5s9RI6+2CyHkwlaefI5PoslqKBsT8zyX9T
MPR0AAcVt6yH24e24X+D1NM0jGpJ2z7F/H4FwhWF9YgEKgypaHk/z9uypdLDs7fX3SOcE/18Ab1k
AuKC0pe8vVxyUsMG3eJfu6LmImQ8tYBpEDC+sXFfvUGqCU+UkIyxgqRCI2x931NoVwCKmY4oCGHX
ynC/GgbjfpZZvFHA5tsWBv9QAtq/1Y35jEHlm9cPsbWRi0RZA1/MfIWTMIdnEbNQrRux4qfA3VWK
f2ymz7SBgLAAjHLO34K4RRYzxLcrjDhc1T3kgsqNgLdO5rxekm1pxEKSWACM40N/Vs/kftEjKGkz
67os81NHHDQHzscHcC5uS6gI0WBMvHtQc3f7vVyRQqgvJXLkschkJdG1++rFjdbPePx7YE/+yPxb
FsnCsMvsGsM/XCmoIhK1QUwkYJMKQ3OWbhZGFGxg87Zo8I/LkolqbEKbIXHUjrLd0r/0XXdvG8Ty
zfUWH3up8cKHYaI8Ta9AKIAhYxUHzr5jg2ciq7QkBhieOVFHDtJpT3LfDU3xeiqTgSuEi3T+ARzv
VTsBBIQFb6O5cNM13wB6Td47g4WE3Y0lXcbCBAP7OmYyqQw/jg8WxP26dWHZujtTq3jBRuvYbgkM
khLgUAqrqPFIqbv2B0x09zSAvhTDpThCDURtwTpalZoeqw7rpXs7AbwEg7/5A3ZKGmLYN6ArOj4+
yUW7ze/0sRvXrdJ5UPKGE+Zh5P68gW2xwR9fnznzd64HaS3fy6uKcCcCwBYIareXKBSgyevALqbk
+U3/ntLxM18+rn4dsnG+ztmsSFemsKADk9eWL6qjPZvk63okw3LXNFDUEsw345g0ihb7u4Y+cWx+
Qvh3eJYvA7yio+MYFDl7/Y5x7NukZnc86IjBf6QdA7liMPTEWu/WSnIFrPEr5McX+mOfQyXm79Fm
3HORffnSdIAnryWjU71BwvohyWW9Dfj48vBJlFgVVnlxeKLiM7KJNxYbx6DNb3xXMtp381EDbeMD
gWPzvQdwSP17iN7XiQkEmkBNfB/BiSKWmkwfr28X5VMxyeJSt+loly4xZoeQGtiH8Tamu1ZPSbeP
/U+dJQFo0iNODgw/sLD5WRs+8eWeFFAez2MzGFfB/0PX1+6SWttuFPvRv7CLtQCn8jVpnktfasZJ
zs2f5p44sVSTbnaICaZb3Ksm4jGRBAu7Z5vV3fmznqGt9NSOhciHdARjmDA5t2v6441KAnbv6nXw
Q/ba0R/FfiZMezfYFLDkkFWGxwr9Av7EMQc9EKxa7E4niVd/wxCqztLbi5JhlTWe18E145pft6LS
7jF8KpIK+VxrJkxVWcC406bf10gmg41q7Cv76p53muPdN081WDCzjnpwPGWjct+hrgmTWp0/nnFd
upkHDMFC2ic+7By9ULhvrjjPolntdF9WchHyLXyM7m9IKir8isiajlLCZhuk7lWK8RbnPUWgWkI2
bLhg0kk9Ca/bl+dY6qTEpRIgV7lQN3C2uATBS6UznbwqTs0QrXlUhroWpG2z3Qm+iTAQ8TbKEStv
V86+jjcu2NcbAvGJU6Fm4p9yyM//aEuUeejziv7MbLtXyRd6x41VZhpopDjmgyoZNOEFfAiQsgqb
MqROi6U1mKeeBJGjm5AWK6EIRoroF8nbydPkD4VTz9Jjjtr8qA8APfOl7OrRjAmFhvDXtQGf/Xmn
vpJUZ1jzn1BmYGoHZGpxr83MlzmmUdREqZ334tzbpJObkh/uUB6B8EYNZuaFBU2Hs8CQ/DjqjmO1
riL5L1TwtbUTLcO3G1Tfh38et/xjfKYcmzCxO/dVR0CayXGh4nJ27AxnRRkwds+b09zJuI5cTzVk
9n5QLaccto7/Sj9uvdlvXU/cmPu6DfF8IVjkUK1YNhDE0/EJvBY9aO+BwgYOsqCInLlBlM4NwDyM
d63RnO5Dh+tB9btyJTcYpXEBOQnStTzoq44bQ40goEx/eYmJbq71jcDDc9skOrPM9DLUMNFSiIb7
ohqQ4QnDunzE0MCibXAmCtuQOqx8eUfRjtsE/0q9nJ/+cqK+gEWFDI4B3tvzmYWU4mblxKrXbLcB
ZDm9m9cSEYvJG0hkC16MAMMP8ae7QQgt1wAthuXTu1SguFbR9dnwQsKCtfowcRTb18lQm0EQ2Gy/
9FL5ySht7/Gv332XAX+LQEDOtGTBmBQ4n67+mOlsJKyg2MOFsEBS82WOfVy1jIb7lI9lBoilczKw
Stl9nB2HWeBwG1gJX9Llzl8Px/wLmBnJWSk61ydjT3IRmfZWuUNqUAW8rfxATOvER5itwdoI2hnl
xJZBoh9dE6Fi8H6MVrIOMJ3uWV4sUXP493BU0/Fau4OQ9MSXW988p4K701rk8W/OhmtcSS8LBGY2
jn+BirdnN6+PHJXOZ4SyVBlpQMTytfXV2q/AJ6xVKQFGREKgYNfzWSxkBg5G4gVbRoekOPlLaCvy
rB1Coqr5Y//pqWU4NyHad68wjETufdYSSleDTAX1s+XIwFk0Nw1SFAWVSHTideTYJSmlcVGCV+hS
Hml17pnQ/Kp5VenYexrUFV5JpicpEoLmAnhWzAbI0YJiVW7uxNXr0XAVc8v0E7QbqrBxSxoRBrEW
djnxVcLn95YZOF6miOql8OtLn8BEkbwI96TSyF77U5M0ICPVhd8PIfnu3OABGux/0horA3gsgYNM
TVEJMXPdz+TOk4MIPd6iOe/oT1vEe1nFLBH/GdpcQCjufKNV+yV/winBdoYcOKhESLJLOux0Qe2e
/AQWJlOydZ066aPubd8nrzgu7IGPzLHuGT26pbmUua5AvW/yGuX8U1A525fcMHo1kwLE6FF45x15
oO7jFMDwxD7mVtg3ipkNTxD7OTKRFJ+uobrhxMpHrfYNWz3CL/2lAQQafqoOql1G9nlP9Q+vBF9T
PleHT+XTc6hPDQBNx8gx2zA4IMs+dJRB52METrJW2/n2RDlVxwxeB2M+GbPywWQa3E+Y5uYxDHPI
VhtNcjChSW79EjNC6UxxABsSzgZlpD3pUtblPckAfOTCeyjtC4eYkfwdhuJENOvUzeBmtVhAbCxe
ONwb2ocZK0yN2k8Ag6jcSZn88EbG+0ZFXvf8KGsnf0KMTg3uVfNQaVGKnGlyra34TBEJ4xh/o132
zVR3OOxSkTd9YvCjHl111J6FKj2Stda9ykFFsAGlUmp9BK2/qFmH0JaXocYVzopw9SKfqfPyDiRu
cLmAu8slO/Oj7qj2fsvfrlfnm1Na5JssJuVkWruWgpJdt/UNOyH5887dCnHj50JiOPRIPciaWocs
7gHW1KmFIY/uddZrOxDwgzvp4Bg2nhUerYIT7+XZkt7o36rRW32//VHN+0Aw/4FgsgmiVjmisxlH
65U4R0XC7Sa5NnVMDdlGwjGPoSLmV7AzLDBIRYC5Sb1dcSLvZiulYHv1aBbrj++URo2I4hnucDuB
214LrvSQysOpEkS48i64Fz1FtuDz7VB7I1D2y49A4RGiSwvon/oPqipO/zQIH5EIrUjcf1wTyKg9
lKyhtGy7TaT5CO/vw7wZDpMPAQf8gGuQakymek4zexqz+B2+c2YNxKwcQNzfgeE6DcO3KWFREaCq
1wyuDGHv0c5Bre42rLQv+oMTmKSkvbgqA5Rkkc9ikcemId+wPhoCaB1koHl3vwGCA3LKFIJ2psIx
3s72Z4FIm1hnyrMBBERSOrPccq7VSTxBhLV67TdiWCdbLBXBIl5c22403J+VAXuskGlKmUWm1Pj8
VXGW0Q4R6qke//RFRcoqi5qOuF60pA4k/SDLiGxhV3eksIg/OxHZaeqEFU6ThV/d9HUNR18UPaFY
ZrDC8Yi7EjjbtBlgzgFrT74KfzFbMfItf0K6ty1Vnu7+HGc4XOp55UfrwkMfLi8VTgBhBJB0Oieb
RibGukKxDDnjchkeWHXJjFB0nT0cilT2aQv15ehOob5MIuEawhTe80zyiEnR1YG2Kn3Ku974V284
breqIcwGFQelDVk7jI7naNly7ckk5/wqckGQZjty2Akihk3EwILlftBN+AA7b2ePQi+7fhWfNui9
+0Tz5TgHHdU+/pV1nAKeOuog3UaiSAwV/eR+Vd1nFM/+IvFNg7ndUQJOhpXtYwHkJUNCbSDk5fSG
h3r100wNa1ePpbIItqaaHWwGjqk69vNg/RCY3CBBHTdEDv1eVWYvd14MLLWHSNP0v3VPz9wZC6GS
W3+I4oU9JK3PAYvTxdLDG9ONBUKabADteq0mkfZObpgw3eSPfGNTgYOYKz1ynT1D2Smpl1hn5Z51
PiLirZQ3zM7IOoioaumgwvCnGogbQOrmxyKxEswGgxySWzlIv8Ho29qMSsfsoF7Uvt/VB1YGC0El
Sy0prVrNxlrKJ75HxrPvCyJ9sYECqLmlZKQjfQricl1eFN5ZopEf8P1XFWuE9KQsCCRY+S1v1HpG
+ROnncS4xZSDtW3YLnIeJfBvJxlr3TFLOAQDismQp1UAAtLYTcGt0OedDgYSdt4i5+4UmqouTLky
29D28azikLy1aLJie+ohPmYCDoPaFBzjTdrRb/rjU59dAxurKgleSnJqiAfmw2Icnq17XIn3SLG7
c0rwQXWRvnmeN+MZ9x2KLsNxg/IOrUgJWDOR8U1cBnttA/HwG+IDu+ij7DObBFedWRmzOGdUQBtM
Z9iL323u0zVs3giEYcoy7ZUV/F9HbEtk5jKrjRirYW6lpa7lSKTQj1jKw+By/SW791eOspnjgi+Q
Fo3xEZKcYW3gKK/eyevQk+76nPYLDNg65VS7rFilIa40oI2Tk/ZdswRaHDwkWDbkQyFnthQS9eV9
sn1t0NHq+TTMCe4degyUJiUWdiOCkJiUXDffs5fXjWcYyM2PGJQ9nyoRYZJ5ZKeiZA5fBAtP0Wm4
6usJPehQ0F2CRjxvEZj8RnO1hQVaxUevwljx4urTydQ79R7WMz+P64YcpHXvto31qTwTQq8vYqKu
oH8M8UrMPmlzDAs6afaPqb4G/eEh8TzpTV7dwSO2ndDyZpEyvpSNxSmf6KZ2Ig7r1SldaqAImBJm
yEPIleOTfzxfQLeaMz60mFIb/8P9/dY6NoIa3Noz3QkyUBo7oDLXS176bK1qUalxJAMQEuNBzMcw
/VlYikT0/Qc9I1341EtbhehemS/YFn8E7jDnGk09ThivW4Jt0lna8M4OrJ3K5ZPNTcNeaUcc1zBQ
690NMRY3le+j1mzafq6jooS9Nyl8EF4DRzrcxik/F4iCHBa4oDkwuvQvQf4cBlxzpkYUpfxIfba1
aaX75xeS7TOcCuG31Kwr4BHjIkchUhVgapp2oIs1idxavecj6cyFcnZhno1S2uLjKLfLTZI92i7K
yk3mB0zm3M+K59pMLcb3r6HKhKGq0okGcK8V6bXzL20OXq29bzmqSkiunhL2ORBv9A8KiUmDoRC8
1zS89Eur52fra6IfKWS36+mH6VmPapgUVaPeERZjugYTQneZzoFk8YkBEAfssIMRIdiOLQn0LcH/
j+h4V3Q68Dx7XEmsxbnsxAaOTfNOW0uxcGl2mF84mXR6oijz7zRbO2VtKQA8GwOoVWV0a+Sjt/de
1QJrcP37mfpSbAZ2SyjumZtD1BJHrLyE2+mDGzawLRByM/JLiTwD4+/ltuB/Q/8wucK18vTJt0WM
VQnOgfDqEy3P9xL6I012wYDXuS+6GoCd0dNWTsVCSNzXat25/yLBzjRXUXbmcnVSnljOeyQOxxCG
O086JeRQB9Wkj98YNftIx5ojmwRbav/bxulaNUv3HgJO5cPN00WHA/DwfEi0SOZnHopoKndPC8Kj
TBFvDHTlw26PvJHUFhevaYvUtsgqx0wdmWbQ8G+GZXOTbToxwQhHijQyTWX/n0aHDycTK704F9yh
7sAkdDYyOhkPSMo7ak8ocM6NOkoeklFEcORHe8FHFiyDZiskvPWJev+SA/9VJUybwqj/DKr2QWmD
E7PYnYVTZ3Dy0yH6sBBtJAxZqdyIjCF5tMVzFA13eWMLzV0RqClBG+kSE12mVpmPAiO1fcP1rDLt
R7wBW0q+zuWJAKYyH0e5KcPIOD8n+xRaNQsKDORvDZ2ZxZRTbn9C6MFAQDfrjE/LPqMI3hHAM5bZ
RPpC2u/fnl1dRQFx29AUjIhSQXHVasr3oNDOi61oJgLBHpBpC4+inphkQGOO26WqI2CPk+GeSk78
X6ItiFVFOA/TauwbDrlAoDE50yO6zkodWwqN5mvsvadZmL36flFfEaN7dinZbEe+ysNdh0nHa23x
8ESpuN/WG12PVw5TY52UFcSoLonWoKowTNhDqV0lWkHgnb4CAmFlMgS2Kuy7bjB4yXdLdPK8zRPn
nx9ELeHm5hyoAVJUP0zAvqLaFZfb8RdlXwy082yeqAw1/Xr1xlPNXV59aiiGDccZaKRBC/OQ26dH
+CDp21yliTzkuxHn5Ad7dlIisGZp65shPZmMyKoLsgk9372Jvc+xjkf9MS/TBUctlWR2gQ8cJkgg
6lP8VWyjUZS5X7JwED9U6uTJD+4ZNJNfxc1Y5+w6MWhZSYzq9tlCCZ8G3w6R4yGn/PB9ESSf/5Hr
r5Ue/1roILMdZzAzmK5FFMVpoB3CgyLm0Hw/wqin6p7HWO+NRMG0D3R2kY/77stVzd6eqyjB5ulx
Wo8c6RIdlgs8UUWs7Vbi530CwWlq+aPXeGCGW5CF4UDqg8DK/n/hLqsgxgcFeNQk/01nTZYVdyZP
6hiaJ81bFz9BJcnTHI34PHDS2alWDIX6hutmD/sOAJamtUezNJ9q2SxfiIeKGEuocx8KFuuD+BKs
yh/wXLLiLSECy6V6wzG1AuG1ueN1HiV0m6pAqOWA+OeDjkhgw/kJdAJoInrMDNhfVf9EkLpHdAlt
dqcRk4D34wwsYcSVIPU+D3Yb6PzMHb2Ur2JjrypCV32e/mjWYP7Fg5XYh7xrmg2KhSEVCHztzXwA
qtpM8w9eo6jEOoS+Dx+/zc3lSbkdAYrCwKpJ3FJbBBrmtbfZqbFqQFCi929QIaUrgUy9AFUmM66L
vXe1xxrOMGuusbDc9Iu7odTAxlTDUL0CqUt3SUDfJWCWsyBE2jnTD2RdWum9BLxnZOYo/dqxhiT6
2rAcMZ3aNux4EFWaZo//Th9+LHZ8+ZvHerP5Y552TMZcnzeLZoOzh27MvVIsBhUmXtg/AzNR6KgO
Qo6oqODWjHhIFZFl/cbtxgLFJ8KhYvqgEFbdmtUWD7QhQm35GuXFeVUX2Q7j+RGx3GGhl3moh27a
l2fDAcEFfvXOTECsa2ekIbn07KyngplArf3vQW0zKugsXYsUPJzAa6TPP8nHy/hHwdH48JvatdI5
pDoBo7wendVsdqkpCwX2PTFZLB342xqAmNspoFlAjDm9lTojNDzAt6TPX37vSp2zQ9YtrwWMfoHg
vZioY0CKOUxrC+y5wo7r3RaNho4/L8oiC/tcU7ONfhlovfQ2WIMF/Trdiyooa9srKDF4hOJZYbC2
r4HfCXNUp6yTsiBV0ncZ/3wtLdEh5pYTQyb+c2R2A7DakQ0fkRESUpzM2S7wolG4onwiqdfR/4FC
wmjkJC+l6I8amHgY68cEfDmkd+dMWeX/oS+8q9tZgWdU6XFb/Z8PpVGPG1ZUu2TBdy6Zep5QUEci
22VP6ofKUE0EVzxNZ3h1gCd4XVVXNlEAbMRgofn/zaGKYbzGjVXYiD1+D4BqFagDuQgZQfaML6Qx
S5nu7v+pgLkH1oYHgy2M2dX2aWoKdKo5iiXN02y1HLsnjGawrauVSpu/Qr81cqJOoHwlhOMC8May
SzJkp674tSEn6Qa1iZm6R6UgXam/Aol+3GgIVs3YfrIZ0oNHh0XSa+xNGqAZ7xe1QU3a+OF9CLpK
jKicZTtkFnA3rpWYVm6+5zneCjbPVW81PL9VF+yrTqkGkdGqarpEuHVhTjVHfSd5FSi4Nt/duule
LJBg/loeiNxBCsHdwUJQRbn4PMA6gX/WS/LUNjzz83EkrEdkypDVA6Bikq4LXwB1suMuY8l4XTvP
pG7DZZgnk5CyoBIas8oojUsboJ0TOiB1snCU1kBVMDUewPTHPRVxoz+zPsIA7PzQEFe+Lw/2344G
etyDItrA+TBXTNdWiEiEKKigD1IztfMVaTQqxh/lS3jVatPCgNMrvqeLPPhtIh9N27J8Y0GiAAIk
nkr88tHToPWNgIiaPoZIR81tOK8bLpdCXKGMKpv8avsAiQNdRaLUPWbrfzfe+2Vnhp75iVEKy2C2
VNANzzAiFA8DrIy1/0gWmads8cwOCL9pTiAKh6CwAM7OvRU4pvq07Wvy9VNpb5nsLi751kc/ZNWY
9hRBInHI3Ern94GzU3yUmeIQHQXl+tL7a+4gOQ8pdwGPNsexJGpkJXMqStY4Q9Oh8P3MAJa+tShZ
djlDMrnbZrVdVjQT3dK9K2OwRnjpEC9d2pc0K8pJOYCD9OPXMo1JuxE8KfU4937raauFqIttmwcf
bky59pWJ9Hly3IpZiffXi1QJKWFBlmPXNVo9KIqssjmZRd2RRVsj27cBFA8BUkm0StfyjJWsm9d5
KnRYq5sEfTnLRXYfPHZU81Vzq5PqmSYl1SwODQ0NV8mWbKt5vFRYhiv5B1bHBp/LoVY6zMgnIsdL
fRazwJ8Uhr2tgIAo0GHuvFZBCJCg3zbkG0/Q/sasb/tU4St09sLZFHGMW1rtawCsPS7wN473jnG/
ygFaQJQ8RpuwXL1lzyhFvfMMwOtqlafXhPKzcCI9zgreFmCUT/zpHMxhhgAgKrIwIhHlo1H7vBG1
LDMSpz9jpifV5sNb4ntVkAvl5zTUwsvQWM1VkQSV1a01JIVt2pxf1Sibc/K7CVbnwKqL3mQzVX4U
NLbxwqNsPe1PGgsPDfd3vgMnMZAsk5RbaipJh5SL2EfSzeZ3P6ge1AA6XOqYHpgwh/N8tZSql1pI
NEhgU0VKye7CTqhG0sI0JRLjeeY1GU/LySUBlifF3wpS5sKn0hrXZ+E2ls3YUy/uLvZ07GrYeQE3
/eil0q5kD4S8wMigrsO68y9u0+dt3Ke8yN61wHxeCEX6ggnZqelBqA/kIWNVSZ+k5Tzcepze3QDU
EINhSFuX2xpYHLMn9ySiqRk6umYNFwGwsfIkxFVxP5IWj9GY4m1u2fKA8nunxhLA+wHyz2WsSP/J
5mGN7y3YRITnGmkryV75wFUp2FX7ceGUdfF+YQ4ipZncqph/1976/O4ftNoH29ZIBIVft5F12Vk6
bxSu/BlYHn2SYAn9tcmSpi1n6qkXajyNprAjYeeBYtrln5x+BRTDIQcWR1dMWNKbNpDhPUJ5fIT5
ACq6d+frk8vzOrcw3pSAJEbPcFZWUZgv+vIjGH8hwH27m5aRpup9yrOXThNbfWBZkzvl2ha7qaS8
mK5tn0zoGPFI5Ac0BXLQi1lpKfwPc6qzBWqAQ+piVEt9XjI0KGLRM5xEm34l59ekV3OdmJi0MYY9
+FTL+8p9GnEUQ1c82xu0PfM7yARIcpbxlddSMLodtfAvw4NAy35S79Wh61zfibGnveHVSgxwObmr
/MJ1rrSAWh5YEWbGfNyPrkd+zaiPWnxW7bzKqofYPbhsg7uEyUSfTdBgmDYgH3i9B0kBENO54pDC
32ENX91AAwJYD1eNhBG08I3K4F2t51WWN4ZrcfU1Tf1pRPHFTOgPDFSGNuVauypg8N7W9Jms3HJ8
fTwx2kmszR3ZeH3HgTzAtISBpsye+0m+Gevu9eJn4pnwiegO5x9OTg7C8LiPvKzrzHW63UXCSJU1
ehbcKHMmGTS8eACnJHhQUWidxk+SHXSM8dA/RTx+XyhHngi6Ik+qaClPNNrvHiynMjsd1K0GZQxd
xklg+Te+XE6KHb/FcxXsk6LJYVbhvJ7Lx0g4xmVgcpyVt6d6ZpEs9oDAuh1ZexmuBlZUTvpbRdCk
RnKS6TnaTkhYN9KXGZujVY/agl3qmLcvvAJ5x25gkh2Ey3shdEkkixA8h8k1FoEef1hHWDdrtC+O
xWt5ez+uW6ek4XKd7bDfgEch+Rzkki3bDcuxX/q0oOj7VQLMezBpwxm8TPb7qojkOKzOXNJUHXKY
mz4mKwQcptWUhoAm2sFxuDeW2LrUmwmnuz02BVrgsy8NVrbcVxez7kyqZ5DTbgNr/eXI6Ugp0qKm
kKKpmj2/yShY9W7RjJocGcrrnIwsw9GuUf3oQmApnmgXWkvZImY2W7tmumhggDOma96xM56i2tG7
4sH2jXe9cQC96FEH67Fha3hqZBD+bJJIWwNxsRuVUxHXP9G0qQcAdNdxcpVxtG+NHlMduRp3zct6
dyB7+Qk0j/pg9nj71dbVoavfogNLOdEkVMUMe4oSjj8OtrNTnwKyTJPV1ziCEZoeuEV2ReGCXAkF
PkUELHoWjgUu89zA7lNG8AV0t046hkIpyByEAu+VclHAwvDAITZT/xR6WAMV3Bsuk3kjlZ/yP4EN
aHlE9sPShzV0rNyr8Ti4kkQfG7gaS8ofzxrjeuHZ68hn4jUPHgPmOO34mQ+CKaY4gmL5J8FAi7zN
5on0vRtj9oefqw1Y61siolZfSOqSwnVwS4j1Fo7APnjnHljDno+HJhC18UT1qWgOkFelFpSyvCHr
zpmK5a27IbSltdzPMaHO95Dmg3GaumeUt+nSjS5U7VBWQHcU6xxiZlRVQCElILUQVY1HdUvcq4kN
/76+fo6T8DV+xX4InK4LQiYBaDuuTwTAOtOhsnqtFVP3MrSXL06Ecw2BI+MNd/cLHEHHaS/cAs02
SmOHEiLX3Ebd1sJpt0NN31fOsydG7e2dOjwtgPom6hNmr+98TAus1lEIZZjYM9SOBR/67SGddHPx
oi3jvuxOrn2aXzxj7r0wUCHKTL8mS+LkzLHrDs4hNnC2X2hipQvYm9/vK4rVcqyQX+lxF5R4LhDa
kjiKpQ4ImRh/ct32SddB5z2AVXoyWG1uNv+ZqvIzcWz9HGQRfvIq68Jxj2p5W2uwsvXr1ZWzSjMS
p6eZQJxZ3a4SVpw65ZMSeJ7UqqeZAZ+suFZDCXv60arkLXbMsYqLNUvQTSd73+TtCAp5sZyeA7E1
h0zoGQ5x/fCAEPyMotHemwKfOf1a6yIuiwaN3Y82npXPevEHCAhGN+QlLc8hCqzo7rMKfDewOFs5
5xUBcQpt/nyfQb78D8DmxyvDg/gd9wOIymMrfykIjQSrV6hDLeDdzySK+dQyYcBk4tq8w+qipBD1
8S8MWGjRaJAhbCttaExEuG2X2+FfQFUc9JIDwAKgLyT06WgcDajXGe0e3MmOsoPHRejP54c9CcUb
e4G/nu3dXGw+n/QpEOdg704MY5eVTNAgJcuNqaT0qJaDKZiNpoH80bSsw32e94xOLznNZXGm7ZrB
3Nb4AuehHZLnvfa4yf2sS9ota0THGL/iFJTjYT5F2bQjzorJpa5wpwjXZVEndLQWaapAtfpGu/Ax
HmwqNl6BzY4+gYyOWQyh+eLg2d8WYcfzTItOmeU03YCb5tEo61aHXdLsLyjSCG35w4f/iA3gLhRg
vFED4MvmGZRZLUBeBW7T+Z98PzKY36rh1/5L5P3pyt+4Ff3QZzpQBbNUnws3tjNw/FZ3uuQirqo5
sGKVGWO98zoW0zNO1LSLxaBzLPBc9u27qvhWcJ9egX5dPQ4iZuBrNM1eTrcS9BCPXV61OF3MsGld
T6JsiQ0PQnqTY025C42lfdqqYSf+QpIQ44IXaB3ZvYVzF8ozUk1100xyiYNsxYgFdyWlGzJXpr//
I8R+8Ze5ntj7ez/3q90vyxhzba7/1W4jDs53rmpbUePbjoaXmFvgxDCXyiOAg5ceILmxzZvWmrWt
Vsm9BJXStmkM4qhrxRO3fjFjX9tQQRaYq/G0VXxboX7bisqkeuNQbwfhF45rEaw2wFiaK74KgB2T
WnW3Npmxl4n1S+gc3+JJQtUzDA6dN7eKT7IKfW06oYr8WPZB6A5nyrxyIrwE66xbXyuw0v9uHfeF
LrG+IxORH5PD76kTq219pHg0BL7VQ8Q8lb5vvl6IxO2VneiMo75prtvObUo3QM8VbjBJeeVB5WM6
7cASs+1n/J+JEMHFD8SGWd+wQwSpyuGtayNRA+BoK5xOnOyAiqYSwjoAuE1+Iw7OucQH7tGBtBLo
4Dt35RrUxB8/uw7oF1Zp7EFHsJEH36dhnbeic3VEWKGMdEXaWI0KP4QUmzcPnA2XZkQovQ0Co7ek
JW8JXn12VKzWDY5AsNb0T8947s+JhA2hthb6nmYFNY+g/kFzK4fPhtLmcKqv8EEAzoOZp2NkIAeL
XQodOc31bBj9CDr6BFyFRu16RueTtQmDOovc8CsOmPl/eFXOLDkU0ZyHWP1MBiPlzKPgFFNAUKUb
vspLtLOs77tL0Fg2lz9YzgL7YgcCAbrbHpmyVb6SRHiofF6nLr373nhQWsFlrkmG7LLKWqi6DUvd
FBuOLIoR89cY4YtLVAWYqliRiK3o9po0iq/WJj7D702n6VqgOdoNTMfxsD0MYi+nCgJlaTbbNdwv
GiNCXP9CuCgAoP0t6V51L6DWxGCCV26dZP2tYgr6OM26TUKqS5lMk4YJt4Bsba/4xmx/0JO8OJUM
NNu5z5X4d1UrwO2mHZ3waZvgbxoxPiq8kVy5JQGl9heMfXBJZ0ds+PcQu+B2dMpFGgQZUxqQhnm2
Y0ckriiPBQDEBc2Ypo4eyFrvY+zhK1Nr8LZWrprXGOE0BfmSi+U4gXEq7V+gtCrjiSSELCEv5mjO
lR9OMFz678tZ5wjNxrvVCcprK+KdOpWoYXqYfGpgvDFQ6CJM50r7v2D9oxeafROlwi5PZCMPqn7b
HrKazXQfwG1P+9GT6yI8GIAx55XAivxCnNYTzjG+PT7RTMVAhB83OYa+0grO/qYLipv78U1X8ug5
wAd7rHUfxHmQH4Zv8Vcw8aF1JbNE9BiixmkZKS54BoN9ovztwIbK1c9ke2/FVIu0+2J7tSnIS+S9
a62H/rTtCp61j3VykIqhNmXSDc8yleIljH+FU4hJGER7AcvY7wj2FSuiJMN12JIOi5L1yXMt3cbX
S5/INew5sU+FaZBl5Bhy/mUiLd7zp4aFdtXINrUTxMTWmCy0ycg1MhWnq8XcbHi4LrTSQ5ffTg7/
x029HqtwGtbaoW8MkUCB6cK+QId59DSps5XUh/KMi9GupXXFX7cGoOn2kHoqhDamN2wzQOzup4XU
9QcuYQvVgGxTFv/gL/RN1QcvwsLlPEH+toGU1VzmxV1AjZ/d2PK5GOk0IW2w3bpbmtgXGTnqWBk1
K8fAxwGV1g/XDTD+L2wVEgD5GqA/dPhLdPi/K39w8LAl6Gjbxy/jAUcmuDkv0dFkF5WqjtQvO1dU
RHSx7Y2HkN5oGQQFJP5zb1+xBSzMr7qy6/uOdx+s55YhA6SWC0+bIFFs1Vevi6N29nz3bMEhDl2G
ekIb3VuxNyF1lOpQdlvakI1lyj9KoQxOMcdDrDGO9UR6VmWWHioQzg3TkpYHcAfmMLmTrbqqCqhb
tvrF2Ua4c04O2XCx2HTIHvQg9jsvG+Zlo08TmaX3Ug1gAKLRj3flHpPG9HrzWPvIA7CL10VVm/f4
R4rXiOKvnZx+MmozTIQ9tnrVWDnceu6Yo0SpeDIVNhOQueqChnyqqhS/DJ89yubZ0tOHaoltlCPe
37yKX/67fxcFg9O7+kPqk/9D/0TT++dLOdKmn9uHn6YxeUDdcUJHr/NDb1B2An3FHYeGHQ7CD1CR
5I3cffYoey0RqaNz6vBfBaF5UWpKgbnL7gS8qqV7MYtxizJEryGnaPxzaS7aAGP8AXfQ4HEgBgEf
Fr/f7rQxiX5mJFNmEPvPyL0yU+rduQzGcIk/rgg8U1RssmXII1OVteEQ7rouWAPMLn8gwSApvrA6
JOSNq1YTPmwN4L5FwyHmvj9d3f0ZSi6wWDc+jGNrP7BUnHu1f5gjcqkUXuDfgWtlU79keh655Dma
NOUlGgAnNq1rez3Ha7OPJ4wIffVuLWz9X0n/M1jHlS5cv+nSscw94DLaierstv6K3E1mR8BoEw9I
h7B9tff1Elz2LZ1vssAkaA8zSCvWsH2CSQjZTX9h2s2JI3RD6y/gnHQqU7JRaYdrFgUmM/PRAq4p
sR0QTSoq1FS05AN9OImEKjmY21+xn7qJYoxOQeYv9Sq6b3nJUxT0fww9Kdy2HbVVaHT0njkfLloj
amkBoAA+dlEDenEvG905dSIzW9UzWSwaL2jy3nBJav8MQJ7YLAXOGmfIkSsJ12PZhBZdcPOtZYwL
hUPXOfdZDiTD/U85PNLUlSdPLGhAuDrGn3jESB0vmO98GeBA3R+7f3v2Kx6S2VTXKil1Nw3UJ1Ga
aoPWCW7gaoFKC7l33P4c3PAkYJtISfTIjScCyaX3eVrGho57joKU6IdhOR+I+yDJzy0eervnSM5e
S9Ty+gvSXlTgu8GQmZMphHblnuCL5t01ECy+bf5D2J9ciQufUxDk20faU0HaKspcamKyy1bbliqa
PuKLzLT/43zQDf8Bm9TZctQNO1jr8QW/SCoX8OeG9qZr2b+u8r27Z206JsLE9VDA2moL1X31LMlo
nyFQ2O44gyfKD4w/Gj3fNdiCzBue086Yzt9xf2wqTtN0+1X6/euBtDTxeBf5yRyVZNMYCyaTgM6h
H0A+azXKVP5TDnvUstFEXANrxdb0pEACCGT4bVjZnygCg5TgGtLmtzRjfgLEZp7ggBJqBUCdpM+r
kxr/zsfSxM/HZiOdecticVTUmlsT529PywplznTIZlqxwU6DvR3EBkHPvNyFHDbx0fijInJlpGI1
kPlOoHpMj840U5yDavQursCF99EAbb/TyZn7enwr4vpcq1GWtkumzzdqCxD8vmXCNhxHbPLYktIV
+/UymU45jO53B83bIc0AK9Y3l6YFkI53NPNpSdMehtNsB/grRnMcO6PBRakND08y8P9wCgzB7tYl
HKgOrpfyP/KoHo7yi+o4XkuN8TFZ1NwUPTLu5KhFWdTbR6tdMEufLf2cIa+5xS4m2iu0ehCn4VZ/
KRcHbDxWN5PPgLtatVxNOpfuoRYkWOe5FdDFdN1kienYciKZH4YP3Cnh/gPSJDc0rBBhuK0xHio3
ZGKfSnVMWBAtZkAkCrCXenNhQdnD5a0MqfBq3/lUpbFxyJOg3XxVwqK66tQUmpixNjoyuEv7hvCS
NbXrlmkrL8U4IBFNPcHyteCHBYH2kH8sExWW65SylkPHU3AIUiQFsqq92h5yAclW3WdM6BRfUQcw
h9RL7xtK/qh9ZS1ZrE7wubs4L+mXDwtK0cGY/+zX/jwoAzuBd/9NPlC0r5xIO4q7tv+LHpJz8ueD
2ncs+eFTGIf/F0QtwK8XkhC0cKDU7hQT0f7wYn4ScdebMRJc3t6yH+Lp1gb2CTiJT1Gti54cQDu8
la9UlQYLEC3ljH0aixNInLcB+jaW2vzpBztfP4MjdrqDPU2V8/o6oysgbJZVix4RCMdEANoLPbda
yw5/BdUGuQ96xMV3tOcvuYDtTMFuFkVysdTR2kG55I82qtQ+ay5eM2KISanYq4+MzqGg7cXU2Cf3
9TCH9gPvVsjwCJDkhNbRCLT7zVj2wXslnMGLMkaGl1rzO8HSaWt7CnCaIEmloBJRrw9tm6p9Nkmz
btuc030V909i58CWUjaxqvcVSNBRi9UnIMTidcnWrz+yYIOl51obpKNxjWYRFipbKWjSmWwQg1kR
VmgfoQKJdb0Reb9KLnIR3pvRUMGHpM/y7gaXKyZ2ic9FcyVe5rrbMM7B8A0QrS1jQCNswwnW21u1
uT8W6yyyaqQLre5YICGyMJ4e7cmL1E6f0K7CtCL6p9n9bMnX351UVvpCCnbSJIRXTUktoCtCFuyr
Fd7lfNbwB+OxItXyODTNOhuRGXMmjAo8ZLmSK0+BsedWoKuERV9oik/IUo5caeEaEZUViMc745fN
QB+5QaADiE96DbCQHyec+uxuU/135Yr6YQ2sR2L/nx0UPCLllFZ3NUWuKhPQlTbUYj7apIe3a09W
6+TsCIoBc7piHbu0og9ccS+MoJL6jotoGiyhsbtzIluVt5vZmR1QSA0ZrrLue7xwk4hJSbeSuhgV
QRv7MVTDFuSvvUjOMWkCZGKbRoF25jsT9Qa+kqsnnMGx8zGn8kh5Y5cRK3vyPbmKbO+aDMLcNEJk
CVpfNTfROg8IUfWWOj+nYfIwL3NF3cmB4njb60QrzQIL/yHe8SwFgocJXs58RtxQjMtgeUAUKv0q
yZOzTKH0fUKFsw+fqcOF/JYDIYT7zP2OO6VAHhsRwjPUu8rF0o9UPx/ae/J4OF6hPAC55q7NvHXG
k2SChTbonv8t2Xd/Azd8YHkN0A1kMW/NCNZilY4fHprce30LhfqmKLRfqiZD8YEWuCgxLKbaEhFq
apSWFLc4usGuvuITM1gxtNPQXenie+lIiGdYpx7cZG/OpaIdAWGPGIIxE3bHY2PuT7idppcO3L6J
5ytZZC5CMhVDlzWbfER4LG7ZJWnQFjvxxkvkE198l9sojcut5rmKhdtfZlhseR4Pjutbb7W4/5kE
nPLTahff2X4kbJInskZaEl1r3jFqqkXHO+nva9GOi4no2OnJ9bAI1PJpQRiXjaijJwry7MOqgjko
jsR4fQbckPsiz9CUcehYzp70NNVw929PZsjfpn+fB5/WORC2St150lfTaPsXxaOJwwsz3H4wLNcq
7jO97Pd+Iovla2C/c3Oll1wg+gtKF8HRM8yF9ZYg72sNVfkON6NeWOAEupGDDuXJcsulMF/3VgbE
NdVqlsyk2Mo3eh+QaL5ZBlohGeqC7AJut68oMavsGYh7Oof7e+BzM3cCinyCAYqgPmqv9OItx3hA
Pt7qNR+SQgBrq9der0MOLW7+2R3jz142ugLILWDdm9tqjITW8e2h1yJlbQAcsZ1QathAkC9WyMju
NfjiKTx+zXS+c+jTex9n+zh7VDMt89V0s4zWWqWaMLpVSsMI0m52Z6xBQl8JMX8BKYJEuZjCG78X
Ds59BYUPRHnajQOKTjE3HUoAGECGDHKbpmKPZaXu8J8ZkTCKLfKwylpmArdYXlUV5iCmUdMEDLCL
7R1MjdLyLVC8jdN8YIzXPGO7GqvWoP5DIvBXi+vm1DV/zTRc3DCsv6CGo/aTGcUbxrLxFNK24TSM
gj7mEyqMA0bGnWdv39GLrwcv3o4/j1/wng2+Ho1AERKMuotbSaqg2EeoBeI/C200Z3al7WsD7LZ2
O1ZPMAyukUiyhgZH/s/sWR2rm7Ec4ZNRpOgEB4TMC7xdvytxhQ5qZLj+PgjyZxrmvASaokmwD4Qa
SHnQ6hPFDTngbFkc8gvy2uzG3wLTxOg1d1d2XTxcHSpkzMk6xo88qGBB/nHgkP6uGnvrPULSO/E6
+77hKcOByFv72IW0Mov/0+TIzB4wxFgnAjSpucI436G2rRVbPszIi3ZWA+I6wSXrbgQdNDP2hiZn
G0TWSBiB/1dsRMzEDpkImo2zVBdQOnQG4zFP/1Tqwow7sssFAEXdzrtOk5Q2FcH+yFtSzw1Yp2YX
e6nWzhtPhhuwkUX60QYB4LocU8mNcapOzPsKZjuOnatr2sB0hirXVrO+GGYa20cTdclVNVYPKENp
K/BIJOHcpnxJXi5IBmIWWAJDsVRuGN8aP6aGid3ZANiX+tAlZphwQbA3hTIT0CX7VIJRQCppmRCp
A/Axtmk/2pKjCGwMGImsZXwhmFNbWeXsQlME9104ZabB/3gRWyn9fcScMHcHsD7A8qhRG7fnEw79
QUjf+j9/Qvxqy/JJnQ2Ahoud4NSR2EUvCCL5gNK66RmQcyEw3sL5OBRZ1DtFcSN9khK10b/TyrQ4
SDNdBI1hGVIUATeaJ9B75wYnzTujqBhjsy5hgmfPK9m5cRrumMNlHAK/QhvVoYTBBYieizWZw+wH
PUzZ3Yf4w30vYsjsq2AtwKeybA8/KzaNpbdR3+j/lx91+kfmK25+NwDGvsiODYLKxwtfLm++ggHZ
YwjYCH6/TsakVD1F86iD8LNAdV+R7gIHH6VgAnJiwjmYk9wbrKBY4f7PKWFUgyB8EM6wLVKK8Jzi
1UYTsmE1mWzwDx8JqHAauq44qmqU8Sbw0ZWCcJtA2qtHmjQ3PDbwLY7abSTOHdcZptiiev9k8hXj
UT1RnEuvQrxTWMCnFVAiFr/JjEVJxOA07shlJpOCV1BMKQ6dZT0oGgUTOdDLbWUvbA6AQ8mY8/z6
MZurcyxd5rndR7nhMaKuWgMJjM6x+KE/3sR0lShkqNN3+MPNbXy2HTEnfIrNBRk8fgErPwEYc+WE
gsvFbZRyY/jaF5O3YrwlIF3KhODMszASL5e47Pd1DLrCo4lWPZnSE5D9yiejFnn//d6WuzKCcuvx
qdyDNSmjLVICMZBNdz7C9DL9NApDZ++FiLtBk6KMOJh33OmIIsDtpp8QFPd7RBC8UZ8IEZrde+q6
eFtK4zzSeXhYHCMFm9ygBSrPpIkOOc0kL/PSWvXLrrLU6wGoD22yd2dVFsKreNdjgwcmqMmNWPIY
CrFjswKQUWZtIXnJzrSkVcjhevpOboy6mr60Q01UJrAEkNyCUbNROnRPYPWqJ6LEh8IWGXrXCxE0
5eXBS17Kpu9+HXVkOwuYRbZLRPkhhf8/UEifZJbejvYpQZVQGQ83esk3RtdSHTFi6pro8oA6X9dA
v+hUUKtjHPoRoumOZdMGTKjEK57yECyL1g8Z/BBAdNrQTIsGiQeEaESrdfZ1CUKX3a7CajGevrf0
K88d7/5QU68X2gl7eFVHdZ9L8h58Du2lyMRQ+0P8W6L9f5WdsH60S7xewK84HnZSwZAu7Lluf59h
sssxmQHTMaJJ2HTeifcX8gs2q3TJ6+KFinOUH16LROBczsYr1u3+qJNdLxt1/6UeHHTHUTiNDkcT
UufjtHsxp5bwU815ExYoQ4+ZsEQv9b/DHi/plCoF5mc7IEdYZ1br9IhHs2jJyAYLVfsY/h5sF29O
NqV+1B7Cf6ixO+LjjolDo3TWnTNF3Y41cPBh2jcvZZJZY+3Xq5q6qlH0q6uWNA2z0bQIsO4ngGhD
2TuDVzjmw9scO9tx1XiYAonS4xiMOMP64s5eRhdSCCzzNXqEJ5UVpVBDopo5fvBhil50y3poTrjc
FxSYgEkCkrm01rL9awzauzwCsJ65t4401DROT8ZKX7B+x9j+seAOtE0T97LIqD8VXOzKA8/km3+8
B9vVAg8u6ipsXM2qlc0jQYsyHJ+od11spxl7EJCLK1gHAxgEp+tPeYmUc9ir00A4N84M54qlj1Q2
WPxbtTyU82T8u8yPH700zbaVxl0X607BPEItEVZArr4tzOC0HB4RB+mQ4wUdINWXYOar243/fQqr
oTKTzsaeBgVTW2+ODZkdYDnYDLgf44Qx9g6muDppdvojxsj+mNgslUVi+nftNZa6LQP07k4FoKLQ
zz/tpJnb3f8jG+QAHrgBpTByMl5GcLUH/ZEfx890NPbXbcOHkAkOR8JWULyMB2HYmszI/+K7SzA+
vnRUTOXjyP1E4Jcu+f3/BYJnFIvmpOcG4mUfci1u6BI7TCaRZ6/JN6HKuPfCs3eiJQ641orKSjhu
3fWGGpxnAhebpdVlKjuyTBNDxuor78Lu7OppNTYHwhMDkUWVkxawXY5kEb4EutIJVTPPtxFnlU7M
mIJ3bGoWjXyYcz7jiusenKJGg+0fdG19tYNJk5/0MXPzaR2lD1JqPdeDqXZnvqTIFMT6wXF+lzSb
Ib2x4PTUeZLuwm9i0KASYhpASUeiqa/n8N2ggxdhdwqyWVqg/gGnhNFaQwAfgS039KO0+cmYdSKR
sc/IUh2dkHcDYF+/EEvzXiB9mv3V3MrrfVJ2uiSKsGA8BvhAS+u0lrpw40JHfBLZSVe01fEdKiIY
EdJ7hoxRXavokOA/Td3ZEkaMiBM5C5qlYXWnVYfBDmf+c2ilwwxlB1yw+llWAhd7gw2VaF7Y5vsQ
zYZjt+OoL7NvImwrDXo6PKXaK6Dtsa8bf3LWGHSdc3KmWpvnbwndau00jveIpMFMcmtcvms3H8sV
rTHEIn2vqGjBl4nubOWDsYEzg3VygKrQOv5InKpJlqBsTPZRbCt7fxFRmt30se20B8XRZOY0lvAS
IEVGKEQj7wrhGI0hvYNSGmr/Yt6L7aOZVF4zm1T5rJV3LEbdrcS0pVNcyutW5zwI+IocBqzMxNZp
DhvftjJ1Y4AW3PZFRgGP1p/O8DbHN0VFLim8ICKuxQMw+2oYkArs6RzzNkTuYjfka9+0qscBt1PG
vN5E1UvRB67B70+UcR8Rk4xUiuWFiRAdVOpjdSkAGbY1L13optt2Fg0vt1PVyccwK1UHUnvYhgdy
Sdqyq+yIiyhiVhA9+guSZrDkkib9/Yv5dKWNOUyP24Y7cHRoA6Df2oCX8ZtfibWTLra8kX2KVTA+
vBLAh7z9PRsLD3ms4LDk2WL5abVtBaCZUsKQSz7Vg6upGOLgHs1F9cnAgRD0S6rxfXz70iEjxEBm
2eMZCtKibpeoLbwtGaQZEr8zj0ZOnBnxtK+hgiiSIVJCr3lCNapKb9nYzu5upnN3OMG9aUGMaEhB
MGL1jQX+kFmqOi3ugN9IZVwMYS4Rkhg+AkSZ1X0qoTeJ4N4S2JpVYw9KUBvRj+gkzT1LmwHERMr8
nfN9ewzyYlSRW45/4ngmGyuwls8Itv7shzCg1s6+6YhJWuXeYNdZ46NiIvoshX79tsvyKcOrPvap
lPgK24K0RieYFdFd/EnRBPYH2ixmvD16pLWIBj7LwLWi2KEINP3z6AKM/EIhSZBmjmQoUcg0XQXT
HoqLfFJm8n48wCukHiKqcSwBZAf4NFlmtWPqAB+QA4LFUlYCMbEUzKsFAxVd3yn5c1WzD0kIytiJ
b77MKQDepkp6EnPHGfz9JNAyB8767Pt+Ks6MxBsW2gUOCQ8IJvU/O05C2lpom0QMEkwOm2gimlwp
gEYKaHJsAmQ3ZfZuzc46pSDkuWs8mD5J+bcS8YZsdzVMltcOIFIu2lDD6gxdV+aBKa/6l8rH2mj7
c7rb5RpJeyHeKkWBx+4PnTmxYzzVpEnhbPk1+GHcV59DwO/pAQExI7H7stqX23JDfXp4ZBFgWP1h
KhvKbUtxFNG091kkVwVQX8vG04w8SPpeHrHYfVwQdYzDE+00ZnvrdBwGNevR8Qn2kLdi4MtTBiQW
f7FlbNNwJKuTAzSgGcRidnojarj9ZW3IomjgFdzM4TvSBQvppEjQ54AWZ+S6yZkqnc+eBZQdw3VG
8dUnKKb9tlr9UOogqE0r5tQAIQS9XwQIKP2nc35ocsxu0ozzFmATGFcAe7MltseJ34TuNMslVTWi
GwGeupJBZQ7ObSPHZtZD9N8ddfphFbgjE387kZx2sp6vjuU61yv61iNBQ415dvg05MMXFRlv3vz5
xT4qRd7YytBDfNYBLghxzVD6iDooPTNzLKHyw0kDWXl4XeEzOqvwIac7Ig05D0TX1LaFXcgWspiW
aGnwTwpuxyy7OA8BZqz7+p6YqJQCQwzJYq1g0dkaQ3chlfYrNs6DSV2HUNsN7uExV8gmQVPDdi4i
XpGGg1ayekxltsLJGgUAH8GG9jjTiPacBJG362jx2KIiQNU3DtC0b2BXH3paQR0kJMaEckCnOhCx
t9NiraTW9U2XEXo8yuRnSHV+mEHM/VGM6YMP+cSqI/EE0xvQlj4zGAk0GQ28YLu9SYQbs9sUYrPV
EAq59/EI65nW/qtbuS7WxuI3YNVai94F2GvtKy0u+iiKGPdtK2FRuMCKACxMVshICdCtTx673sGY
inR2jI1v9eA72x30cvF7Wq3G0S1o1K3ImV+qv9OujG+YQ1uTdJw0oKAnfyHukUZJ6FnbxARYPb2D
0rC94VMfNMrpjD6NvcZ9gUbUtzBuqgXPW6XOi+QWw3qmvB16AXtrXtY+nXjtS4ddhvHhRUZIBhjt
CHWB0kjn2xPUT/VcYuQ45xis0fLZaDs3SiQExESLZeuoJPeZzOo9Z7qhyDKUwbIzku4BcT2cITJL
LZY8ulziJZ2BpjoLGb1CT/wZeBCOXmFBCht7m2XMpUQ/CLHy5MbeLd1d4u/DP9wlfF3wPaGDa/Wu
U9rzEOWOGO+zCcA1IIOK7VeUPI0kkiD6lIjDTcW1Tzh1ofCWBBOu1DDv/qmwDp5OMTUF2NQg3ko4
/Fw1WfakcCnwgkLrBzCGQu6Z2/KHBOhH5Vx7s8pglhY8GVc2SclCLmrZklupZmA9zguAtf3PGQxF
Mfs3m1/veU7amDBUWZhzLgQdfDj0TYp7At1W4s4hE71EclB2kuvyGhy96Ba55x97oGdsgoM9+ph5
sMXKTThdG5HcPKaeU75djQBI82jXyS7/5XkyN0j3yzlve5Lf63IXVxbb+k0Hxnu1xKLxIEy+Nthx
oN9BJzKNORNUxq6TsvtxDCQLZdq5VR7tY/Wai+BtkDnBTOMpuLxfxUy4E9O1yGT9yCEoKDUzlXVc
l7TVPIsjweyUfYs1wFb+76D4LvEFHyZVwYtBa/1jomkiOFHJ+lUbss4nJ94hr9MHoQ/MU0qs09BZ
jsUCIokkvDiGqAw9uOz9Ta6CoUXmT/rhFYHyk2s2i9opEPkwb8D44I6J7EJ7mCLm5ew0WWvwcjvm
MR0LuZB9ElMw5SI1qkHzQ9GjgZu8AwDtQBMztdKl6ACiqs/GAsaXB7BiR8ChkSfh8TXTq6aOJEbS
45b5qnFgLvZiUeg904F1daIz8iReiHfwq0pndrjtYzDrKO0e7GgO2ta4bI5spOs2Ay5cAA96zvzq
tfIwKKGEopbb3CRwZ4BZbt9Dg6mem4A4ARSi/FMXpG0iwtNbz/Kv0I28a4174j3gOcbyviy2tPah
n8u2oBCdV53dQbDQNcpO0Q7zfz0wo9qrPEgknVQFN/vuN/WuzvXcB3H7PdXuUZsjy1+8bGRcxmen
DbntSYOIvY6BfZ8tjaHRfIDmJ04t+wvejfbc19WmjQoZXNdrBOfGKVFBX6+ldE+k/WC2AIn3C5g4
uO42sonhckvwOt4T9jav0cg/Bybz5Z90yE0WRUjuNpvnXQjfNO9QCSrP8t9jHyhS8+JEixqKoa/J
HQlLlCQpYG3aZvl1BOv36RNzyrSP1ktP80DEmPjC4v/6vUPj+37S38LlSNHsMa3BHRSob8CS4QDJ
kJYsVxmweomc5D9UrX1sTeMOY3GycXdiTkFa5iUxwrKulXLh1SEEk4C6ho34ZHtwvHGYTJndsLtq
FWjRhbUCC7J54O7Xxx2M8ydTgoDpFyP7ta/L5Bhq6aHpH8GtwaPDLsadl0WMZ3u1Tz7pLHki3zAa
22WXfBcVoCmIhtbCUo83aIZszELfF2+e6+/Zt/dX7TocflhtGJPxxsrGzTDcE8/BGKNHBwlXdwRi
oPq9eVpsu5QwpdjYhlIJ3zgIGRjjcbTT2OdbhLKFj/yBqgFrZhDyrNaZW4AqUXkOJWS6O2HREiRQ
bGTcd4tz/n9VFR2+UKbaRbB+0ks4sGoGT8KVwMToqLSS+CJTjxNI2HPVksoKH1p+ahdGvQNNK62Z
qNRGQFM2YYGMZ1Em0pS4uHWLfwV3eNX393megnbGS0V8Bq0TomBt29hJz6+arrB/0vf5uP7UdwfN
C51MLbmxxNLz1s1p5+lGJTTF2O8smOhD7wu3Km6WhzdOCLpitHek07gQN40KlYvt08sQLeayHUbw
upEz4boaPVYVAJOLDw3lsJWHcuw3YBSAHaWcjN70mo9wSEJo2Z2WuuDr8F6+1TDaQIL+gGDznFKq
W8JGuLibWsykq7E2QowhYB8vdAdvG6PB6HsxkY6saOoV+LGY9v1H8qTLeaxSN1BHRqRghNnZZ7bM
dl3I758NEsfK3fGCbtMCNQ4QZLe/S89GgrAuSuM7/bLcn5TjZa2RigNxhHT2hEsTzTQK+d2vyLw6
YRBfIsqyxmqW6m4ADpHwQjwjBdBE7+4HEcjVi0GaqqNs9fUhloBI04n1tKorUpNkL9f9m11vjR8e
chk7E8YIJSOc87aRL/mGAxV47JV2cUcNzP/b7q9qPvVRsmKJoWuxOrQD92LlCmz4BBUYrQVrxLui
47+LHAQstXazMXG5cn7vENDoLMSJDilHY/y+87p1xJb4cp+21sz9gXeSVpVMmOuON2v8QNnjnXB5
mlrTgH29R/YKPKtUaRtfB6Oj+FrfzdAN9quT7HT4jyTuwJk25TvZtTeLPdFxIwErbUTD6dNp3+kH
L55gySZcgzmQlbyttBmuRuHwaLm1ttzFYASITbYx7F7CMmlOAyw8rIJEJhHLHAfAf3VwI3EbXsg+
fa6ZIG60nJNT/+XgggDdkrxM6CBZ+IV1GoSrosnp6yz7l1kY5kYEvpjZIdIyi2YVFOgQwhjUy4hu
mmvITmvEzRV5jKILBdvvZGyvWMSoGWfdVxwxhuyH+s966jlNUZaJn/QAdQSe3wjOkk8oHnehrBk2
nG+vtd9zdDjxK/h9kOEcb5oQ7dJZf7ZmDdRgWDfrvhXJ+TLairdXzQWvWD7hObTRJoUvBTNHt7dk
0AWVtBZdRG4yiTzRy4ld+6KxejiCElHCtn57GFGcYvn74EPTta7zEIHtyZQcwtKOGpcUVZuYFqo2
6urr4NcIib34oTBT2JBOLhdxTpzsKYHnJ551LisPqpaVZsMJ1GnyQ1DDLIfsR0wFuhsX0OGkXQ91
E5DyZinkEOhrZHXMnqcKAGr6tF4+mYMHx4rcK+yA+rKzTTQjvi5yQF9y3/GkF2wAJPDwjQZkpRp4
pho5bU+q8YD1ZPtMkytBop4cxZLwV7YPrjMX+UDbp4EJtdHSy2YXJb+MwqmuKtxVOrbn0eLBYtT9
zxyHnPWwtrFOEsXpppKHBacLnakzoMT+ZAvvQE4aEQlvGw+Iyu8zczb9Fg/txLgBUcsO1ZZijcDX
hz4GVfzfvB0MNvWtxOmkZTraaMhsbijx+TVrf/vKgQ6QAkHK2dAoTSSvVtyA1Y/4iHC+VcrOH3dP
m3mYvFpFyeHE9TmK/JOmr1zHKXiQqPS0FJlvd4Oh4qgS6+AYbCZihCtC9s1j25++sOnKdCn7NcJk
eoNQin2x5aal6d/xF75rE6fcQtfiU5BZ5HQaA1rTFe3U1Eo7d6jN9aZbreZWQa/fHI6gH1/eDE3Z
NqDJkOeERjVCmvq7mXvkDA+wR5VUtv1BKcIYx62AaJqgvnz0EIV1oNwmTOrfKFCfkdFL2naCVNgy
pQ5Jd1Yd5Fog3Z5lgC3KMcKCHZKsBBWwKnU6ivhMylNk/te2QTnIzofnZVGIDjiimX5qY7Mv04eO
2LuOE4hZTGtOhRlk8iQd0MC5AqpT5EyZ6SQ4HE8ewaDPSRPlwUJJr8gxzzHBgFOXqKynUGYX7aG4
u+cXVe3UGo235PI8Z+rtx1PYjJdIQQNz11xoVe5EbohjstGT1+/eKJEi3qHgYOuZzJL5vwzSGmy7
rxqwqPd+tSAmP4hSb9NHUnzjJgwF391o/uGjn543bm+uAf9oS3IS1za1yZGE0marTm2YElzBh4LD
H+xht4s7xEHMlaxUfHzyz2zIbRNENSzyNf7d/esS5iHFEyC2y/NX92DyDe+PuNjxNg5VE+ylJKp7
9AZN+sLp7jNY2IgSYOTQhuORWlnxTzyICK/Uq0NERzij6NSfaTKFZ4F8NtUyPxOA4qyoD1dXssX7
si2jBaYGAV3G7flED+AYX78cbGqwwf9a9iCK/Z2o8pbpEMvgbHETQCsfRjq1QbVJleLPaCRN4EVg
2qmomSX+/Nyc2upTlmw/9jDo25oirDniVpi3nCiJGnnEBte0rRBE/1MIrOTlJZSD+Y6XjcykY27a
8jzk4zjOsdtbjI3Ubdl2bK+0W4DLeRHzZKE0I0363So2iEtdaNjEzVjjeVW6iUNzvYrVHd9fbblY
Vx8YTxj8ANCxV0RHh1id2+QiXpFsGzNv6BUw0iq/2vnk4TZ4gkLOPlJQHeU+pKWpEje85iKdmL2Q
lCikMsdSVc9tKlgCQLzbEj/srS0EKeyLukZNCuYNIJbgWeQSYz1hsZGG3995VeAZY3wLs7CWlbMQ
ygw0c2cXg8hI/A0oIUz1zERc7/62HMTDDnGsG2WNuAQe8UhW5gFN0GQm/5rcgRuZAub3SX7mVroA
jazsDBhbMxFNRMMTJQZADLexsXVVIq9CbeBwDDDDd2UNJlKbI4wkCTJc4iiC0MIE92k/0jBX/8fm
bc5cJeFTeWe3DTyPqSKdu4I0Awo2BTI2Q0cDGt0jqnMMdVjXQjl0ZjSNpyp4UcJ4rvMiQEx2l2OO
qBT0N3A3A7/Yyeex6GY44+AE9PwRL+2FL05XvU3inJoy0QfeZjNtI335b2J3mvxqzw8NWPt8JlRb
g/xLyEbsY/B+2UnEYZqLNDu4//y0ejUzrq3XiFSiqcKF1nzcNam7akyMZOugV/OKUB8pISY0HxDl
bYFs10MWEWPEqWCWMKlESjagOnpgnmgHlyEnowe2cLhD9hIlrWv5lnIrRkYdRPow6WlzVzjJLn3V
r3ugypDFTBOM2ZByFSGueuJ557gK8mYdok1RFdwuC8u/Ox4VvutdcuDMrOvPdqOzrwLLUhNafRes
Jv5FkJsP5gQQzdCtCu7odcYHwLpR/Z7DJAMt6UyKj2mLGaf+9Wr4vY90Rj1e1ktsHez4iWKCy2T1
EnYfMLnFJiO6+TCtCIt8xLBsWsfBLnXwh7K8F05RpXr8k/UaTq9oXB/uy3nCbLNGgJs05xQwaxsr
OlnSzuPAY5+far7GciBT31u6R1Fm/ThTZOICpb/4zheRD9ruo7WetuNKizce920ISYQuKfmj31Bs
/V9YjzGChRhBEVxyvnIJXUawKlJyi5h6lUg5pX1vNhjF6G4UpgaH/pZvnnWlu7cN++y0BQmn/qWB
rYkZL5/fCJ5d+fI+xSy5AMWGou5lDHHR9RcqlLv9k/COjx695uLg05TdeRMGeT7JqyLCz8UgZsOv
mbGMr+XawipuefhRuPCx4FyW1SzFahJypoCZDJvo3uDhJccDABCp3sVNd5VY3ca0BqQeJGOOws+/
FU2vTjES6fQBVVTy1XLwJM0qHD+T82RUTaO5TRT03Hk3IYAiQzWYPjoK2YYeMKyFdSjkOwludllD
5N5s0G9p7784jhACarBnjjsEqGu2aoy3O7QfUhpQsxrkoNCGZbkBAeANsjPX7ouSrwGn5SRz5xSi
p6nHGYz8KOzHyv63VaBx0suYPyZEgpmjZaTgfmV9NBfSRDF8/wKhDSy9ZNGBAum/m624Bp6qI59n
fXap/f0Jmyi3cpgW4ppywgIm0DPANx4uRTVceHZ9J+BMGgw3PtPft30br1j+w44wbpifEXPZp5lw
RcAg3fPIcaXnLb9YPaPiVQe8dopqvp/ktaLiD3Ku9cGWgzsGFs3u3s9np435CxJN2Y0mvMkZDv19
a3VEaVlZf1OogoDRzyFzRQ/E59kk9OJkGNDe43n478l+7LsMPE/r3sxem7KRBgtyqT5XHQGvVM5Q
iY7eQxqXgmKwDAXbn6ajPjOXrTmoLO3J/uhS5ljXFBhLoNO1gCFJXdD4a+b8fPGUAZTVB578A3ru
hoqGDvuxgj7zG6jTUXo+DK59bvtzgqJLFvr1JI/DWDKrL3A4JlSKfQrAgBi8GaFAIgqkG3botk78
dhMqW5Et7D3EDA2fSwgGj9dlNLiEIaoxhWLu6V+K79QIRXI+JBAa+M2petXEal7M4bEey2+WNhY/
KatE4Cb3UpLEsQ8MCn493DxICSBTBCz5j3v23qRnsFlhOTIsDNbYNGZsEILNG2sDhpu2e2niABFZ
FjfZ9IFJmQizkb4yQ5RnCtXQlmNa2JXTuL0517d8nGwNLfRc2dBuV5BIzY4mFYmlcIR5mUGQiKT7
VQCwy56Qtabio9TfAq/lkLK3hC9bQoSIp1V2Zpf2P7PqSQm5AZwkn7udL7tSpCGhYzs8o3aPjd0Z
8vsCO56uBpxKyownVHsLM7v5ClnlUKtOCCzLJZdWIIoPNQRrIuBIpcimRNlHMHpyCC3N3xA5FhB/
O8v912U41H+jsmfL8nrKqru9CoiE972ugjozM6VYjWZHhWK3aiPk7KmVjAZ6FSko1Qx3LgG9dbK/
vmGw4+pkjmVzD52GKHztdrdHxwfgvAT3mvdYo8GAIAYxsVWKP7IE4kZNSFTJCPnUDNne5Y1JgGR9
VuAdebePU92qynu2M5EQLu7DWqRakK0/XUHxODj7JOD87hIz2iLADMGAGgGJc+13jTSCEIBxhneU
wXpe2gjIZMmvZL8XE0AINs1rfND1Z3IkJbg9/iIthTW697uUvBdRlZNBg9XM5gT617/KRGB3bKO2
LC3vb8pB3I0l4nj1mT83r74wyehoRre8g9FVKG25N/1GDzxYrxy3zAF1qY18Pv/X9OD8HoW0W4uE
1Q/GoYbtoihQTsu5Mo9OncOwNgHsD479jOSAinJWe4zBhJXNC5b2ndKsTc+KWSYIyGTIvM1m/gz3
umQu4VjP64tJnAVJAW8OAgs5YooPcZs1QJn6TfES1m3b78Xtbxp8wu2Zav+bi4FFPzHcrMaDh2IX
/EWPR65yJmU5dF3NN/x13Ov9odpHLQFGLYtOVymAnt3xII9d7vhwqRpNTUu7lWaTRkdwEjwWYYrf
CK6nGeaJTDv+CnnkCjWhpCPNiHoMx40y01Y69KMtez286vkmBvmULz5Lqyj6VpRdRTXdxRwMhNXJ
zkXm6aJ9nX0/f0BqG+qOUZzQv9IGvWijXxWmLQA0ME4qz7Dawx2A7/ZanuWK4l2SaiKKSl35xFIt
RcNQKqwV2RjFuGl8KU/BegNAj7WCp0mBLVXXHDp1CvKYuU4C/vddkvWZ26tQRT24BSt6Zjrloftp
Qzp8tlwNXsU2sg+gJG9+++N7iVTdeamByl6rIZjdbrBn3XSsuqO+0eW9rqyIelu4uKl57HMtDISk
qyOpNLGr9EhRH6r7+BcKTnQq7tksQ45/28R2rIJftiwzAb/HfVg2I7lzoT4b9/hMBDskLzmjhyRe
AtAc32mayEhF6WXwiYdslfiaXrSPAUenGq6Zo8KCA/DQ34U8JabY0rTn63yP84m/bAZ1n+zCdvy4
j83v44sNLCg71p6vIE15PmusB6mcnn7LkBr8HVwOAKyBp2iiimgVITEV4lZywNVhh1nBiH10vSGX
HDXZo2480K1TdJ14e2JpSWictIrPmzHHnXIOUuCw70oQNXKLk09EK65BID+dTn1CS//lvj6CUU/n
nJKVIQhKXn5mMvdAAwIteN7KZZzQRfP3SAgWe6lMwDd3+Lfo+Gdaqh69ZkaVlgSy7dIYrzlbJ8ol
nh5vHKAurGRUl9iEEKGX5+Sml//NXI1PgcVJ8G0PZ4POcmWKt/WBV4qnLT9i3lbMsMNbhcMOgAdz
qQckWzN1k7mNslOHTspSSzu2o9O3sKuR8/pZLfgW7xXbLEfE9lO2Edaaw1K10+1c90Kis6sdG+c0
1wl/ppplArv7fxmwqMnmWorQOVpXXBgEMfkWqbInyScq8Nefh7FPROtCb9OXeO/I9DzmkwkTxaEI
6LFxpFFL4WgW+GahsuerVe8lgWB5Vt1xuWJlA3QCWxHZ4nJ8K8Sx/uRxNDeFqa4S2p1AKPwA5RAr
DePFu1YaM+YPuwIDqgYVjfw6HgmCknu7SUMlSDKaq9PD0AVUGJx04vRh04gtr6H0SvfZQDR9wZPN
DJq8Bhb+CKnBbY1Vhsx5wzooeSw1eAYOVs7+KmVCYfJQHeazoe0s7uxj7QPMrFf6m/dmwESo02XS
mYavhIUlAtZwW5IaYKMh1Gyku4JUBfBaClQyoF8GJ/jl3YfkcbVcRFPhOH7e8Kgd1iBnGGSaNJFx
qZJTfvt8fZiYych/JfTWt37+E2/l9UQVJzdhhiDM+Lu89CKAhcwwFtWrw232j6c6vGVrHxA6dV8D
c5BPl3bc+GRvdUsHDSW46jqizu1KKz55OLTAQxV433h9IABBBd4of681lEheH4QfSZdIbHpKkjLu
BaLBQ12JpJ3amnuAq13sgzj/N/DEK3YfWIjJU1SzXH63DOhxImmhqK55y7aVN7PgGr1qFsdjzboW
wSNNYjNHJeb9HsEmvm/oPU/k6hDnH6z/wj+KOWA7O1U3W8FEE9FD59kiro5zItkbayatFpFizOWG
Jhd4j0ijrKz2uAjx/U1yIBLJB3U8h/VMTByqHwogyg5cypTeWsOtUGA755AvLXGVEyZUY96Ci7bw
mkNOcPLmZaDqy9zdOb1Chz+MGutxBXoAaBiDD08JpkjnVf5N0quczYtGF8prWNpAp0jrOgZVt6TS
mDlzwO2YgznZCeVBVOh0d9faY4tJ2r6xiF+ZcGbSlgjEGfFVGPNrZVCxZ56CiRBH7fbMzw8kbdnp
LtGOX0WjYgeQcA4gqU6yh8F+18oQ7iETs4RO3chImL8EPGUKtbjJvmj9P0+obeaGMuSeXR3bnI8P
1JRYLzemjhxh6cgG5mUZHrIvIDOOj+LoP+ObVIOSzKfiUASXZ4lYFyVrCTXPCkE3SFdvJ95Qpcc0
MyTYV5z0UD37J05rZwiOo7pQKxcEYxXLLV6DtUZCK7hhpYyNdthMvf/US1sBY8g38ewR6QZSTHOP
6BUkAKo4EpdO6Cm+7MnZQNJz86Fyd/W6H03ySYSxJArcVeoDZEzcWPNxJcGlmqdTuMpPbZvov4Y/
ZnC4aMbzu+Cw93z9shmCy4x21wWD24HQyqCBjH94zss3Um8RdCyl5MtpLbgG0GtvPxhZag3nDZME
pO5uPPnnJhFLmYusSsbcTV048DjpI/m84c8eJMvGrYZUFXhDRH/j5t2UKGGXErkdlQcpy7xlS3QL
6aUVUvU0VNnX21OCdw2TPgdDJOgfG6bA1sNDSc/PYFC8kW7GIhLNlwprVS+n4mkpmVcDQb0hkN1g
o/VhbIMb0/km5Op/JlSUFjJGDpXt67EOELZhoOs2vBcQHFRSM3SN5Ax+z5QfaTZpQIcJHMRYyLHw
+7W2gh0VhGHcCxtDH0Exo8vFlGG27RUvg4/7Da0c+PbEVdXG9VOJzwyP4U6SIjqOzeMIuiUkL/0y
c4Bt32K/dEIJESYR/jvJsrU9kz3tNLs7Lnmcs+GggNLecVHOuDmvHvQxoALG5EdpPk4XdCa2W6Jj
PCFixDL1qI0k2FOfHNZDZDQbZUgjKyoaWjqYkmGEg2p9K2d8qixLSkCEKtlwYa3QcoT1oZ50qesV
dQMX6yNSVDysdB9R7A+zIaIojfUAxUzkxj8wmNgEiNMGjqbGzDmxGcEyxMopje3jiAzUBUlbZYn3
wULvenptjV3seAAld2dCajsv/JR6Th1zvt0GYU4MfJVTFokrW4JuyBDR9Tp8gOFNt21z/B26v0A0
JEnQ2/pyuWERSuoPn2gnJc6bNstEiaRag421Or1eMRB/EzVXyNpl5/apQhfaWymH08BR75tI5pdQ
LVxtk5tJKrRTxwnkUBr++BkDZ/hKKqhrH2NOxrL9jJfNWDIVFkNAyUpRYgvDVgPuUtd+EQfIYJuJ
KF3o84XKfId459FIxhtKSQUEghsjWN6QPrzXTV616KjiVjxedwQ+4D0KXfNRC3MU361IsdfXs7xB
IhEC/4VjFwLXON3rceUsDU5xti9/IgplRIFA00zTOBFrz1oExahy0cC3RuG7vXI75Aq3gUecDlO8
wx/Oyvn2uZVNoAXb48BrcAbXeB1fwFnOSdUseDOoMfOY+DePubgjRd2OE9tXY9FggPLRVDo9+tRd
mhzV/ElIEb8X9Ve7OKSg7RMjME4Xp/pL8k1BOdQLBhgEaRox1sn39L/GnrMDssC7A39CpNz9LvhX
bi6rdDMljMNaEAn3dMjj25gpjkRrYnhzPHParwzmHN5d2WOfZ6G3Jrg9u0KgYFu0Oi7ghBWlZA19
tWKXNI654Lpvyd87z1bvYHrR1UWztvD792vxppYcsCJp4ZXm1OU9obu8fMViAaL4I7pZacgFT1YR
qeePTzmvhWXIMxym8IjCt9sNiiwYri2IbdZcDZIMYOF6Zq70MdONcOx967QpMPVDqdoAXHtqJ1lh
EUISoF5L/60HSvNB3bPkizTyFqxyIW00NB/NyemxCAGVl8bR7WbjEm1+ic9YoFyJZ+L3zvq1HbaA
vtS+dKdkejFICBBl5dqYAfNo3WNmDr1PefMrqYdfxwyctAZ4c3XmHUErsd7hmn1sV2cgOYvIsL7b
JgVk+dYySqLEPzNEM68ZtGTYPFpdgtzUBW5s75m/SRIHaEw1ymLF7I7EGyvJWM4WdtMjo4/eYyZb
6dd5vCpwuxWmz/0jaeaF2/wRM7mwQ/WuPfpjAorLv41Q2+SX2h33eU2t0IwlF5LnZ01WHRMQHbM5
lPAPMylxcD0YN3dt3X6rxikQ/uMas8hQcKhkyYx20vsnuGwm5aa9CFJehIUxrIeVCYxJsqaoSQHv
s9bL5TDXzgdZizct4WKtUHv5I8DwtnDesrFGPLicOOz/oG3ZculoUC9V2YlDLXJZhehLZTNHq5oA
oS0GYAAjozrQxvbP221SQQuE2MTRqHXFCwSSKyJ6kulUl3oUBy18ss5vVPnnsGz26JYH2baPTC9O
DIYAUqLsDktOfXcAp5tbKoxUMTInZhpt0XJkh1t/XMuy7liRY3siQbQrNWV2BOjyGHKM9eLJ8aLu
4WlOTp70H47Ci/GkxNzQ+nDBNuQLW+ioEH0XGVusp76XTCj7jEj3RBaPpgKyMFH0r0ex2D6H/wzW
hllRNTEQDhr7NygXYJZqEzYL/wczBJzNHfDfVuRWnnPMCUD1YjpN+/yqFpblnepYtuZ9pJclBJ7K
8/YbifI41MJPrElzAMRRin+Oyho4ptrj1lxxJRBVreCp/JkEfGMhDX1eJk8QdUF3eC74YBJXXowT
f1WfdOnhvTbHfNsc4cCI5avluLf/FVDCf9Dws2/iu7sXiHs42OfAn82doLBJlyyTpzRct+3q3g1J
s5qHd3RcxYVZA2OmIdsMWhPuIxz0B8C38ALPIlT+HnBf1xvStmfUNDjOwEW2ZNxNqd4a2XSH3ElB
b3tuy1Tw0fmeAxvdlHAsVsbUypUZJouZroz2+OwDw5wfWVpBZzlpoPgwgMUcq95s88jgZEmewP0e
wpvPYGK8WSDF4kYFZKivBF7tHy44gSW2svgVJzd6vw3p+FmPnpabGpwiHfinINS9J4LZ9GOKA6DN
QHHjciKEjp7kiYADKx7EwIK9qOQnj/x7vfQELxPRTx94OvAbJm597CTt0EJRLn/X1/KnAukW7K26
EX2DoxxzeTY7iqgQzY4RVLKC+K/TZ1nr20cqiNffUMs8jqINmARPGA6qfN8kdGtqaHXTSbNjIsvD
yJeCDQNukos0Cd6484G1AI5YjMzd9gT2z4tr/uih//nsEtfpYruqpLbeLk6+L9y1h19QceGMNf/O
dvnoTfRmGhd4P9R75voKmQ/m4bWAUOHPArrnWJCNUMDhJ4ot9Z3e4DyZ2RSIPr3Ba3BbrBpK3sgK
TzRvd9Nin5SaiGArP8qFXQkwxkDPcJJlXfsQMVhIJ3UXpUyzCFIikJ0srrcU5Ii62VVRebCrLSf1
oZ9wPbFbtKDp9JhfmbJ7IjOQlZdWnyBI+EhH7PqgIDgcWxyuMd5Cn3oGsh+GosHu+EmLjXW7D+sL
naTfW/Q2TgVwATCHxlis9V4ufxTYRUxJgp+js0mUeedehAafpRLGxu5B6wKg5DTdGXxHsJTLY9nC
/gXk0CNzYiu6Hs0Kh5bve++qIrV5Ped7LLJTChLdg3hzlCNbORih4FbiZl4iM9NlXXp6oltexp02
lqigcNbGQtqppT2yY+lgZDzUoyJQBjhFfWUXDPVdxkzawz+tq4BquWDEISRMiedpR8ODZh1k8CVU
xL+ebOnsczMFQLqrH2nWkRn+REDQ7uJPh7TFsUSIJIrKNJZ2jLErZa4m7itFbrulcdaosnKwACTB
uRKPjK/FJ+HROYTCz5dRNl7BEAGYKQc9aLNZg2AehMJxnFz+B2UzBEnF9kYqFsjo2EHzphgWs88T
uBveXRSmjxHRwakhAgGFAuGuhOi+u2ihySE2nnk3AG8AzUocUy154JJnwoHrqywctFeWYxkERl9l
ndc12c+QIOVngqM3hekcmZ3jbJR0yZlV19YoVE+3ZRpx79kHrb2OjsxRdSNcNHmx7xhDB/G7WV6u
9JKz/fwK7ABLxS/pOT3VUZnaaPK3P2AWCovug+r+aA5KaZLpuwFMqFr77Qe63KHV76/kXg3dwrTG
BXjs5DeLPLZ3Y7jpaw47L9DasoXA2NUBtM97lUHry8GF2cKNIMSD1lqRb6NgmzmjskMc6BqLLub+
sfKimXvksjSKbPN6efaQPYRivqBnnqZVDfk917ul5wHHz7flysNEF1yl5BCWZQN5AjXC7bxRcI0u
nCc9AISNFhhr8Z7GeP958AiOp166OS+0IYyyqh3zc0p7MOl12sbvl78NZG8+zOdo5HI/Xey/jQJX
8MThOKTQ9Pqwbjw3G/VCwUK2YXH5bIWB9YL72bgngJYX/cutbNDp0fX0YB4zX7Au6pdIPlUs/XCZ
Ui76lBeq2sHMRfcDdUA8UukdWuEEYyyVGhmz39yX0GeFMkfzFYBk300TPpZxegYlIebo+Xpq2My2
fB6H+IRzUHT8+mN8Iuq01CVcA6wLhwpuXSDBx5iNXfQrDflKIFDDNG/bowHoi9YGq0S4+atT179R
ZGt6xD+b265hkYsP4Rq00hqyVXmP0G/23IAfzfmvp3uofhtS85dYQuV8jIOvPqZnkEUF6ZrPa9pX
IXyhCB3/O43qF635++YiWHn3Kh0Sw88lBaEt2Iy1942vXJyQDmikvbhl8f24bGOxM7Va7T8Pczf+
ABNqAwkkU4nbJ3LEAiMmQvuiYLR6k/dGDVo9ngGPhcAhM++QxknO0FZmOr5IO809d3kWIxEGnI2f
uS1y6TWQPUpJMAmLRjnPO0Z2PbWbG4mLLXU36VOgwf4fZA94LnEj+p2m+RtDdD6VyeaH5peLDxBu
w3nlFFzqaTB0ZSfN/EXoqLANlX0AasbDaS0AXCEnFTHj/Gpaa4BGWUv4TcVOViyZETX68BO0hZHh
DCu/QKs98yWIeLTWLky4GkogPB6yM+j7cWxZi4yzSMkuVeVOYT2pLHeRP3WSS68+GuprPtuYIeB8
kVD7iIXBe65VhJ6Mwt4baD97VxbGJ6Ge7l7WOnLu/9qeDpDfWdZgRIszI8oNwwgtuDIzm/dZM31a
3Nlw+ju+Ls+EuOZrqQBqFWDyGMUZ6mX77jA8W5ba1bPA91JF/8CLl02r5HPwjLbv6ty/RC03tarh
UX8gTsYXFLTD2x4geBcfuLDAkLCXHuMLymOz20pdqQYnsFG0Ow/Nc1i4z7mrMCjEkWWxG5UOxiGQ
7X+5PqGZ8lzpkXiDY5G9YEbhDfaMb2sVEhZsCNa1xHAL4It1wRnQ4c32ovVYqT7FjeQvW9bMPnWx
TMDbKVdXsFpUv2fltUBUGNwyhSNJ43gWjVrKZvezi9SPo2KAlx6xML3diAsG4QbwtXcx4aSIDZ7I
bfEbasS+isRJQge/nsPncsU1awWfNGIwCTuEZX8P0oxqS7k0w2xeTE3OeX9aefWbeQCMrlCKujfc
4TNJHbw4XrW/Aq+36mKmedjHbs0oXHN+hLx4UPCZWDTtZf0Rr7wxdjSQsTJXgiWH/rSKsySn0xy7
zUT591hRW4yjrBvVIAhRiTCgKlcj0qSQa4TlI/padygx9or7eFExYDe5tHqNvh23dpRTOrBjXWEP
vNsKG+iqmvedpWaC7D8De2VHsSCDZolz11vMcEefFNvnkxg0lXGbIrsRwchF1WR2vC5ocfikD6Rm
jzqTAQUZZ0gQaNMzmQJc9BoBP/dYw4nVPJvbqU6FPIYSDubqYKCoPbqnZ+SGwtS7E6JMNCRXRrQ2
DRwYMKfEcE0909PwKT3kRw+WctRMs91UuEos7ZF9Efmj/E7r+Vsly8gRAinptaSmZfdnNbmJReTE
0/3qDihJSltuTfwZNjN4hosaLXKugLIG+uU8ZPSlYjUy2iSAPR8yockbJa59WzxQs1I05ZZ98KzO
z6w4ewkyt6Me9fGNQ9gXl8+jqLzo/reaBKM1VP1eAdqwYhpMwvcf6eYcVU3pVv2ilwzoDrDduCa+
G0ugB+D/d0fgGjwYhaoI1xhK7VjSDde/WQ7aPp7xNOyBsEVznhRXx7Gx0Lt1R9joeWkGo0ex5H5e
mqk/J1keIf6o2JKHtZbRNYZEWqYxTNhC4rs/QG5ez5c8Gsh5yu9sgIWLNJRSEK33H8CNGdyo5FCW
JimpO+Lj/NbHd2yaHyaBfaxydT2InVkS6245jFYDCWARme3KT7WavWBa8mRga7gXlbilVF4jK/fB
WMiTZ3v0oYB2boZcDmj2jyOtvbyjDo3idGVSaRz4OqA5p+HnexzsEM1F0B1MpobP0hvcT5NE54ft
hWQ3EexQL3w0KirdES6pkta1vh2Kg/2MN3JqcAM1h8WYv1Y373bHe4AzsclKi4+z2DpdsLjh6K/K
OQH9UL3DXRK7Q7LPgihKr0i/MQ2iTybu5rLpKr1QxlBOueJ8oN+Is7efuWfHnVdkHk2PPFHBSVQC
+1RrXSveGHw+aWkeXsSC/s1TQkCoJAMGKnzdP3dmzbd4m4b6LC46Uqtw+G8sobcz2LuXlGNYOeSy
ssKPrJFSd6+svh7Nc04BPryEM4GcwLNatTif049rCgsQJ4uIDnA0n3PFumpEn2IKBTa7281E1hiQ
cOA+2xJuNS4UFM9YCdG4bcNM3gd8LXO+Sit/NpUe8pxA6OeKZoLhPeRDNtDOSISZvHIhJ5Ob6Mkt
goQx1p/FQkbRElBicVImePCLRNo5f3Ym3ATIt81yChrax3O460hebP3uE+VnVrJuG2yWH0Y2eZkE
Uyt/s2iW6QFdUxza6Nza4onQLQ+OIJpyL+SkR1kPnhcfWiVw9Nhk18NkA74WII5rXFkombVPSpdj
tvpEsSBdn23Faf2WmU6dYoqPf3spnm3/KK/MToq1JKr/hy43FItmIOTrsoYN19YI22eHdh54VQCO
mBt/TkYdzf7VsavrbttAfQul49LQNzJRVoNHXA4YmMHNOc66zJ1YyGzd0oAvm6Kic7rFbFIu1ta+
d11+igLCSOl9tfPb2fVaPrbyHRF+1ezphUTY8JfraLVXRkdaWgT7kFS9NqxluANtyPepxBremyT8
cjet67s/4gvoS3Fut2jMjWXqmu0Zhkf2UMsKfVHce/LGJ+kZsiYSYPdLtOgfSisPdm74gO/oVvU3
6aRH0A7smMX5meFNSQGImNriLirRcmJA+jQmCVZZGh4/yThoderh69GC9x4XMKNo68mJYj7jX44Q
uW7bTaXClCmph2tdatolItNJOJ4sZjR5CkfKKrU3SOxqr4qcqrX/l6yJ+LKqyz6mmFgb7iDX+lRT
FhUiGcykPAT78oZraeaAYDawiOQd5O8LE+qpVojZNae8iH1u+jOYaUMqVp5zA0/j87RNnqbKEIrD
EbIBw+hUeTBirNqoVgH7MOQ8cVGhEqb4RDd2AfllXHgR0RBPkoXa2bL6sDsDeYvlZq7pteU7E9Dv
WYAWO2MJN/mtGSWKJwe+I7QWJ9/F3nytDppBZdbNgCpqX6B9tZHzqezepJfRyGy34OT5+CtoiQgk
dREtZSf9OI6jp3ztwkYPKw3zq0XPAH1MTCTiVR93XM4cqPIgIYscN/lJ/pWorHxaLYvcZqmw8tAN
v2oaPt9X7GLK+rLpH43X6cT/6wIzDO+nvi7NXLTujq3dtd9Q7Ut7yq+ebqdeU93hjK8+H9GlStlg
S4wvF41tcifzGeYVoRHRTE+TfzvRK4SiOJ+bZHtm+qxNcoNWyJu0ROY9QNktINqWHMi8GpQA9Cpz
U0t1ufhJX+8Pqem7tK6oHHaszWTfGAe3rDkX1CQLHgnO951ZZkMddd9rna/F9cWRqDG4iLXA0/bT
2ZuqZ8rycTaqARPenOkkYbNlzTqfb8jLYbf+6bY33/qNtt3fVgZxAEd5j4Z/5hq3IGyvve5boHHw
HAYUjlwCQA1s6OTkwrTkwySFwWc4FOqoqcEuh9nitUwUXxU5MEkMOq+AA+4bUTW5kRmtiCxdhHyR
VNjxYlPfMy0YHlJKdrbxNQmHdz2HK4W6SZ7okf74ob3W2oDaM21rbSv6Yh7Pp+hAyk5jE30cMTIZ
dmnZwbaivndXNpbit4TMWYOoyNG4VQsOSe9gLxWbvM2xAokx1zE5yViSJN7x0OcSZeynwMkeGUzO
djU6pvNJZFFIM4Kd6sK8/hWG3RYME+7kLIdMovC6rlHPRzCWLNSfeR6AWHI/dgTsmRCrNk94VHho
7f6MvOry9wtffGzyalGWurpfAyOKqCGuI7MPPabeVxK2fs2w+GaUk/F/tx3X6DLTr2O5mNRMtGUs
4VaFviwCrQyMiS1ee6JO8RKlZKKpSdOpRIX2Y3O9ki0vJmRGpPIEXTzRNSeu17rJLbPqyD8zCs94
s6fusCAAe+YgZdJ9JQDspyFq3hSrhq/0PTL8ztTLf9Je9R9OBpHtYmWcEKv3J3Y8vxHCr4jKl4WZ
1aTf5U9L9tSdNU4R7NUp8AEiLXAY61jN1X2t2ncmUpXywJ9qFsKo4v1p3LWdD9ftlMc4r0xZunNG
qqD8EdlLWxPSUoAz+e4YYd1dBuWC0s20LovveqDDYc0RgjBtUzVA0XA8QMxpYCSSrZmYpdGOpToa
UYCF6ZyIgPnGIVNZWSaZT1+SJgXGEE7wdWh2fA7D3FAYKEkRYU9h6pd81kIxiMfrz25v3tGMpZaE
fVbDaxX8Z6Dfax+DTneIV/p5nbK0+zeL2VyUqYiGVJBPxW5jTbUAFrRsl0XdtJbxautpsY9312lK
kFAHbml+EWDzm5/fJ+sqbIbvi5xaI5UCzCfMlnxNxwNm0hf0ppbzwJIm5oS9okisav31QKkLRR1G
WCdbOcAePpVZNJRvk7eDjRw33CyrX5NpmYPJFONgu9cu0yHd9gXHJU//lx6XEyWBIhQk7UK7+za+
e9ajlfWsr5g5YavBamck3UPQ2W3Rwxs8wgjJCvTAwy2ehFTK3Q7bhfHDxOeh+dgIRkMi0s85mmTw
mA8SEBJx9ePXN6Dg9iYETa26XGODWvmW9q/EN+Ogjn8Wsoquz6wITduXU3YSu5FcnutqMrwiz+AL
KrkiKiUG0EGyaqbvdVyxWGlDhUedGeUAPsAD+5Cb6yvI+MZU3jfDcLCY95t0IdfEjvxss9SoHTrm
2nyR0xTRXE17asnLNwA+oYi9LtgP7JUpNlrvNQqzg9Y4cn1ws4kl19bCiqg+KH8oYwZzZsdp5eOP
8O/ogTediA7vKvMMmdcgLkWV33wNhDja0OOq3weFOzR2Qg0wvZsvxG/pDt5r2n18Z9tp69buSPHL
mdSLhQLDXjGj+4m73RgI7pP67zOy6MLPY/3G+/ml55mZH7AHqNYnCoTWd/ONhQl7vFRBlmgy3gIZ
RcWx8BwxT9dhzd9yqyMq23LAJgCyf5npnnjRD0j5LAUbdbt14tk+DZ4zw7GVYbs2L8Pl3juyiIZ9
Xfn82zXFDOKW51xomjPoYiY0UIFnXhq22+LA4hjBxrorxsF8GnqpqABrgzJcruTI7ddrPnMLMv7z
IvuIxMT+Lp0HqMirS8bGzgQfWMXTRBIC0COBaH+rE53P6K4w2xaJePLZfzU1KAgLIODsle1jMx17
fWRHCBUtccIccrX8V620ThJqhoSM4fR5oJr0L48/0MMG9lUzbGt4rsvrpyhaGx2Xy363KKMSLLEM
AqixFnHNgqXzW7fbTVL6q/SgfKnxUr4/7d06iCrk0R0L9d2vsbCEQfkL8BGFae8vB0ieE/0N7AU5
0EIUBSMlur8c/ADS+MvQGRBqp9I5zo5t1wvFnf5CWD+iZvgUmNfK6WWuMp6NWL/uWoAOi4eCnhro
d2Qp3iXCqwTsPKuV/iOg7IThh0VIfy/bF3R+z8u61n57FEy5aGmDCF4MWSlD6W03kEnLNrbRg6dM
Uyw+CnfpplUkq3w5fPnRDVOBZwSihKrzX0NZfcicc9ooYnUpCiB7pUVyUYIj7pKCW+1cuyvF/82g
Feccd4itWpBc5k/O7KQ/z2mq8GyxMt/qVmzhYhMi+fPUAkA2OcV2ngxv4uwV8s6q2U5GwipEVAZy
u9Y5Z3SiHyUxOKCE54WdPG3xvTQT4T3gwYvSOKo9Lzw+s61qyUWBwki/+6vPTU5OAZYg12UTJhVU
3ly/zSyRn1/LeJX+fhc+9r3Yzz196exhTeQGYEp3FnMdZcVz+PKf0QoRarWbqL4PHCCsElB57/or
6XJhkkzBZ+1PUAuYlEnVjPCNjsl/G3+nnZmj+REbyFxyEgfntoWKBdH5FUlr+lgcCqte01WNbIwt
6QT5sHAxV9apfo6l2OZBsjcHUhuopoQmWXNXUD1dXhOwC29qZrP4RY3swnKh648OlznJBfHLEyWr
VL5AugA6+Zlyd6HjOokKK4QgKqG5yxc12qOi+oC0IpMg0BAYQMqc18P/O2ou2zcWi5J54CZU3I0c
saJccRd8RjoKqpcgGYZ/pbUTDC71Wz3kGp1CttfUajmUyj9uYJmDz7FIUoXIxy9U38Tp9PxhNs9e
VSDwUBdMv431aGnRRPdx+AGisdpdUa6sKhkIzLCxMC8sAnwe+uQ/F1hOO1TuFZfbgJkTbfKeweuP
o4u7FJlUxzdSTU6+tmaHHIwwPe7AnS2vldjRFLVsJWUS0sBt8jVxUvJad4v4TnpWEdIsHnjF1SAu
YCzEJvwfn7WYV1SMTU5qwClCy/oZUqYPKswpYKm94YufnHBX9t7VhUcH1tM6AQoNmb+gXh1/rTrp
amIxm2hf/B3oqJLR7jJ3Yh4ZFXtM4wRZ3O9XFFKedqq2wXa6l8mVhk2kM/lLK0MofaTZFLEv5Amg
6wtzycQf9dPcOQ7IDsezHuV4M2u2iL3KFQMN6H9ajf/G+cSqeGlcqjt+QsEp+AgUdl9v4MIKvu4g
wmcJWmGlgkRILB88fuRFMio8z7miCZAzA+e78EqrL5G8edKZhz5UzrheXlD7cEAsVLkcmrgnQncO
bZJm9xTyf0SXWOtKr8b0Psbu9BR3ml0joUZLhgxy26hB5KOFGHPXH2lwCEsEr6PIB5MQ6zW4LM/f
14HTCIukObg3xREbmS100wlkX+E40mMJPG2lRm9vzg2OdEhXuVHT1Jnq7EX/i1ZFKtFQBa+3NpS1
dT9EXQnblPKuFYeQwEZ56D8rKspRtLgNUk2ZNlUKqWEGBcG90OuXzN42kpoImxbjnfBZR3DCJOl3
0IY7vRDtxZk/0TEELETXDj034OVNJQWzrmChyyjU6wO3Sgq2tI6Evp3l95vst3uFMl68IDMHv2fU
fvgZLwxHQVN6oEib1Jj/XcwxkzmAv938lkrwzdVA/ZvPYXhE2Eg2bnbEVnaMRfzGlOS+0RSKVEB1
kTiESyYxRYqeWgC6rNUlxf/0QwXVIzUQxN/wPxdMKW/yhnRGZWHhkhP1Igtk8O93RNiEbFLGFdbx
6hvcoN51R2GU8PH9qZtGqMlXENxgEbqLbBMs0SGavSiicVqgPObHO96tkTn4Qq+DKQI9IZ5i7XPb
p9B+9Gy8w3Kb9FPRwGL0AxyLvA6KIRS8fK4lg2+8mf+po7vGcXLxvaga9gXW19VBFVilVAtsvZpJ
ecB1ToakApXoGSOp9WrmggNWrW/nXjILj2vLGx6aqS89O0lNbXeRnZnUa0C5onDVDoIn/xmnE4ed
Qf/M9EPgiDq5geaHXVFiYTmZY26UdGB0zVluSK3YGz9D45kQxWKaI5V302IsBnwRYutss6o9iLVq
3R6xPBmZI/ATVryf4fwJU+alaYMet1CBc6eJuTSvfl/ZwF12Hco0QtCRDLGKUfs4W+Ix84xwQDpv
CVhq0ugvKq807S5F2kmiemPKEQoWP8lO9NE5pN6n8GZYfn18ZRFFVbr7oGa9NePeLvJo0Uoty7ao
+WkMXShYHA5A/LoXrbjtdJ6aTRzQaWGeZ2YTDVIIho5Vb1sQRF4UNPvjjwZ8SH14u1Eny6KuexMB
AMdWvYUkk7kj/uvUKMuJcb28tfecHYhe1ybOMyvF4Czo9NPhao+fuKJArBBkLeJvvW1sD1IGUY6/
XOn+R3tVt9IVbIbD084kcrd6doiGied5eFJAwENGM6MsXJIZzkfN7QdFeoHNFOEe177gkiHXFMhB
b7yZWE4evys1iKetbOPwQUC+oSg+po0Bt74nyX6XyspExYjzXve+FLSJsu3x7hBINt9mB8lBFCLq
JhhGbrwA/TD92rwGMBJskDFOeyGOSUBBzbLFNCbIVGPeJIL1Df1d/9p8d6kt6hn9A8feStjnQIVX
0+/jKSS/hMH7FPRqz2ZPeo6EML2dC9O1e2PWIxYVfbOfGQfKO9ainrcdphPD3geDXrzS//X+0iVU
zIXszLQuhDQ3dYufYi9swUORebrsFISV05JjaaQv+JIrKRKRfQ0aE5tQ++ohLNrMEBQxijw1JVpy
9vDus/0DK1AUuFAFt5IdcEZfI1BM+WT0NCQ4M1boWUxvFptALDDa6y0qzD55XBLnS+kQyaVY47k+
iwXGkgKucNJU1liL+jceSgEMyg/DpzHw5pwllS3Vxf/Zcp9DQfVDpeRnxKuNV8HyP+twr76uTpV1
vVSAf6CEDEyurmcAgYIuS6FFVcgO0XEDD5AHPxd9xEp/Yemon4fkQicrCOq9R+QGyOKJBCM7OFhE
uiJjv6fo7iXLJJ+7OQhvQS4L057Ym7tUl8bPjH91cD/LbPd9r2iUD7dGuikYJYEdWn6onVrNhJej
sgOVrEjdvLoAIRHN3/eGx95bz5Kmtrymoa3+Iv66VEIYqT15u/kkym6/GYX3+GJ0dwsX5jnSFzDk
36xk/ggnYSzXzO6YJTn5e9v9iGsDkhITyO3+SNevoZe6o5U550G/yAn3+rXWo798beCCmYB3igwj
OTxnpmPdn6TfydAedCE9tYENiwrmRmTlxF75AxZVQPkRvLF0WK198E0E4BTI9pbl6vAZSl02AcYt
44wYt/LYavQgxo88enJ09UtI2bHAbvPTElfdr4uiKY4098xYCedO3abWaSmY/ikpXF1J8AEBzROS
GdlBPhx8VM7QeLjtQUAUgfo03Wt1NJjwCpOdNHFguVytFn5rMBq4JORsm1I4VDICEmr5lWILTM6s
VJbILEf0r4P9ZYXRKFJLHkLIflTFCdtdhpob4e2OOX4xt8QgJnmpejVzOe2qC0PFoH/QHza8qpWd
M6jN8KDrRK7HQkZy2Z90IqjhQDdkeao3ZufqEtiNkUpKDwRxx+nqEBaNVGE2VR+gmdDCBc48Fpsu
i0eJCl85NwBcrcpHGvUr3QoUg3U9DA/BTjuhSGpnx7wpEvfwo6DhOQRn8m8mCJUa6opYPcDlzlGF
hF3OTwGAUTrpDXJwPcSpYOlg0AbPzbQrdyRPZHeUA2gYR51htgNqLWtVCtLgYECUbbR0GeweMLJT
i3KOPbnJYalLR3B+WsBsDfWVyUbhPsG8BcEHkqpXj1hyL7IJMcmDTD4L0iGADN+JYUMYuF9eyzSm
/PD9bfF+1Adv/v9eenoOTDOefAW5hTQfdT5j0VWEXjqU3VyDlY0c0fsqo6rEJQCVcw/40prYMpQ/
cc3yCs8ygc+NEdnnP6qukMwvMLzRC2qN1oyMo8JRRFizjnGX01ogj/TE0MP1K3fpl6r2CwSx6Vbb
qEoe8LJXmP/GIzLMUOkoNz1pYkfBLHAwVl/v54jSgHpnFlDX0x6lh+L5lIJbFiNo/yF/4kLOVmZf
iRQE6VDwe1GDaG6UTqinn6CKgWDeE3cCJ+4gxQmX0O5AVl93JgY8qCnSyPVtXgrfjBcVbX7QM1EH
Dsz+eGFciLGDbF1ruf+sGkOYwGG0zqfmhGeI3vFoXQaRvCm4/msjuxPA5csuwONAEBD/rPeR9rYa
7DhXWh90MkxHRSktUVU1+7cWjoSnnjjNx/owOR8HLEFYyq6rHgDGUi335mTM5imQCxOwbYWV4DEp
kI+4UiJvBrSlvTX3Fm5I7Y8ydP6WUgZcS+5Dh3JxNcMyo0bxtDbrRj7aKTUKrgBB0BTeXsBMb3/k
JcuQOQoWN2mSknEOSo6rGWaJrQXGd+XFh/1AKjrk/TOFzlNn5rk5IDmmi5blLDC5b+yyUbyRGd0k
KMfC+/bu17nJUW9Lox40DKjFL61noTJWbdv/FE7KvDj50rX9MVBAvivrtTfDqQhFbnEoM6uqivZj
GO5ON6deM7lDXzFL4HXe2SWuFQEI64kO/mzZFVSMnKwc5sQ3OMCZrHSxoiJujwaBNkmg37ZKXPID
VzedF0A7cE0y6AszLAwDt7+JJZ2sWsTFi8tiJYyFYfyF4xT3gEyINISCFAqqIg+C3eKlz3oQfNDi
XBhPYQBaRzgaDtzMJtEsqf7LKBE1GndG1KBehhSwrsjhJSI7x0IxtqZKR0InoF03QsLCKfuEgyWg
//DeSCmkwEq/frjAhXXs2WlhVIEiqBlArb55pupHPvI6QDkM3imDX9M2TlyhymZBTYPwECpPTkob
mHvKqlhHAviBW6aewyskwVr70WakuTzORrAV4Wgf2EkfXu90Sy65CqF2R+yjRI2JQxiF9KQLdWtO
pfAFjvOXR/y6tVz18pMyxudaSU/g+0AbxOhtGyHEn4kwM8x0P4D0g6kUt4sVCbtT+Z7O05sqBsV+
elDg/+OotXjVk3bSaWyFyXyUb1/BdjXFMAFPiSDN/BncHLC3hMLlyLdZy94YJqS5D9bBgPtMUHMi
qcAmlq/2uatytMBxlvdwS9++k5Bblue8BEyeeKgqf4f+90HOIwWo6l+d1gbGNWAwLLlmpUfwvLnw
m6cEKDYt0b4TNt/5LTOm1ribztjB/cDb3DCNmqfvKreuYSsMU0gNtDeWLnz9YN1OeRcbRjnDf1Us
Y8hkWhzNXI19ekYsRDY3dZV8+oFvs4LbD8o8fMZdA8HY83y9KyFdHI4vVefO+P4MXrQM8OKVJGos
3uQT1RchePe/sCe4veGPOwBxgAeETGbF3h+PrLcimp03A+HVgnMEzBNpQ1HnMuVtIRQBlLsoxGOe
HZQwysJcxcOwWaRfxnno2S0ucAP5LYee57JpccgpUGtX9bdmaFB5DxAwgTrovZdHuabdBIe58EPe
Mzc4KT49ygkQs+5Q8cIxMjRCR2w+JhcDi+DLtcFfMlY0UbKfSoPq1AAOhhBFkCP8BZMC9nkRPBPS
1geI00kHl5+DC7h8VfprpcmkU9mvquyed5qEmdHr3nkhXGWKqbSkGhBnTtHfgCQE27h1BuF52P/6
ZbqbAEsUM8QZ7HJqMAprn7g2jGlMiEI6oMnkGQqKCrWoS2SQdK1lhw2LVH6UyXctzJ2bcbiBvpLr
maX2Jw5+xYIBaSIJi9XwiONizLimsDIbd/SWx5lKZiZVFnpv8+1yYPpTeA6hOpLC+5tNxgb+YjTa
tXkeTws50hypV75IYzarKS+VrjFnfyC5ZB9vmAWRCaByyGGnHbWwCB4uUy1FFgvYmo7o/u1zTZyF
EEXgXiClDIEk+yHS+msq6WyJteKCO1xhAwih6xAwPQuSeabupejxHLF7uLkulJjhdH2UHTW+I2uq
EC2n8ziqLwHme3ZPCfvWhkN5sqgXx18NeJ2TNMw6el6K+HA1OpExGa0zNZCzrppFleVE5uKuTh8d
ecJHcgW60azX4LHw3YvNbF0rPvW7kVLo6FRlcgEkB4ag1zkMyVikL5lvvIaWZ60LI58/s1CGVmEo
Xao7ntYBIdBITRRjIzIMTf5GANpxSdEjj30PRnTsd4O4mqu0LhxKSw98AyeI3QcOwNchKviHtTFv
M9mezrRmHzCBXEce3BRtosh3DWFz2MdyQwG8MPF8C/klnIIhz+oAhRNR4RJIzyQf6P2aryCl5mAE
sizPQA0PD0lXfwYO5iNIDfo6KdVJdwn89ZlHwBM7rukn0KAS4Qfycr2ROW/w7U1Cg//xnIOH6NfU
twbxOgrFuINXX+Cy0XCxS9XhPTH1iIInORof9SxdwF7+aaMJ8+oKCAhaU24EhlkcGkfMaY0PrYey
dIflm8U27pSxBC9X9JRXMuExPSavA+deYlZNi0rSfjVHARMPZ28HFQQi3s6UNcd0gEjpPsO5f6xC
Vx63eS8m4ZYgekscNuk8O04kPELfF6ywyNzIERh9E3YJ66ZG92pLHbB0FzbrFYfIkC0o7grnySwj
Fk8nqaYvLpwrQBsl7JUqCZkXS2j21EzCi/zLvFYv9yXdQ6RAZ25mQOfA02XJBd3k+WNA8PjVbvAd
r1R7Z+u9/f4KsQQ1rMPzroKzwhVIWBSuKZp3RoSdvibahSPJPBqKVMM8HIlTOCEeLQVJkTnXKChv
CyOZqtG+kmC1Gev6TC1kShv+qdCZIIocv/702l2ZSvXRtUrZtNT6hYsFU9o4g+kv+WF6mxeZNL4r
gjuC2LYcRlajaIyIhgrXoLoO/5SoVfuOLcQnpNYvmMNPZGVg6jPCDwpf1DHm6wjpJG8GaeonRNmv
aKYHtxzMJHGfsB5TxIBTgs+sJVWq026Y5jVzrW0HRDO3CNW5JmW5QInCjiRh4J9D082BKi0ZBzpo
zBQzOKr3w4ISYPCLozNV0WchGixBNLizOyOUAQ8NuBTjCLuc06mNAnDm+zTQxFA3FzYFgWvu72wn
LZGqY/oCaskATIBoSmqsDVYYtHf5MXnPWGXntmn7sB+5ww/F/fa8RlEwoeNxzZGjXqM7iw3rzGhQ
ZPPPxRhQvJqP0vBNn261rdCQYWIEGpOP8GfIRgbcDvvrNOMUapxxcfsiWFxP6F8zSXLV9tTrAcfZ
6bH/vCRpSW0ZQVWfj5JRDT+0UTMm6M1K6MmBMgIH7o3+0CTxZtClhKbrpiHMlydbnnQtZ/NyFQEG
MEuCf8q95GomFPPG64ocozPnuUh9hd6NDBN6sPth4tTCC3LTVGFAzacw+ksaskxIYycHSzUJGmNc
BI8UyS+S8JUSxCUPgBqboL/WmsXMbs0xXUw5II6sAEck3owNvd/xV4do/eicMT/lRwFWRIEELZUI
xmxsPNBUsyLh8cHphLpBSDj8auWcpoT9R+XpE76KBjNlTGgQXvqUHRA5Jsa6LixSSTeif2E2+hko
JD/BJJvDlKoZvJ/1tKMNxuVhHGfdcNx4vrtYhG4UYIYJw7GkI/C+Sa2thRCeG1rWh3luWlS73y7Q
QE065DcY1pWS6tph9JURZzw2yIefdmD6bENRpbekTne2Nbkjj58HTwvpYzAOfmR1MfCI+/Z7f4dW
6q0B/lBvPx4OBHTixrioTni1WgjCimCQgNcWzCKojGTMBIGcpfCUZfU4Stl0ohqglxtT6emHmcPp
rnY1cEiJhX43OseCvfhJYntaW2n5V/hvJc0R9QRLaJakI9oYXuxRDVUepBkGtBtQvX7fO+pZvQl1
WQDmfZlZ8GdvQJjo7azO6HyZNgs0LHXHVNDfekXxYKWlYnqb8DQ5uiOTHM9p+AcRkAzvaYE+ehqe
WrK8qprl6A6rWxbRkAO3wzuaTCEcCCI6tQ+CQ3soWqBTBLJ9UoxvrshZxtk0X3yzllTp0gUmBjGd
dWb5elVghcOG8z4sl60AEew8GtK6/8HHwRBMeT4+Me8V8q7uiVm/14Rt32OddtjKcH5NciIZb4jY
RDhBTeJKaLwqikovPmrq6/nAPesdPibbeBBxGgyKnl5a5TvhwTh68k5rM4IYz0bF+7y5akeTSDsu
RJfu2qNkf4hVaSKbQRMIrfNEzkg9CVIc8Nrmrn6TFen61rxyyNZ3nCxHnfyeEm/rxHIr7ZMG770v
w7zY1gGSW8LZ+itgn9+DbmMG4xVDA2X1/ggk+lP9o7sHgQd+hWAh/scqmAx3xU6R5yO1CbxBhQPC
HOty2IZIvZrT/eUaxBdbzgecLVZDpBv8JcFEPjVwu2CcIudFBh0w6/jiGen1U+2rgXVxug3B4jSv
kOnkCGLgKKe0aFchFO1i7hSa+14+ZTwKxMyibLVaGNtp3FAD3Iy6yqLQqspa+L+vRsYtehqgwOay
ppDubc+42y5YS1FIXmiA3OTz1qGfKscVNYXqrChR30FrbJBONYtg4jp60blO3IEltJFY+QS0rHHS
VovVF80ay19UqUr0eyACFfGivmzsy7Utrs4/0zyIL3Bdp9iZXnqHLM7hFgrTvPAYnVuX7mV+5RRO
9c3euuzt0SWn5gPQviUMdK30LnA9R32ALYcSjuRUG8VhQxk65Uf/rmdKV1t686zOfzS1ybdi04Zi
0EBj6PKKP3Zu1TO7GHcmL9ml3rzmgoEyodpXsCkPp3R8UXPXcsYY/yNqH0dawl+c1hR/UGP3YH/e
7259/Anx3z92uJf8m0hu+clqve+OvXORWEZUz34kYpKTKXhuuiL0hNGhO0L+PIlwmyekQqdhH3V8
ibqAhgN12FfsbC1EDPwGsy6amt5zpFALZyQva3e8QpvT3m1ysh5NE3w0W1FBILuz7Vi4AizL4fdS
r3KtuJ+EIqU0KylbB0LYikI6c6uDImmIaX9RJaXZ9W2dgyoliXpaZdB0puf1T/QTTcStL+d9mtwM
pzwIo5IG+BJQpjB/23BclJbJYe8O0HMkakLagB69DghX+pyJBaIxVykOu8/pTlJjmQCvU9t7vQ2N
rHXvKPAULTd8VmdLCMoAlhFLLGrz5qSH5AQCtt0kECr5cRzj+7EwkZJyLWQixkK/qfwRo25R/pk5
I6HxqwbvNaNx316X3ETvo2pk2zk0tL+r9X62FdG2t3jsHQA1A0FWM4VDRX0o2Ie6hxXaCuTgHa1/
ooyugAuSqzkwTF/1wiprwYFs1QcA5WM8s0eH+4yV/wYjUDKDOsXnw3VZpSJVEflqYXscCanNpB7G
ESvnKFO5Kg80fCagq2krJQaqkZt3AkhX+9EMSb++JvG9ExC70Xjk7lDPeQdRkpb9gTkdp5YAvNmg
nr98BucIUHZ9h/rxOPr/xE70QagP8ekzGSZsaKGUC5QYdhVKG1ySfNKjEI0dBSnkI3PYTNKh6ABN
sgADdUj8GjYGT5pVMPB0F3IZr2cHn57KgdH0O3d7FYiq2MVFueJK8LQWFUUhbEtPSxA3waP4I0N1
wZJk9+03dhY1Mea1S6G9N7G/DjYr9wiXn3uKQ7dlhrp/CU60GBohJuNbZxIpqO50++Z3XiIUSxzw
0IYekm792cJG4jKxO8kWO3+2VpKXm+lSJegpIKHaloyngrkeT8opL6u6rMOifCKoq/H4o9X1Sze/
UgqN2t4OXe/zINC1wFknSExrXuQsnok7xvHQeyw2KSZnMKAIm08rs0FkLqV3rGdLEHyjvSfxPw5O
42PNs/NI/lIgSwSXnj8sXXqOtfeMS2u+0GLTVLBLSFaYfPQaHYAw9IDuBorfzjDEynmeqZUQFum8
MiK/jcnIDLgPcA6GCNm6flNHsA6OohfIjB1dtR2AvzxweBWnKc6eIccsCNCC8mqwSUXM/2E64tEB
QV3ZnJx/efnh7SsvYAx0y6WXJSYElB1VGKO8CCtV6lGKJ4KN3ExkMNcfh/JSbn/4e4//JCTV8zka
QYffIDyyPEfvq1xUy+CdLen/MVJRuszqs4plD5FykvgOb/cVK+tINKFtq9uwXDrOdz6UBhTyan5L
Ud5rKPUasULIFu77FHJcRxb1kKhxGqjPlabWyoBkaabSB1vyARZUHcjzfRUGUAWXf6DiVN8maARs
oV2xa/qNwMmov4W7eavUpESP/Srq6paBUPiWsDW6/OdjqN9Y5MYwv/Gu9sQu5PwQ3eLQ2MqkHDZn
L6UDDfvrGuGuZ11ZyqyQDgZoaJt6MxpTx18lKN0n2W9F3szYYskaU2fIPgnXprfMK/RXMY5sddhK
96jzOdE340lnKKtGvqlwPjk/Bqitrc+zzMjyHXZKz2P/T+Df4OCu2CtScgvamIJvLoLtXhuibgBi
iCkS7fcgCg5RF8M1k1VOqVpHaF7Wtz04XbkkNbJzXD26MxfYaq3HmIRADgs9jDL6HD8IFkXDgxm5
N3tM3Q/NyR8D8c27vinBsR1/e+Mz8gq4i395n7EjoJ7+/bqnAWALFBP7bX/HL2aP/RSz9zdsT0Ex
tD2WaZZm0XYbNtkg9mKBf5z4vTzgm4VKLs9VbTSYnUQzcZKcu2jz/Ng54k2uglKek1vcXTJtKz7q
8SK4z1YtEiiToC8JZITdVIwQKtNYx7+ZeD3SUVxucIb2yc/pCJ4eqGr+7et+3TrbL6X7+aPg6eXj
hDguvHexZEi4mINkkXtCOjIM6xLY9TI5ezIBvvp1I8Xz39WEbVc4dqopSOxm1lKIDAjPpRPKeg6e
CaTXoR3nloh6CXTGvhIDmUtFb981+ALmul9IyrqM8B3UoGQbp2rQTZAUfSaNdl9QRiPz05Ku7Twa
784rzCckIX3BivzkzxiCam04c3DfcnBrE4rTvpvcoKxHQlwUjfruOqTgLy63YTajaPw54CdgHrb5
LV3g8r4wOHfAriMKvIOJTB9nLm/FtvnLUSOjY7wHY4cTuNYYStL2w/HXRoKu5wdlbPPI0biQmJDS
K/2Rftd7BBlITyHYQliENRpHvUzLSyazG/UtHy61sSMXMr400ob/gXGXc7d9P2Xd+9bYv1gM4vAi
rVS7WsfMqrunrbSQJs8Tg9fMErOUggqeizGocpJB1BXOT+Ecn1FW8pucX8rR3WH2ZuAz1gykD+hS
tvPhGP9VuzweqaXt1ifqtOiX+szSw7kJ3/D/pmm3FDxKNGxmHKRrxn9UyfC5ud3rtIBiabCa4kWg
BS3MwKH/TkFpZekP0tHV3a/TljaL6eyoFKe7tYDvB09tAGZ6ZGN3vzsFUO/tO76uUk/vtacbHqXY
GUFgF377riF2ts8rbYtQFhkOXJaVM043rmMhd8GtsF99nkSrVsnMWmV3n7ngm3JCzwNHgjQ6cq2+
jRUSsRjKwFJrmUHVeCWKg5+OcSMaN1BwRz7Hwq4CnN/3myhM04fCeTAjDBJuE9HrA5KkwZ+nzMnW
yuCWmyLdvlQEbxyLo8rlOEUqRzVTURAQGkgm3N+bIjXqV5H4FNKmmcVrylELmqNcN18lCKvYIX2d
Jfsmngj2ouydlEcMmTIUMkJskWb8ZO/YPXGB5wyOv2+lkV3hZtxqe+gtZHE+UCJb+2ojLzJK4hyz
NA7A1Yp8GUPwaDs0USDOXkdM73nwdJ7mrsEau7vq07oKH5taribRGXFU9qLcROsB+dIyvnZbMvTl
Arfv69ZXNq3Hf0jGF0kEP9BNQMa4A6dANskq2aVdcnJrImMOWRR4KBEfzJkmjTwgzZshADZg2pAA
go8l8dIOIIhqD3k3Mr3IyainiUBkjDnlsVkNH0sFRy5eVJIYNFKhcobmpK0LVg6+EBZSPytzaanT
lpb7c8B07BRQWTraacuKH37tcysUfWkU16aq1juBpRYKvzE4K5CRVUvDMLp1H6uTQSz+VXwzuAvD
eFfKEKKgJnAB1JhpMlsgtiso9Xjem4EHVLEAoh79bDU77yErX+WFDgGM9C9jugB55DO7n7qdDEro
tKBtUs9m/CxYfmMUc1acgLdjWhy+1QIcEpOf3JTRWOvolw+reia2IP+adFYfFB76AeUMNprqwyAf
vryZRANDKP5Q8O7rqWEdVq1G6DqzzGRr6okPldCZSDT5v2P49dwl+A35I/nhvQMUlVezwOt6XAf1
v0MCJCQGvZP2b8D9LBra7XQ4igl2fs0cghCljjKgYHcy3sIH+yxoQgqulhcY5BE7P14aGZNyMjJV
X9B3tdLF2RNI0GWGFUZnw6UCDG5m80J6eNVLJAexUpnztWIllw/r+JPDEjkF8PUtRR3ld9nO8jj5
tUicPavDTPXAoQhC9/ayzupQwFK11nHSDdURO7O3c1o9XssmGQWTCgI5pPjciFEm2aMvsnB/+xrK
9Ln7BpxBfvqXaQu8qezD/b/fnyFGxt/ynsiyuOiz1KBfNA3zLD5NlBsZl8KDNylStE7WomsH3KIx
0EdiRqvm1sy0WQK/qyeXVUtGgXZV40piDYJA3QSifRADMZbyUPmUZ+xt+9L2Af8y4Meqt+XpBTOw
yBElqj8ZPsv+d0dDzqbiGEbl17+5/Jz21Xu+IL5Jnvs5rz3v96meIRzRIzZRTJXDXPlnnkMLd8hW
3vt+lY9SPpilPAOqbk5hfXC5kpAd8qhXBCvD8x/WOoxdUv+fQR3x3WUzED8qFMh2DKd3vMLy5s7Y
JzVRyY/78prVRCCybhjQwXEIraMJEsstmYLk/8iYgaNOtfvxlw+p8bUUmccbzyEMWKPzHYxgfUTK
M6DHvN1IriMVb1sRPORLg2a3QGBxAo8tZuoq3/JV5RRnufzXw6kz85E7WVL+VYq2FjtMixUZ9Eut
SYgD1tANfDzbpuoGjdHiIho7XBd0ffN7OlkDnj6v55scC7tMvim/S/jufvFlx3bg54N/F+bVKish
osQJW/IEuV8gpsOa2LhwewADnkg6Hd4eLzwWFgMAOXV7rcJULjZS2CY6EPGkGpurz+mvT9JhvbFE
DzIn7K0i+nlqQjMZF0OWqyCtBVpl5GgO6vql1qQe7rHEERpJv3drkZRlXM5expAkwMKzzv6IcNk+
/ypkHGL35sPEXQtwBgfnCAyX2nHR6o+8XANr+mjMozQ/WtsWkptkTgUXz4h76ENKBasJQo+9GoyM
x0UocMP7lIv8wMLBV+FGGMb16U1AF8toWWqiAYCr1e4S4rArRsus3r/2dEWnqk9m/HvNcbhP3tI2
GyIhGxQVkoWRg+5nOd7BLTxPSuJJeWqPLBUnvLpkh0Hc83tWnzVebiRI66Algb2DQ8ThBh0YWudM
aXzJCS6b+bb/KeFqMwYFMh/4QWrUkDOFF+rjDvyu8H6nBtyWqjXmh4jpknizG5ZN3eKsP0Zx8MW5
+WH5sJYPXbvVDU+Cw5DsKiKgDPz87LIj+qm2sOTwaDf6zl83LX0AVYrOC+f5/yLnSKqV7O9VrLV9
PA/pN1SWQaQAXRkXkfBV3AL2LAPgOBLg/NeIJDW/uOT/4SAlNjceRmRlqdmz5LbD15aceS/7vGCK
feSfsjxZFPz0iKuc+qzYVv+3r6A+nDM736sVfLWsPahdUVvnZYCafm2LfuiSqPyVx0Uzu18M+HNz
I4Jpck9SHYLemffdIhf/ejK4DXcOI4RqO2RKhxlI7VsbqgY75gVI+7j5A+EXlvaQ4siFKN4pWwck
hM5SnH93iEyQgXRlq0waKotLhDVjRfBFxhfLts4yM5VklydK3BMNzwuk4IjALmpvihJU+HRZbFZX
xkR5C58PMJBgKimz/Pwk/VVfLcwUCQ8N+AFixoRQm9osZnScpVGfV9Du76/DG1Md4U+mcQ8c5cbX
qFxz1R9ol5JqS/I+1jEEPvlV8jZQgz6NdwKnHURPCv8Q+2PjewpAhax6KwHUGVbwnjE79y1ZxHaX
Zj8bO7XWu8Y9+Uks2XH2IlLEcYYEhzSUlAj/2vac7GROcvlpLWdw8h4FjiJXx9AIhWdDeiX+dK/a
DnBpPwhXqciAxlAYc38dWNtIakTUL9xgYxrAWZ4vqnikCT2fSBUPgQmBKxn6uv0ofNfR7ui+rrAk
c4zig8lDdh/fLYUB/dvaLPKopj9mCr4T4ijCQarsPbw/Nf/Jb1yn2HMliTJJ/FSxGv5lYdROqcuj
e7qqsr9/H/8bHrzlx4sYWzJRHYuD8ZKTbcNZ8oTzQhImOGXMfi/p54p8qSBDmWxh8sz1ruXHgSYh
JlL5ENSpuJ80jvwJqY/aNT4kIPTHRCNk6fbSwX4BqEFxANnKErMCbMlEpuJtW6V9OXK81NyH6pCj
AIKyjXtrhc7OSYN+mIastqeBd5VVQFO0GAtc7UBLLLLsaNdBS+DbCKdc+g1kL9s5KGxXcXdDv6YB
sNGSWI4pShT5wX17y3ltE/K0vrg4750NHoenuOc/S55kIZFjw39tZgUt62+LdwVSFGdfwhJATBcf
Zt/8Rj32VQJXVzOmcupzfGOmenyL4E1jWLoGRr5c7bSpipN9HZNCpO6bTjmKpN6AJSy8d64BrmLY
7cF/s/GVZ1AG548yjXJnrIc39S+tBOmcsZI17Xn+iWe05K1iLsq+jgH/3QUV6PuN69Uw8KtqqexZ
tLY9FKLB2FbHRJx2phbT+ubLu2ZMm+Tw7Q3Xb/V0W7wor9gd212NIbtj4cCaKckw1obcGDk/K1YY
CKKMBWKWQU1WoGFwWgypx4zoey14T8GcmvJCkinh+go2iDuvtOWuNfP8Bukh8R/aztFx14uXy/uz
JRneusx04OVIfby8BTJnwRup9w2ocmMzRFaPIar/yAk/NGjQQcMR/Fu6onEUQtqlnP92rW7W9AGZ
hENdYrgOyWCSymUnrf0Y9NENC6yW0VWcG6wxFM2MKzJ5cGJgMukX+VePtspHu/0qBTGtBhWWGTN5
wwQBZPUmtWUteWwLZttPb4uVQlh7WfWUdWj5gDacAU2lQxxVzBozsgzsy7FvARTKtsD3crGq+tbH
kZ2cZzO5EIOWP8M9zQatzLfkDYijul9AY4rAmmz0fL1H8A07oI/lXgAvpy4GoS8ZjbEa5EZbi//3
5lxIvHD8MinsYszqVUww0gB57RC0zbA3ClspW8SIUon7mFriVMy1bUFwc9vgg6v+IX1Ph4XMwJ6+
RpvumPzg7nvjCYozqAlWRVsyotojrwnLkRBTE3RZjZOxl/qk8AfQdS+hbp0v7VQxkz9tmsP9r4Ov
qmCXKcOD6vCTD9SY73iZomuCTye+hDvJM1LZrY2JzwYkoyqLjkO1ldtaifQZBOxtJ/FNw1XzdhLM
dwHRO4U+TBD07Usiku+F8zTQLJvGJbPZZg+T3PEoI4fgQG2Vordj83KGwOcq+3GqUOHBYa75s8Wq
aSk4PyZ/0R9Nb8MBLIWeOBFhc+ipK0TxecH16s+tYDmqh95WqFpSTtxpQou2jKe8ECkVUVZqwGRw
UR7HJ0rmyW3Rr89tVzRPVsk7vtqi61xF3KtnvFssC1//UsFCtLANydxI8AaPgHnWmznLlUC+fUhC
gTyt1zIXrxu5Ez9/3wda8AlHZWS0vRJKMigyCfXcB2EzPO7U2oWHA3L3GBE8kLlYOTA7i2pWNSfw
joUQ5oz+xYdXfLhMCiSmhFlGqHAF7zX8q3+QBYmnniVjIi3CGIt9A7Qu2xlBoK0aDplRPlCe4i76
a7TJxoNIsjhTxhR8/PXq71AOYzjncfh+XKwKSJMXsKbmmwvmnIjHN7bCAu9gqhB3ILvsRvrj2SM6
TKAZe0JtJb8uONFeyNQbkf+5ExE4Gz0DLMQaoDAI4snaDS2UnxdFpK+Y1tNJyk0ORxtNDWeTQO3A
8Dp91vmB+mCNLJtjHbnrd2IZlA+o6BYlDOZnxU9T1cqRcI9GPnGWrCphZD6gAKxSOHQdBw3Z9hOy
r09vMxgt6Di7rImx1iZgOcypRMHrsPpbH/eckXSOmSZxopAbkd0rJE2A3okPND6tykDTWin8UQ4P
vgya0ChUgvob9leRxX4+zEKEVt/DqTcW+VlQwJzZN2gmUWEm+UnDUearPH+OvA9ZVJB7KnE1Bomx
g4ZhyqZ667Bi9MqVaZSHXqaN35wnbDji2X3V0E6DLoXH+IFHZU3ZbxkCjVSN6rhRfi9Xn4RhBMih
tCl0ftLNHXng99YP5Ut6MXSHBeADNRpNcU/FCsiMc2AfpdNRqaoY7TS5L7pj9jGRpDr9vbFwx1Eq
u8W/Yp8isrUK8NrYeF4NJLDv/vacQSEUQ+6GgSa8HKQOy6n5os/MHs1QCzVRtsqQ984paGdnLr8Q
wMkDLVHRoSJhRvgUhxfgywjxdjNingNng3DFkbVq014RASmZBHwdOeWnZ8jZ2/0m0jkqn67Q8jPZ
RetSJpXocy59t9OOswebIN8unNt76mhM0n4NYUW5XdT5YhYmPJRgP6XDGnXyDT2ssTH8uI79gQcl
4IdvFChkt/sTLe+2a2wXEcPx5J5aXS/ihndyUtA7ZXuNpDJiTJIsOBn1ae0T40TbtO+VimvnNBUC
qVRyD30jqVTjDMRidaYUHqzNJrqqIxymslgrMh1z5okSGWPh5sdrs7DGBTh5zEpixbCanSbEW6Yf
VHPOX5/PxqNEhm54+fMrxuww04PhquYIq3n4wAVzbhBdmyZM8nw6rciylzilHkOlSkFzHzR/6KRX
Y65qS2l73IYk5hijL5CeeDsTYSQJBdUk1jJv5JhkUDgOkg24jFqZmSdms5pqZwITeE5PYjqaHJrA
VOeRjr+1lX22kmiOL2dAJWFAvs9reFKG0gttYaAQ541BaTVqWS8OUTUHaE4EZxFEEzP/pWwTMyQf
fErUCH2WUS2++4ER0mYO5cGLaQPVzKRv/EpnMa6SQ2J+N7fZtpEzHlg8Z82SSNp0rSC7AMO+Vc7A
f0l4InPyCP+0Jc0t/1kQlyjl+QpHIwtp1GTXgWNZKX/l6Xeb1cfpwnB5ZXlg5S0zAZKGszwYSLSk
vJUs3KOb6IxcNuBjpNIyIuITun78983goZ3Ub0odMKVqwQh6h9ZO4A5xt1P6GZhqPgJLyPTkB9K2
1U8E3XJAy9z/PgLpNuUxSVownCR4x+qJlfFuKVSJtechIjsQ9RzhqoN/7dai1sRNDBKmJW1nzvOu
dAT18/L7s2zVzKRNSDOLECsVh4FYQnkDTTYgPKMg1CLjlZeVEvQK4IOzqM2VoKmpfX5fqKd6qy4x
JxspHnHfyfB67Z8mby07l7CelCfHpMhjFeuVphxEsg8yNd/IzAIA0H3YEUaI75HClii9zPL9Eh+/
jHQJhAgfW9+rItVnPA+efccusgI1kMCONaU85eie5CG3PjmRymfFvQ8ha8k8HMg4Y0liRIvopz5h
SxKj1g3+arbKI3rHiREjxt1PmNG9mQZuGNSeHrX9vm1WbtoT6I0PMqxf5nrr1S2oo6rrjK4LIO4g
eQU6W5NLNO4XDmGwMhN/fX2/u0RTJ22qwolF4vPNFg9bCwky6mc9g7c+Qcn32qRMN4nUjHLtrpuR
Qlb8sKUqlwP/CUKgOPqqL44u2lAFUnDzgZIKzv5wuXbAOlB4ktCQmK8Vmp3VKPdS5iQtaPhUmc/s
vTkBje/VgMxmIqICZikmFrmRlruJkU3hLvdeBKiLrHtQRw9GDHDs2jAflGu1YbA5qMEzphSBMzgR
7K858BQp59f48vNtuNJtt9cCMhShmyqJ8R00rZYdqD31iTuKfIZh//pLoi4RZVwJsNyM+yY9lspp
SS2UK3DnuD1K2Gwckoj3Q9xhF6MFUMLwv2cQ6XY646dWwtgBKS/c/0t02hihVdOIodw7HzTcxJgC
uZ0uIC6VRJ0r7b8naKo0jQBvsrGiLDObjkTbrSdDqNdjrISqc2JnzFKFayAnpiKx7t+OxhfTOdy4
QkbZp7WgG6cl7kZp+sbgsjj+At7r/9y4UW2pc1JEJZT7hK2oPwxZZApmuinprMuVq4knss0klHFT
0kVeyCnm8LC2Ju7aBR0eCqXum9vTWB+Ty8xfEsw9mjYKNsCO/A1TYRktq+uRLJgVPyv5wFrtYjdn
idxqBPH9nq7zt0X9ewK4OOlfYThlqPFst9qQmbaX/XWxJkxPp1Lk4c5a7hTagqDJw2ha4syjaarl
SpQlVvBQ5YzZHLdbndFhAu3Xt6960Ku9qmCFNuh9IchnPG9/9WoVUcrx00GXtajQP1l0DaBRCIOp
lUFZxcEByxs+UM76KfbVZM2d8VzN0Ttzb6uFU/ZiCw1BUErZQr2euG7nSwrfiaIGwjr2qOS2m55S
Kjulv7AsecBOJYzW+//ruih7U9dU/9s2T5r/gTrPWh2LJKrTV1k+xOmA3o2oQEhpO9rePZcCz1VM
oLdsFvlQDx+PqxQHDsQRJVy+AYENryHCmsKaN5XHYYVnOKkBBgXGptOJHTeLAIp9QOh84FK0+hDp
7TnaeJH+nVOBnH3PZV4/YBDP8RtyBazDmTXtbkRyIgAXVEzRp8vifaQBdVx/qwBpNRrMqKnLvUf3
j1T3FPZHjFYAF7w3/Odcjuvi0T3KIZ4QBnNBj8k1ipeRS5OgtTFPWXJDYAeWqS5P9pbjL/lGZEmg
u7Haj5/E0xEbuqJ/4GZrb3qHz93FuVEv8cOjiTxl9f9BFSGXy07CiNuOEqjGLANL/Wjasn94TrgJ
MwW8xLOV9M4djYz+cBOd5coQoxExyFV2MOVloCSG0RBpkY6w7HNg3TVgiH3gn/a9tT7xsQqW6fhU
d3KAtEd5vzvGRkRwzKhGBQQmIhcmgsW+u0Adws/cwxMrSnL3i/8mXPLWvlAEzsjJHBwa3vuw8jGZ
tGlWGM5PRtxWcNPJjjE7TCmqUaSwBdz6rY+b++HY07xUWuoUfVizkiJcFF0cceAuoP3Z0fNjELQ3
n/XzKzPW4jKCQELhEau3SYeKbHN/s2PwoorgTuvhEau8EDE7Qe682gDMCPxCUCvBzfEPIijD8mVf
u5Cp7P+CzJyKKB5QwvnmY0/ZyFV6SpG7XDLKMAFo3N4P3WcjfCs4pnrrcr/8zTmthaLFldPBw7Xb
WXqjiFfaFIHcZapWf+3WXM9WiH4ZLnFM715OGwnx4jrL6y/Nh0WMMlxc0htBt6MOxiBU3vBp0b2Z
B+SKnsmNMBf92GnpOSJLnflyBz+1UN0wji7LcwnrYfBRyrNvby4BRNVLfMamZg6sDIhNd/I5jg0k
UkvyUjoKLNwy7JfewBUr3Lya4qqI3SDlnPkzVI2rLkiSFvAWjmttpn7t396Al7uesB//P7ccMPhB
fFvD7BO2Be1/+BC3+HmtclWVVWHPWJXBNN8IVfsqzlXHKqXZN8eTbaY+dG/gCEf6J5Q+/yjx+Vbh
faxm9iUCqMiF7vEfTsApsmPjTfyDDRXAhO7fnKpMvqI50/xmVLdXTF5IQ0r+J0HEZ59ZjWJxrNyP
VjXgzTfv+04x9YH0x3g+YZjoWXoIEOHNLezroFoFESixrPWcZAudMtR6HfQt1K9i5j9n2bqlvieV
EKU3g6IU02N9x4aFkC7agbeL8+7jz42n1sooBaV+kOJHlZEMeIswk5ZN0PoHTfKqon/Nmc6jvGom
Yt48thncZuzN96Rzfp+W8JPtcYjyTVvModk+KqdI0oBVRv+DCLBLDIi2NDnrDyVIIqhMS2x8H1zt
Ena1BtP6Gg/T9SbWRl86X21SU029c5DHoNVSt31cYECcecdTjvIisinkMfN7Jdm/W0zArckzua5H
aqGQFsK7kdq/2PQXCZ3ejMivvD0HIDIFSZU7HQW3WqdCEnpUNHP+bclXgg05yIEC0EQyr+xTimnk
ZQItOzRGYdDWmxF+oG0egrqU671OOe3/zfENZUwupCxbG68Gylw4puzRpQW80BYQbR4dd+qaxTrs
aSKnl58NaGP1PNsevt76NQXvG0tYjBuFl5vSrMiFuHTbNv0wQgT4XxzfB9KHcae0xiPGyf/0IILH
jezO6RcJEfuOPE/sBmWUJCkWJsoCXRYu6jUQM5+YmmylcHRtEecB2u+9wCwK8S10nu7TL0Hv8dlL
ykMdZyVlVnC5ifeh+WSurYJ7UEGkkwQsv9mfsmvK7MTP7H2SBPTU2Z49/bTYK7fR2boY5v/Bdw60
i6UUpfor1n4xgjogWNmTowT6W9LsR6q+rqPn4GiwlbhKXHBMZVVWDjkTxvzGO8CSO2tIwoESRIfB
eri+MRqIHb8x5sqXRa3KjjaLO3YD2xQDjtsvn/RuURI7KQMGfoNFLjvOmXBM6xhPEFmrtsTqJmY8
EqNuEajx5Eq713fNMVoGk53KBKaBpiKi8p3+9AuYxI4qF4QPKTzcUpbHqEoNsUJx4A7522yzrstG
8LbW6iKx/ym+WnpPpMdRlpGKYsRovbfzOu6oZZhJbpbf/oQrBPrsH/0AU5TJR+dgLIiPrjKVxYxe
8BbvBmQ1atOulcNr5sk11xOaLhMeN5sRm8VsnbmHbppWFZoIA9du3jejmnwZORIEp/xIBIk0eeA3
d+iMMsChvXjxJjRQUGFCRFhB8psnNxuVBcMJ5L+yGSt7lfmgo1YtVeQ9BmiSpT06P+nKG6xgU8+b
1DXLaFdcomOuY7wArskv24Mw92r9SXRQ6YcfTSBKOTefkMTspG+wI6Ec9kG1BL5T8qoGahDJIegN
Dwudamk1YJIWISN5g46ITz8/tsqq/+1c6eWOyT4PMhuY2cwJd3pIzkl0jntoosFKMvNIqqsQQA3E
Kfj5E2WN2OZHH4JwhzODDqmG34ASf5n+Kz3/f9dwSNEWcohU+OVrH00ghX5+YmP8VbbJDnObkIMp
Pb7k87PXcjCS06hDwZjQthakXQ/YHiKqSdSAxLzZW9gumElTIEPTKU1QaBMhJ9ujSi+vl7WDGp5A
+SiBQ/QZnst0gASeak+kZa5V4OVnJd6Tv7BC7kXhLm2nE6SFHjSO8zvoiVchQnV7R/KZXEzlniBV
lVxNrtXEO0OXCVwX1Xi+cw57a6auO0OSlJc9L33IW9kTUI8NLGuXrSSDTEmasBP1yXZaeLBlbBzi
OUQPTyEWfKfcXQJgFjw/jZhHLZwLoXsTpV0j6lt7D0WAtwxifaZsQK2RDg59zxx+K4Ep5AGeT2fz
qLv4UWXg2kOWhlVaRgvjRiqXev0vJZG26sZwVS1pK6GCrULVcPiHHNUA2PtfUWx51v0OGT2sR8HF
5BGAYEaTep/+9T3sCXrotg+O0UmXXY4HDC/m/TAZtxzAo1lMz98BuVDoQqGpaP2L7UezGTFoG/rQ
j0zicP8wnTj01fG4gPMNjwy7ITDRheUWfmwry0WdaqRFRKOVntnBwEkxwRSvqwXYK+yjhG6LknWo
792q6UTCiNjlk9PTzAbcCH/3HKJn4eP1Ctq9kEIlM4iQ0vcUml2IE7RdLQ3pitW9WbxSZAtHoTFL
X4hF2omjSOTKgg+xbtRF/g43PeEbgLqO2rXxLQbVd0boG7ip4W3Py6eEoe1T5fSqrfAtItwjaZoJ
Qi4DACBoHcFEzjfaHmSZA6Olqi1JWV3A8umSbovb6gBbnSRgxSQFvx3gR++5rr3d/PPUAgNJD1D4
ACa9vpdVK0dMYXDH3e0Bzf5ZGFq7kjBlMO7w5f+zELBnxPNdztu8mCq1qd6Ik/W3f1PZ+IX6pgtY
NLnh8ACmzcKPJmokOnhWcX0e++fGbWV491ErFocMGzKdZo/XRwYLcKhWsYgzfgP8Jtz476sTcRIm
pbKG18zHjKFWBlIRPac5xL5iTZn3eoxzuKOsCANy9gM2pecQcmno4Z0s4dLWVjGE7yRoV4JmFRvl
zgSRg4CcWq1RpESJd73n+5zpl8F4oizEgZ7Pb1FwaX/zGvASrXExyyR9q5w8Y/VAbH3MQ0UsHqut
Tb4fxRsuFISsV0uURn2B/4WVMrGS+48B/N5Xt2P5GHOsh/ILkQmWQ0JFj3x9+UjcmmyVCWSFa47i
digEUyeAQkS5F6yeR34PcctLSWh4j6WRjAQz/ea86ODDi9jO0/95tB/niG3FRRdYmtYXcZ8tEtul
LrxhjAgV2kfENjqaNWdFyuR51raC9hr+NqGQvMwtvLzfLqEtepimqHK/zyCm85bB7hNrhqwmbvdz
DYCWy2Grn0qlnlM+nIwXsEjdjYHpQ2YuXiKMdbTjUfAggyRR+c5JR2BRn/etPl16OyQr2rejy7Ut
R/BOZ8+SDhlklBJrKIGMkuVGRNPleAUZC+bNQLVOblL+9KI1VAFEMAfkUdBZ/ohNjV0htueuUtWI
BYje8wpS8rFrTWcO7oOawIh18X9w+NYTHZGBfLdeCVt2oDlzKbUbP6lp1V87bTyktCQQem7j6mUK
jYJLWrjmcQaImhC/kIUE+UcAXgoCFuxkM9AGPiBQSLxjmXdIwN/TJg/KYwqiA6hBM2uHOz5Sj95a
46cn5S0fzNLkTmXf5WQCkVwIFmLOtXbF9DGIrYGky0VPqfZMUjpBMOkxzpyWgDDddEnjqPqzEQrr
WyiDbAc4f+/jk+oV72W7AgzSRQ/+ITFVIwISkDd3NKQXQE1ko/uxt6lbqLAgkOlUsJXayn8FipLv
e032D7Rn5dv9m4ojl4lwXNJhs3tI/sPIbdfV1WE1jDFYh17vuZtJi+sSlJiFU4U6bycmmQ+gyYI1
ZpDX1MoYg77RNyI2UWfJmZzWIoL34i/urlWhEoyPqH1w/8rY8DQQ0ud73Af+Z6wZvlm7yizdICKd
2kN2vUM+QJZztn4L5s/0Uy+ViKRVxDewS8cuHqFU2Ol6Z2AGJy0mabcwxevyxAOpBBna5D/TDNIp
7fUogW89EI173eD8UHaOnRI7RlN6JKpWnz17eAMIIS6uepfnSPceVRDIwBddw2LSQNPoz4N0pDqa
1AcRr6rjvVtP3D7Kz3gpERVXqW6j+Tc2CryMigbP2I2ZI9SjtDWEfeTwMWM31rHho4PTKJYwK79p
W6bQIg4kp75ZBYI1jsOK7JB8ZNPMkd5Av8GmUmcZnBpGU/k50suMw+G9yfvYuZIeu0chlcBMji0x
WyYGbv4azvupSknvjkiqA13YkdYkhh34nrVhdudj8fSJ0YphoqjCvYGPvrE1HZfHVHpDI3ID4zBC
Atlc4jvYhgBjfUuqHnMCZY1rJ0gl/bo+q/7u+IxshhE0JxgmKjzy0Fw5wG9GiJJfrWIkGSxWpgbn
1lL773tRAx4bYhRb74vnJ32w8gI3kZj4ElqKg98i+c32A2H8wRNyZiQJ31Jl5xmSaS+seZAjxQUb
3+dkTL0/R+8G/wCUrwQyE2h05Q2ooLmIvgAw3OvGCB3DPO6oj2agEIVpwezlIDLABVePvhYcAPRl
lNH78BdzNU2D470vTSWkAYY81Dt75ykGXEVzgHVn3NO6M08btneZ+8xeKLanCaR+LZrJZpkeyBn9
d3YkuFEpbK9sIh031Rs3LE0cOJQhZbrILD62/3FaH13CmIlX62UmeyFLky09PLk7pS0DK5S5cLsu
e0jWgmUefJxRHs0SngETCX4UiSUex06JGscxyMyQfawvbet5Ut8WP7QlDr41UpjcXXMGkKWAaBTw
5xR5hb3zqf6LEFwS3wXqD+FAin44uTJi45fSTYBiyBExZsm0wURQyi1sKhpuGc0qd976Np5apHBB
ak8/mUpnMMbgDTsAYAzxYbBCLDZVuqIZqOv9hMS9gfo1/BDbx+WnvXyyJRd4n/jxNRmc5calrtvE
S8PbfHLzBe2t6yTlE4VJiEqILMW2oF3qFWaGoddPgGPR4xj6ysN/c0Js1s4rdgjKGiROEJmGd52L
pgS25LePczxEoE1qsnaNMnx1AEjCl2CHSeghJs1k0wYnWztldNqzREav8Jx0Kijzm8AwilXpWb4d
j96yV8FFeRH4yspnL5jm1ebfEpH9vnF0+IOCIWOAgFE+Ql0zz/2eDT6YpaQ53u44dqXS9hcXJ/9K
xWykv3exKjvvSw81dsUy69766r8eEQ2UHk80yqf6Gz1S372fO1Y8oE08vWoc2VRIbZE4zEWjoeQS
VA8wrvdAMVb5YX0xOrIusmPVyGvxwPR8lCHkMATssq2cuZZVc1Qu7CPev4c7gs3+69klsZebk1di
tDvDhmE7zJjl1lWNZjOf3H6dGcCs6cMTMNf7nG8rst0mZcU79aK3+eNu51bP1Znkl7802enSNNPE
uyGqH9mZXZmb9SrQOsE870lTUtY+OQSdyIEBkH5z8+1gf7M9h426iKovT+M44nbC9q8AOgE1Rm1N
1m7NiYX8Shoe/HfORhqAxXj3973ijfZ0m77d6pBpvjZ5d/ND4f2vmGDilGAEgUMGIVCb64bGar6t
epcChf9X27HRjow0UgAz4OliCCp85m0mI1e1eK1GFCTCL1+tkUJk/wcBmUAV7X02jeZTntRDM8z+
SJjwvkqnECzbseQ+KFKNt4QM0NC0dyC3s2N906xf0P0alkhHjfRu/ljS5Q7BQxi8UPLSZIYBcE3w
FW21XQhn1o3McX4G7UyYVWp//rABuwPblpf9KeymDbN11DY3hybOARjTZoBxEtth55wTtsfvxS0E
KujSLe8P6hkJD0WTzgLLdsE6lUJ+rOtalFoZyjUoV60svJ5EbbVhV9EZEt3HG3vT/JGvbGive6km
xNp5P2q6v0MraCVuwu/eWp0897GFmV+t29mLUB3E8IvvOJBk90WWLMME05EBy1tFCJEgVfo1FXyi
bDyXhF27cOKYuQut6aNTWLRtlMYHB1b6lJegmFspJKiqrtOpVLB4sJEEsSGsoHvjRQi+KzBlRPV4
KTo24ICIU+nY8IgzvdmXAk3TesZG3HXuYyttOtSziA8eObBAXQFXK1U8NlA/vCvrtjh1jrclzG31
mnglBIabLG9xoJ6o/Wg4zpBZLqkk/vPpgSQp6Jbp7r3GWua/PvStUlk8lm3HjQizqmPK99FWDAdQ
0MUaIcLXZQAHOeyDly7mNdeUJ76WNfOjlr3wZfRDEE+l71VDDvNjxOFeLphKi71whha/UCto3FMt
bbLPIgh32d2Os9WLc/LCl/7eLNP/0EPFvqRcVl7oqdOxMIgAKSucSgxr+7bopgpXNHEN9geaD3vn
X/fAwbEwbNqnqQk1E89hnAzzxELZRvQT9b3sh3RmJtjkSoSKak26pU/Yhtp+p4As/O4UEu0/ARUV
j99WgBJjJgvlN9OkYpagR5zTeMaQlNWRu/75+NL3g8ovKHOZpwnxJf3Bi4+QkZhDA5c/d29/xagj
NmuoLLRNESQqtueiWrcEIoiReDPpPgThKK2OG9qi8yeTKXt8M5U/fpfbb64DIjU38TfP6UcJOGcT
Wro1IVCtyYmPhOOOWF7aBfITCql1uukQ2k2rz1bDmCcdvai7xNXk1QijptNqGjNBsN+Mz/tHG3Xo
ri+BoFZSobTrfQVUc3uX293/KbTaoNc8YnprCLtg57u2sSRWMfzWjG8bi1wHW4MX+Y2Pkhe40FP9
oJ99Gk0bh5wnmy1UJwZmeQjrbyppgclBqJB2Wx3bDgPm+2pzztOasnz4/fogZjXGiZ2GfpN7eDqb
ymjU5/jw4gK0QxIvEt46ES1OPYCSYb05m0xjoE066C9pKZ7OO2lqhy6luIAn5BJbegY96muPMGxz
Pxkz3r9jWY3vut/JBhemZJGu1i3TbUAhshtolL4K2bUC/fGm4VxsHjZZWNFqhxx94G9sdrV07rIn
DJC9MPwGxG0IeeJi6+3d+bqQbPfebDf2EINfrpGJIvk95VLJJPxXsnSs5pOFh5bUhQSC2aU0ZDBw
3XjTJOxV5JuuhOSI2JyhHN/WyMHfLQDaXDzbzHmP41uAR1UgErkwK8nMcYjZCyilDKssynTH3O2p
yaSt6Exip2XvkahSjm7jOc9JM35QOPDuWDbmWc1rcRrGQu8nuQcxOFHD2wJrollxNQLPglJubUAH
xz4jGiBnRUC9O5Vtoklf269SIfsTT8yijVbukGOA3tI00fJV2FQ25DVXhxnYW+YpB4dJHRc2D6CN
CJuP3N+Df45YqL234yINTWyq38whaxid2/z5/SiYgbO5kKDRB0EYT4nLMfKWw5PnP7+dPgWwvV/d
qkG2bZDSdgsfs3vaxTIQni894uXZ7vzQ2WDxz1xilJv61VYp3NwbeJ3Bc9eMKz8kSCg+/OWYrT0i
FKmGMZr0XXpiW4IUrY53ioawcCsCPINxBnDUtRC+MdYJJ0pLqEkBlbXT27ugDpZjR5PlZYZBSpUo
LfBjc9yP/K2npOZfEZT80cVbojP/xIjkvErFxJUAJU0whk5U0hgU5gLvsst73BYaOgwO13B2x3An
yvXr+wJTXyVlo8lKEzvuLDTlg9MLlQDbzcN96Ej2p55d7qycy+/mCwxBKn8yq+BxVxftH3zhy+zn
X7jDHclt7PqkVszraHEl4jDm5toln9hs/d70WQmFuTkhyKt0wX/PVhAb4LxpyjgElpzw+KiZPQO6
zI7oZrvrEL27iLQGL/5FEd/Oc/hk9brSAT8+zJf5j5rHibfZgOaMUlY1Fqs0fTAg5viuoR+bh7fH
gGM8zC36gJ72G60gXMRbTKx9q60yzn9zONYBHz+vIj67KhWrc/7JKXYk+bQEsKdJRT9+dZny3U3W
qIMYxO3ImJ60ckAkCScz4bEEdcxG0MKMbeAv2diaWN/K+4QMTonJggaiynZRvcJW+FoCivrJwt00
gEvwiQ3yJMAIl4pF8CL2o/vEW+YapuNEZuqcvGt5BmlNZlMjFuQxnP2VygaybDYg3iidi7BxbR1V
DmyjR8td6oVqSZdPaVZBrZr3vY/zW4YW3OUwioo5XnsjwHDILIdbvIQZdmXwGLHX0pn0zJI1IkXq
qeOwqwmwZ0E9QPlvJgo6VOh+99jDVMxP/7pwAEcdYOWXGNcglSbjVpgj3jffDeRsjN9kCtqcGZgr
E+sQ7v+cBBQapa2K/OUNpu3jmMU2R1VTsXFr8dnkGy1UW6+em7fRrT+Lx1d6Mvcjw6ybDTPS7VmP
eYeJvJjnGIW0qTeycU15eYRYR8BObmoZYoqicph+Co5DdBVjEIb29OW7upNQ34OIBU9DTtiLeuDi
hrH+PCl4EiT6zQ3oMCyAGoUqQLsW6uHR4/h12FufxdTdQdunYgFxZbicZCtytNkInYfiNtWj/fCh
BLoEVF+oHRfdM2iFUFGWmd32If+l2EBCSAhfLevvvRGAklIwNYzhmVmTiZqZkIyF10Ye62Eh/2xn
L/GvnspQpMxLEoZdcTg4MsqWWw+fnd8KttsY7Y/UbXwkT8zDm6WpMFIg/HTgsqkN1w7/3HuUWfvX
PbHNQbtmJCf0jQe95yl1iAAkHH0jsVVu8facsknFZi4/e8I7uhjNQfLU7iVp9LrVmz5W98aXpX6y
tlk/6ltwH8AvXF0vxbjTF/BtdNGDbhyW4MbdO9ipwCpNoYfTaJuXaNgdYR923ZksoBcwIxgYgwL/
DsE9dAbujiK6ufPx3aqrGWaSXcat3bZxgHGSof12nri7JL8Z4/3Fm7V0qCborG9InJRBlL9JMxOl
HVHJLgSosCCrZ+hbKCwHL2d3tcH7y706levg3xWPZjyHbqMze/HEyQaaUHAreXhzhBvz2Zu7nEb3
YYBmW+BsPlvPbCTA248ThWb3RU7kdekSD3yalaW/6S0XEE7lTe5CZXIaRatUbp5tsU0GVc6PA8Ls
SjE5ru1Pw1jhFVS5QagNmg2wNS6QgvphhBLMwT5Hb5hwUBFnraRFJJjWIcfqueRAuvjkaRnwpvmm
7eN81zyU9gb/dlftcSykIcIpfzfeLNdel5iEcB7JU/Sc+0MvxrLOiPHMbuOa/iZ39e+hCA5K1kwo
VoXcGxpOPR7X+Tu2N6YS5pqD3Tbbq7bDJ/OmFjTfhI1RXGrC3FitC9M6a4K+TnyUB2E3cMba2lOa
UnC1UCQVnJcQwRG5d3uPvf9svEfVK4EoxLrgLW642PP1vlOFqd3Z7MrcY/Qs1rULl3UGRUinaBv/
nQ8OqabvyOfXWSxFoOGICcgVatdK6cM5M+SNQChSM4pvUmbmOxpJPs3hoeUYvZzzg94iRN5Y6kc2
YsWr/wkwzBqDE2/pJQE2LLsTEIF/ffxN3q9v4k+64OLrEv9/QSlgHY8tuWVk0d0wpFdG89hKaffW
2/CK5a3wqdJQM979cVnb8n4eafw0OciZ0Q/u6zb9p3msFB6YifMklA4d8F/ms8EFc/mFKnNLY+ET
xqHNqOZnbC31mehJ4PNF3zTpmFxZEbVX+ILVK5amaRbjWbzeneVaq7fTGudkmU6XyW/Nnfdt4nKa
xOyMBgfV4eC7Yf0pDthexbPsmvvClQWXoITWUESnoqj82EAcNgmNMNuV5eF5g8Yqr0LXtBtRMczn
kclgl4XaZStpCOGH8Me6htc1bpvLFEqgyuKfDvC4LSFS473iTEwwhC9wHf01FNNVqnECVMP3jWW7
tFvv5YIHlhS92yAjIRNgGysaBeoUVaRFo7dgVkxGUDC6LOm+eMwQNyMuxfds5rxjE/6pukP+MVJg
+1dG3meHAsxtWgGQvbtdmkWsRLV8Dr1QIvn1204qv2SJKOen2xt2TZ/K5e2cMHLd0cAOmh/qk0t+
YfzmPPMXv9BhJjnikAfDAuh3GVPHPowhokUCIarUsoKZWUyU2HE7B1C2IAwyH4W/hvxujdOxi1mi
cZLXuS46HiF1qb5uWe+PCP5eaENLKo6JTLhoYFy4uxMwU706lyDiZ4wzCWHOY1z48HmCgMmDY5mc
RhCx4RrKwpMjXoSD5MMFy5vftyUZ6WkVuFBPJ9deddFJaGAwEJOdiZ3M0jKa92UnpORhqQXvr5cs
avNsZYlWn7r0uL+g7fvrhYErGBZ1VdgvjC3Hs627Zuo+KlFXRVhcPSE4QHu/WqZJbY403gL46W9Z
ngDcjrfl/htnmQaHU4EhLmuHxGiXo/WCtAby0hF9Zp1hcuPnxPZ/fU/wAUpWKY/r9OkAuMu2IuSS
Cou+vmTz7vpSg0UTMmCRMtXn56tOlgNcmyIJX5Tn+MO3DhLmEjQrIhfFG6B8qmATetlEY3sm7A9I
JAtmkVZLh1SyGEZlXAFfR7tgkgSchZwquIusta/Mpg8xAmCiGaMmR/ULXL9vsUVsX8EOaI0KnFjv
tibRx/XxzMav4wvIP66fqChTodvo0Cm4nhZ+XBbNPVIo0yb4yzCTaDytzQLZQHFMJH+6hXNWqOJo
GsFwnOh6O/aaVoqixM9MxX6059BkhB6k/LuWaNpyna8xtqK2epOjkqmQ4HxJ1hJb3oq74AmI7yRZ
anPtY2Xe8gNJHxJHkekRlkUCOQ47cv72r1Cgx4QOKofaKbSx7PnUHRsLxudkn3SD+Ok/8hFWhgKN
5Oo4V0hDxfRcGzOlsob622OkzF8wm/3Nd5/D4U2koW/418RWL874SXpLkrWPIBn9SveZNARcTJ+3
E7yG7+qPqgFSECLwo/2tMKjzwILY2OVxblq2/yanIk0GngHntWm9o6+E/0GRzPcseg2aJjfeBj3k
VfDXIg0JKJzt3fRMe1NDtFq6VSlAi/wnKixIyCg+krj+TJY2MtFmNjYVqE40Healkyy7wlTOyX2Z
2HkdAmqwKCurPqZrPAGwInep6P0gHE4x4qTbQIKbaTUXbBED7cBF/A7F38pnVXSqgBIlqMfeyMq0
/f/bilPg5jWRVjthVxBlUJQCCj396j2rQ6OYo7ioYcDRGNcU0IqlKVzBpazZGyZwGDXzi8Lx+ZGD
50/Zd4TkDPQuxs/lqTH5vDCvpOP96eKijKEE5GcuEuXJGk+OdkVXRPUKY0X8z9uZbYJad8j3YeVG
HtWVLNeXEd2i3aVO8tgYyWbQVt+haV/o4uCpHz3tpSGTnbuF/WJtXIdKCqrpYH0Cds+POi8zr/pn
tJBcUjoXi7mdpU8XJMwJthNPbzX6yhWEYGFHGI7cJMSPYfjlcBbYi6hfP/WXncgSZK/w4bgv8SZJ
UStSlwTt5zOqQkbS1c79u8H3odqOrGFss5HQ0QK23gJ5lp9UBqQXtteoTzRsQ4R+PWT48+h6WDhs
e1rEehdTbzyzkr7SfQWsn8i5nxRBAv61Vo1Kg261WF79gFw22pQ1lK+spdIzH5w0Q6e4n3QgGbWW
tHvII2i72FIMINWcVgZkde06EAexbF8CPlTTFYz2JeYAbbIQacORovNiCB8vn7ISoenbcXIkVH8x
rFHVHGzmFCEGfZ7qEkT8sI+CTe5RKo9fKLCJSnjG2l8/R/WUN0sRaxd1mVBwTsMMFmCfQS7Se6xA
sg94a8NMdrCLeIAQCqDy8aDS0rXex4vJc4z6K6c9jzVJkfE87G3L8EA6V3plg4nIPgRr34tKrhlr
/O7UiFYEuMSR16IGnBY8gBmMzIPQVFprHmAxN4Z5FPRq+nFaEB9+n5WxTfeKDeCheoZUfJRysl9B
9v/ctJ2q6qPwvJRVOyTzfO0Mosnqn+BctwLjKK7VoHJFv83Uzu9s3b/knMzAUXNEK7R4WXMBWsmV
k3+9EkokiAy42c8YGcXqjZ3UjhcdG7jsM4g8uyPhmOWnwowFkjQPmIYPk+DVcXEPP0Ehz4j3zfQV
z1vgF7Chgx8qCuCNhihINnZnax/9z2sM7WqqptSLlvjDy7V9O7/NwmNMfg2A3zT3/LCZO9f0cFm1
AunoRt0UaKQq5RToFpF/BfT9WO4xg+6VzShLcJzxrzjeEEtVwd6J9TstbOzdpEg8Fz/XrIZMvrfJ
Qq1aiKR4xR444sh5XJCElbyMln9r9rQBG2P8ry8XB5P5vMStuzLLAgoxsEo0Xjb8BRlEvofPg1LF
f7A+pRHHROM94wKqmeWAdDm+GuEVYznM5r38QBG9ZWtUj3Dq0Onb8LtQ3Qo7kc/xd//H7KvpfG4Q
u5nHVELmPXf+l51serCHiLA4cy7tpDW9GfHoZVlQihc9WKFToo23bhWyKS6r/KIWGGdlmEOvLtXT
B55QJb9RDzhvtRy8hTxr45Q+iHNKRs0kWWXbnrMsqlDLwcCGEP0eOnPv6+RY0+lAo9b+/dNZ8hM0
7aNcZiFIZ1+5W1RXgu++IDsnpHJZ7yrGprRDXrXNO9akwTl6pwR88Qz1hjXT55SAd6wE8cphg/F5
L4yjQLiJ1rrb6IxI0RXggtFzcpX/Z8nD705BeIc/APi4t/06mB67OhUpxJU0ko/avZeFWXqwXD6p
B9+t/e/sWLnTrZ6bQrcoG6c4EQJD1f37OozpusHvP2Z+29NMSms9kT4Qvx+4DxMLVOPCyPIztm9O
8ggv7m+ZggwQ39b64uGtW4scyR28q7K/1MfAAXHN5ce1+A+vep3Gr3irak6pnDY5DBgAkZkt1QPE
Cg8pAUyyG1vcRRAEBBt/CNsvqrfB01937xCJv34Qv6zTFAIc/o5brrFwqqEqEFpT3A9dJZkvEZKl
KQGeE6Xf8iUdrt8lLe7YhUKIPLxAw3k5rTZ0YzBdyjWtU8dNOhY5AlwkeJBKiY1XHoeYCzgyKsQh
TB+a71HHkcI768O48R8RgaJgYtiHIRdlzROloChDJHzR0/HHLwK4hr2hPXBSkMOMaMNAR0Wdl327
LY0YLBGJigBfyD4BfDFzInVje3pVD//Dj2vw6klxUCryPYBKsyTZyw1FzpNEfTNP7O6PDQajmh3l
ALi93adNB5gnVXsP91iILT2pkhYEU6w+DfEpZ2G/3tXF7n8ETR7QLnKGGQCwZYNqiRJuQAV9OyHA
1lVdBJ3XmSNH0c2NbpZ7Rmf2VcdRpbSwUX4IOePlzLQJEiBwMJY/IuAK2Ta22i0vVtgu6uNDrUyP
2JRuUUCaJyQTh1XE/lksc2IGlBndK69OPRmo90iv8gfzoDn4VlL2VYA8eHpAIlbcC3bjWbKTK5Yr
QGmGQp12B1w2IprehY3W5XYzwRN39Et7Hyxwgc24Dj7ltpRN1Yp4JK4swszSzRNanfTCEnGCjNO7
dJhoYrrlF6KE+YDeGBR41bA3N4cYvly78vyqCT3Td8pRfq0Kg5yxOYQBF2Yl+PdtuA6lzwRmtwQ8
qddcWG6TNW8Of8lPiW2kW73BAKtCePw0b9O4O2u0NPyt5DLK3c1X1DJWdUfN14bjypUkwxmS1dLD
z1f098/3ihlp3UAF7OfBMqvhla3O3AenmFFSlIp9v51oKduBGpSDayZAJdOSgl+VqAKd4CWhS+sd
f32OE/49vHw2ttg4t4gvu9SFVsQv8kknwD+wjoGWnAhM6QRZYiMVX+ladOe8Bv9tnEqaN8SFaF/0
eQzvfA/S8Rx+lrgjsBUNS3KrlZiLgqF8LnesVkQzPhWse3xLX53+S6t3VLePF8lGm+oDulufXJCK
7z+7v9ajw4+GLZYNSXuxN7XHh+nvp74pg+J1V3jZvUHjyGMYAG/kq2+VT/a40ErunPLx/qGw95vX
B/RXxe1ifmjsaZqNj2HfeX/1xsp34pwpepDP9lYAv7fffrgDiksiEvg9U0/9yBcCVFP2baoao4M0
RRWXV1xPu762EEeJU3uBFStvFXzcYvsbf/p9kj9ak4OyFRoUQulvzU35BxqqPNc+IWH7zjFLcRjz
XF2l1Nyyh2Acgg1IQtElmXtA2Sp+26R0YK5667zCyHotT3AUsuHfuLZ6vkGjK5OBJbMbfOd/KZgQ
t1IVt0XDnt1fpv1EY14CcdGZW7cn+0LK1PaigPZF8V1XgtoiDAV9Dg55oKexvGlaieV6PspFo4RB
gdDcB7yzqXdK32VogLkgDnbsT0XJDvp5diO03nte4HCcqpm1i13Um0f3+T56vNDHWXKgrmJEgfOs
fqCbAhJIOp7j3pGAgWINcGdNv8u3dJfUDlN7URuAESia1iu23bjlE/0k7HBg2HI6JjXoFrfxVi4h
7h2kZOc1ShzVbp05hQSJP27O2PStAcof2ITheDYtfTnlZy/RRDVWrAmpMMyUHzfDTDCPVBc2zbEH
N/OLcz3l5/EK1UcLb9bU37z/Z2jQvv5SfdmBF44vFe5iHruaw5qmUeXtzooRDYVJl9s6mzoxQi5K
00RNeYfccpV3Tr0tRW8r4X0AAqTcNLPFYAw9L89PSWuyxtM/e1f6oNEvQQ0lNJ5U7+BrQdKnBUkH
QW89YpsVXgUJl2wYZ8O5Aj6sVkObB1K7tGFV/x2n9p1FyP1lGP1TV2WRLaON4Iuiq3/2hFizjsw7
uIA5XyINZlAhaO7yJx1LKzeqRRJ+BVTd6txFjnRNZjQO1FMEGQ3E9DXdvLZiNgD8nv0Rhx8CnWup
oaeCEim8dyo6L/9fBMsNUvf5sQkpTk5ygzD/vbbMiqn/ipGQslDqWkjFAKhS40n/TicJ9hhD8AY1
eYeNYRgB2n3/XprpE5qoAvYTmGfTKlcL6qjFQVDagaQZS0gggHvJN0rVuuFjP00R6SgKs5BgWkmn
PEO09CeoX0iZqzo3pIRn5tEkkAWJPFpOTsAbZo2g75gXNITDaO0wM6lENKAF4x8i2XUaHEmm9qwR
sjzj3qtgNusIycTbhJh4sKOSGPNtQDp4HjsN0cYVOB0CjWnNsn9GJsiYsZGkj6COL6GNmq31ffjJ
v8y7MIDD85L6nqkxM5QIDf6LxVfB4R/SXiHG+2itGTF0fLugkB67mX0Nt3uCrlbxxWT4irhgBdLY
5xg9vcG4B+IF/nf7ZpUMGMCExBn0BxIMRnkDC9QG8JqInOuMQGLZqSL3tWy8hPWwZUcmOKdPsTpr
N9VwKMK6B6dK05QJV2UCHZv8Y2lS2tD1u1gOGes1HQ4Xpv6y7jQxQlvWXYvDAN1HIUbMMxrZ9s0M
uaq+HVgP6Ql4i248tpf8JSMk3Ys7IlVAIkqDx3Y35J0/0h9SNSvMVfjbdi02xgfBK+yyg2KI37T2
COXOgc9Py4OW+yhz0N8QUl7MVg5wJ5e770mcbqu0CBir+b5wWHr0hf3rEuqd1nMbbfTZ8zu7koix
5NdfuGzUsvZrKrxCMidB/IXxXBTAnI1hWbtTXZEGvH//GVMVNJXaUj9ydj/p/814Hn/daia5+n1z
+6AK0zxxHTGmV+s1myKaoSC38r8H+ye26y+9bDbM//rtnuXx7GpqJNu0JXsyNKUFvyRKkLUsyFFY
7UWeK0qUqig9afqMlBS+freyEgBPT/Y3Na1QFf35D1dVlbgAB7Ug1XmjmzObCe/S0gK+Sq+FUQ9Y
sLHKptSMtWvMV1MhWb5ZVzczjPQgr6WLncimQHXeyG/U8RHb9VAQ6KDhvQxZNNFDXbMSKyOrM3k2
Z12Sw1YOQ2Zf9OpywZXW2KbPICWxjil86qFUhV3G2DWA1w/7cPjKWz5S/KW7+OVLxN61BwgV7mNF
Vk93CC61XAMiwZr5DmeGAd9Grk2KF/KezO+Ph3eWHsM+8HEpbrQIJ1tu0VTQvIv2R+CizmWcJfTr
IlRiINgLdu9FOqTQzkkFtvs+d+oqIfYuzI5ZJUwoNSogV1lALwQBRnQ4wdy3Eu6fOrnL0RdXg9f8
4VtEOH4VLMA8NB14DYnwcpSX/f8llb9CV6fXLPzSifoI3C8WeXyIAD1cJyqAJFP5r+eFO3THpEB/
5gY+kbyvSdkKLrfQbq9c16fDvxF3xC2QgQSaYOC9V0jf2C2pdZa+3xhDri1sImpgrqFxehyKiT6l
xaays0LLwP4+YCgKB2GwndvZm2fMpan0qJh5ztz+pN/CVfHTfe1fSizHoFVi7vEVf8BUA/muINDv
gyTaqO1pxujWFSk3Q66B4mnGnu3pHl482BMLLANMMkN5bqid2wyGDEWlaSsE09E+XD8GWVRPu7S0
Wtn4TKrXybi8bKm5y3l/tbpXzg6U40/AdNEjfY+M4aDAeSAFkfYgNIB7eQrMEzphiIIv19+3WhdM
NrxU0hlyPHfuvCfk/L6ox7YijoT6DniOlE/bY63CJJtB2/95/M/rEDqPPKdkQ1dPpVIrRDVDr9PJ
o4/+EY9Wpl0xlCYEs2mo+bd7NolF1DFYMiOu6FiQ61aOIJLzgMeS5VHYRlihWaxFo2u+e58g7yuX
IEQgJZKg+LuSekwfMq+LQNckUGw1XvcqzOd8IoC0j8lMxLN2bjzs46ozQFTTeY2cOKp6/6tHDHZZ
sKBblN0VtWuKalLX/GUu9a4Fok5AfjABQKkzQrOkacSeqvFnHv0479Ctu5y3yasCBl3PCGTBjijW
AWY/dBLsRDjXcNJuPlD5t1bisr2qM75JLgRrYJbWVt39AsioXWApk8frc1BwuYE4jFAC8M9dclyt
FGVa5p11BzdhYxuhj/FNsvSiT0X2a7iYb49WMsmdtSc+aIp+TJChXqgiRjmBEWzhyIpHZShn3yxp
DVl25DeTd+zPhEmuvWrZH4ADQJvWwm/rp3xMH94eoDBF+kznjsSRxRjuFtjAyVggvAImdRc7NDcr
3J5IhbnK5kC6ZhATJ4KZlg2o16ie/h4+j/1ZZQnUe4hJp4ZtmfmTo1qKJDd6NO7M6/l2jD4suhzL
DNYHFRIsyFa/v04CyhtUKZGH5dWZ6YlJIpBz6N/4cn0lojQ+U3HM/PPqwSOPwZDAanGNzNTz8dAH
7CAPxKP8YYNaPD85uvZ6oy8cBpTGGqT6U9+IKQvuTGko+cozEdCp1pMwR6RBfnoqvzqxqO6txvmN
CONpYTqQPImqojgQGL0Ye/POH3ghgqTPE2ya5aWjmCVcB6F43/C0Tzzi16kYPUwH/g+yqX2QZBFG
j4ul7qFuuxqkfpth/cau0KmnN515Df6njkMGZ3YWDsbonoPcZFcbcSMrxQoIMAZpbpIj4JsyrgP1
QgYbvQQxcEPa4CSkMRa51n/DvJaDdWPomra70U3uEPLIHBWaPFHRL1Vp82+aPSG1SVJOHDTVVbHZ
ljEODQphVwqV1O4yC2eB4nzFq1sBbFuhP+wo2upvP7l9I9VC3cFdTflEP+oL/k2GBcuzYY/bJ/R/
q6kSZKm/xBI2TYqizw3M8Vp3AyS0gQ/FnkZfdXNUI5HVC8y+yW6qb2mfsZI9y/b9+HRcBekFKjxC
GTkGOEJ2w6UrVvoqGJOstMoJ8hEf5lNuXSR2XJOkCI/eUli5LBH3Bv+QFDMmYmHHxmvU+neVSUWg
vQcZSjSb5p31rAm8ydxJbFpbj9rCugt9wik0wulkESkVPj7rlHIrgf2MvzmWeE/kXwatK7Wy031E
KWdzLquAxsvVG1ig1/ivVSz8eXeKmCbAj2wg5UxxsuIfJMDD/iYNSMLHq/DXT4KG/RsXfZ6bVyVF
rHldNjQrNPWv+4ISwpjnuCWMetUnJPLHZ3yJKn56+FAPJBZb8E5QYf2mN2Skr9BDNVIidpALjTp8
fV/LWbVyAiFE1ZCUyKULCS2WsF6eoVa78tQBHTUxuavhiC+Ip1yOgSw7uRX5Gf5MweZAPwjML0lz
KP8+fa52unpC5vsVspkghxnw2GMmjBYYPF4eHV/Rdt6NExENwkHhi2iYbMZy45yR+GMvdH2GvfEh
2wr4IHKJNxWGRb/gAYuoBKUQLDBQCmBlohyyEvP2cqyhARqZ5cnKgofuR/SgGNSQa2pjbRgbwzgh
/6no5dzcOYzNiO2MumOTTGx0to3kZxQ/CUv6BCJfnFpam1cZxUN/SUCM+EvDv4KprWlZ6y2+lIty
X5YzdwD9PvZMRWM3y8sWMCyPUfvt+8A24HxEzDP6CJIkFsKaeId+9i7Xy0GKQfqLUZhkr2l3XPqO
e7ZFRr9lmKIiI1CfANLEoF+57hXct2i+BqZDBWRbouiyDLDS+O3VyubPnOW/pZ48gt7+GNaD36vC
9YODRYJ6C8BYec3h8cHxloD3ydvZkUbNxNLSbEEFaOM+ccp7HEDiupUuVAkD+yMsXHl3/Rt9DJiw
pGFrpA2XM5qwHbg0xZ9dYcnNoSZWmqFHR+2sdYkMuy/V+9nwTeBMGvsilq76q2stP6VN28eNC03S
CP0zM2FFpFotAshC553/aWDomNIUiLjIa5UA74+TT5Q0jCUiqNXwuWb1QowdygaOmJp4LQwHDBGZ
Ldovox5mLqIMfDzJm0uG3saCUf4XwcWiTu/Q5MGZk+nlcX4S6tZCfENTaTfmKC7FZiMHec9hysJk
r/tDTB8seQB9K/+daWXh9d9Kw9FkLbQMXhQxiioTQIg1bB3xFmhdbkxQHNhOmbCTPf8NPif2KWmY
eFjkzR+D6TuXyy2Qh1cQikZn2Gttabc6YA/Hb24GQLM1qhLbiJQ4LwPA7dgxBtfM7I9IttaKnqED
51ybhwcsXH06ul5TgxhJpDaiQSH20p6Xw7/M0k5jwuZX87nt7j50Phv3ILyxyze6dfHg8hsQPGQ5
x6+m9ue+nxBuklLz3dcpJYnX2VFKqli2Hdx6IsHvNSYLlRlb1exd1QadjgNOHN3HUXgJTKvBIgZF
iF14h+KbGiKkA7/h508VERQ6UyuvbPc6xxsSKJE/b0j9XjL3ixBcWRXgyVj1gey/GIGK1KcfxWyP
0LR4sGL47FOkTxbiKh/ZumhNGmRYoYBqaYWk+Tb0kQTzCWmdhUre8prZeTjN6kYVhvEpaYEF15uq
jNRv3wFMyC2x4tHKLzhhHIqBSEIRKN1c3FIS8q0yIPe0GAIuBnos7z6EyLgRBakusiayvf6VZkdX
ncwrxEFtHGcRvhn8Z8s84C/GMzemaMjDwrXVkN7Y/m9UHYdYq6hpXZZz/E6xu9cyn4v26OsFMiLJ
OChAtMjxMIcISWOTOATG4tYfIHLBDOrcQi38+h1hG4tCcH6172ZkcfbKIGB1N8Ur8DMf+oviu7oI
+4s1/KvhR95dO2lgeT2TPBL6WMHocIHrqJxDkSZdmlqoUgBfEDCtXJgglrw64GIbtWvvH1OMEFn+
0lh5qNCipzAB/pfD5UeieuInD72qeKrIFJKoJFZb4+bbb0s1uZSJAz2DA7GqYFIwy7ZOhCiA4wVu
dwurg1qAHj4OX1dKlbxG+FP7dM9PoJOY9fRDKf8uPVj+j46euZ7woI1FjZCXb25hhF4HeYT9zy0x
XSHeasJ8DmcSR8NcvxIwslyR8f/Tz50pwsfdyWQXDOCbbtSJ4F2sUkxmMhIapckTBamGpSZ7LrsM
r1Eio5Yj5+iRAc9Vx6pb1ASRuFu3jz6KmPDSqhuRd5FwYF8iYs/Ylk/FX1BJAETWTsEqvPyCJWl3
Dsl+TbtaYS/89/zL48yL8POzF2riGMNSy/7nPAH/3SRF4F/vynbbmxzVXtKFEGQAuhuKR3qsNIPe
LADDKao8idA7L0TLXJK6AeO90ADLc153BC59NBz4/jaT9LdzFSMezMEhS7AUgjP2m7OioiTMiEGA
v5L4J+F9s3kpoGWdJe9MCeWkfJHqx1VYnRwENvnxlxuIPpQ8k+hdevdwmRC7Aigr4BoHA3VGb09k
gQQS31qa+51vRRnxx3u9Ks9mBLZ0bV+cZHCACeIAjmVOtaowkfd29EGkr5fJURSSLiLkUHYgTxZt
JlMIpQI/kxmksJoSVv6VZdgzR0+TAZDcbciZrai7PB+oT0tsOSKnD8ZXYurZ2RuzsdLylitcsCzI
BCztUidIVbgK+bAPf4NRhw2cRmI+ysIgxpvc150E45eMgOya7Lczg1dRvRWYDLVqZNIM3oIlTYow
kfdD060JWb5czr6Lax/V7TCRTzlB0+e/I65vh9w41gapRqicf2hoFabybefP/zJZCUDkETO3EZxm
69MtMJx/I8NsEgYHCYol23LrFr/16OmcNbsy1Lj3Z6trVYikw60rh0vrjxUs7muQsGFQymBVMNzw
wEXVLg0bEXWPlK1wc+Y91mr4ynheU606QEjm5t1FTBctWIei7PYaecSF4kXfTbc5JUmdMLGH+Mbl
A9ZG18u/6Qhj7D0IP4Dv9t7VJ+szARBwdA9MMSkTx+DRuy/nXKiXtPEhi5WZUiA17IZL6mb5jfQk
jlH//iq3ih/YO1fMnSZRiZ+fr73oxtURSwfe1dUCZv3fH1BIvRpOsPZBi/w+jl+wZfSePoKadxBP
0A8pImcHX3ZWSOLqLXh0IW04G08CTz1RTAQI0xXGZAkiUf+EEjS+F1HJdr6SDP7akngSQ6tADcjG
LQ2mlSan4i6w4a0rKOWCLPWvKWWmx1xzA8U/hoMgFCjH2I8vsWiPoUSIiUl16ZdVz/tFaHphrdt0
of25rje5IQNV4+H4ZHVJ8G3BbN1AW9WoQG6oSQKa92pS3gKuTHcU+s7NhpzMpwroacj9vMQv9Acx
82m7zkBWyZqsHNL0VSUGV21ZH6KKV5ig/0eEqzIq1eSc7HUeW8UIqadk/s6HjW8EezjCiOVj/ZD+
Y2+6yhztA+xBk2eADxRwzOjortYvEFtHurM5kB2hRYeJBZuirl4hah6W8X54R6uGQqz6BgQLCN8M
Fgo4GZ4OEWO1XlGItMi75eCy9uqocb96ZZeaOnPCq1nS4iaAMmsz1Njz+6f4+TH1Tg9rr6tbJjkv
YjfSJJg+JzSNiQPTdt9ioLa0NSubCUgjHBb1EGFemiICQOsPYgWFSJQ43iV+fa/HWbxs6lvNPlvd
Rxs+uGTxOK/vHqC7/z1FC3hJdfQCPHO3zMlGfax6jzh2nFl1jjb/HMGRuyjWI1huj/ht3L1g8+P0
aRVDJRmYvO1QKEG26kEUU4k8noCnGXoG+1pgNceI46vM8Vfq4/Vb2QLJPqBA8KcZsL66hUJPgl41
Lfc8j1TRphLc8yV8aNf1x5WZAFp9GPZPneIMjlyWKrcF83cG2vER6c/4dtQfJ8s1yX4H4bvpHycH
pKFAQdRiSrMqBnbyjzT4/jY3yzErnQq+VAJWQFbNkKTCTaS4XFSVWmxd0tEaGFYelIcB3OQy8+Jx
3vNIHwL8SBnMTkxqF/rja0ZIJO3qDbWC0lRUgmvQxYKt0XdBv0PaPoc18L8x3+BiLY8Eo0O1K4ol
AFv8fJ6mcfVrekrG9T3IWtHIwQ5rjHLle/P+ELqNmfyee1wLBf5r1Hlhiia7k8ClfhwLzaNuIvvB
CBsUCPXVAnUdv32necczvdb2TJi0KBZI1TF8SjEg0VXguTBSdvpxkCwUgBAJnaQZju7w5whiDcMK
STwSt1vBDtO5io/VPK6z5Bi0oKTo9Lo5fz7AJ28Bkb9GELCYVe9CxL51NT2cDPXujMNefFD/POH3
jd4WeIDYeKiB4B+9c4RE2Sj4tjY0+2Z3vBkkVKP3nJqjzN6PtdVsuTyUkyL39MSTsQzqu10CTmOD
NsvY13m+i3nKZ0gmI/1JInGmwelpndXbYivFwybfsVDEhFURxdx2MsNqcCgcYkVX3x+2eIq2oqH7
frxtIz7lCQkFgfrjHOHzhTjx2M3/+jYuJOinfwUFeI4/gWlZvsiPLenfXuP8F3P0JcF4Hcn6UJtG
NYZPKxneNSqfdUnhHoJBc0jIPGu/lUPDlz5z4vcawehMw6LStyKRusn5nuYrMtK/+W4U/JuvlSZv
twpX+CrJQddIM6vBPNJxtGjqsO6CkqCc8sjp0DPQODWinnxfpHrDEU4l6rUH2qLDKAJLA2TwIW4z
3DtJQ3e5jrYdcliSpXgODecXMYbdaPjBHdq0XO+lrQAJa0gM01wa0xrdTOeVH7Z0Tku+S1/ft6wd
hUaPLzNTW76ORlSVOGm8slGx0NJn/LlBtV64MlkpBU1kUd1ZXMJUB/Fh3m6YiiSH/iCFmSpj97p/
Bbd8hn9egwU+AgSzPCduFHBOOcDlCWOmWSGOd9KN/ivXOtr5XEM+A2+IFGT97kfo3Dbu9mH6FKT9
erArbE+N/lCKLy5Cnu2mV7XpzL47l0ob7GDycBObL3zZnf6uQrGYQ5/G1XxwDWvl+VdwRqXGzMaC
bAo0pClwjw+EfqsD7N50+OHMEuCZr20duNlXzJdZFPSFqV8I4gQprnjJ3NZFVJOyfpogRhVYDh+6
ZT/XvDw99jMRY7QdTOE/S9DFtxwNGJVpsuZMIa96Ap+62efAsiaRnCdCk0B8zb2M0E8Y2UH1wxdm
ukX90Qwu3xtP2LvAR5GGF5KdMi/wdPGWx/luXU4sDEDqeYmnSNBfNFM3PLQ9dHMpVyqsXp/Ip2QN
XHgrd+U+NudSXlitvs31EmnjrYDgiTVfdGcRFQSrUmMmojPIXTGQbIYX4x08Tm1Sr0Pe/AEihy/m
tqBZKMxISyU7lF7x7E9/8c5Sqa3ZGF61I4keTeFCAvZvUkjrbWLd/eZ3s1GM9JbzOQ1yPU6ptsQe
o4OVQVkQoY/He4PNZVE3nitUlwakHVWe9o5FPCPGINJ4SaacHpTxatOUvZdpidrVZzyHUqm/2Hdy
yKodzvMyLuX1futr4PncSVXl9Jeo4AkbzCpoQDb8r8Eeoq3+R5Vw1nw0gZ3jJPs5UpiIlNP4gTAr
0YhBMgCkFCgYdzzhquEU2iRZj/lWvAS3PCFm001uZLJFSKtsbpQhyEODpx8fe2/73ej7FkifsnB7
W0YH6Uj7HZxLJmG6yW0+JE3j71NKjtQ/zJZGoij+DszIonJqFkAWPHK/wJEI6NCMioNmi1a7sq0W
Lwlt7tHaOW6zVevs6DSaKACaSY0nVCZvQPZaoH4i9W2hRgccLW2cKYCU7dvVkRvOCWF6lnvxTgMR
WoDi9SV3RXMo+3fGZfyaO8PJiefa/LuPkoUxujuLJPJcPaDT7L6m8OQT4UnMyDh79kOEZBxNfNn7
ewVn9kmcBCx+ePn6fEQNc4tUu/MDBD/VKqEz87LqvFhCd9IXMctampL5DOClMmgy2BC62wT3FUAd
oFuiunjfC3OxkiMGJSp242fcm1f2RMTQIrcyEB9nvuozdNrxr65EVtOl0g77/+WxT1SPeoC1CyF4
3ERMwv5lglx9Kv6gO1It0EYKaPad84EDOg5we98jG8livBCmupwSiYaDf0CZ8haSb/Fm2F71+JF2
B8Yk+z/f0AnigdXc82lXlur3MUEFnVMZ1+UFrVqZxAlMUV1Fckp/R06aVFXJPEosVAPohop8bp/y
gopSp9ea7ywQLRSPDYji5aH6C5N8JqsetTq7B8LwmmO6V/xZznGqRDmesMpdDyfujxgzec46T2oj
c2ldJwwoV7JaNbRImqnSdnxI8P32n1ztpm737TD0jM1Y0bJ1rxdfUPJSikHz2IPGkfSLatSrzHU5
XC2BJ5UnqMwe6gV9SPNlQMjALcRutDyMEVmE3ne03+NlKW9Ke0Aasl6WpJLCnUl6LiXU4VfsXAZA
jiIqISvzT+SmY27zgIHfCc4JxCwo7gvtUUX5vB7+t7vQAuIe8i8yOJ4Vx4pIuNfjQ5d9w7sCxkye
ZoiU31Ul6S7Ucp7JeLBjXXuZtB25TkVdgGSz75Ds27mSErvC0xS13LNpqgm+ualBysAthpbiTQVf
vjHsTQV7dFfkF7d6OqRNnKSI9cdgQzNVfVm6nj61thjl22ibeZ0IR60PDtADKvbXJFIcbO1NV/gM
IMeTQOWC+eCBZsKim3PqNw2lKEUh5uZ9ZdHLKs0gWqz1/99s6GnSAghqbO4fjCJiEqHV8H1K1Bvp
MA+7zXAlk2BoxWAu/r6tuzjd3miouQylNi3gHhEu/1QIQY+x4dIxgeh4idThqbgNIfhyMzyS8XD9
y8NrLiV2XHN0A48/y+A72g48Aoea73co22ji+b3+HOZ9ACqpILGKQGe3ZveRfzKNi8k+X6mcV9v3
GvvgITd/0tB3v1X93I+yKeCngiwuhkg1DjB2i7+stiZ+HA+TxEQFSn1jyAFxAzbvIo5uWT5dICKE
mijCsvxEh93okoa+jMhuDRxi4MprmdsbrXD28+7eHIjWeZc2o0FMCRdWyyYxFwBzQKtoQc/S8W1x
ykw6OxpIJZLdHBbOdB9MetqkPPQjEdzldf/WlBtIBU7ipNyudp9YVBbvA4eqOawMzPTz3yEU1LHQ
9aUZZYLUceyusnROaAEJif8oe1HA1men/sIgVmeqQYEAHyaDi4dLv5SosIxnPdYJfdXXExlo08yR
xqe1KtwE5b5ieeGY2L/wq/uCyBxSF8dKQicFxtx10iwzDiU1i0rApxXiQ/d2OAaepKU6u8whua8C
LR1XMNxkuhEy2YwCgjV8Zqs0orzK58RRnfek8FkjzAqBd53YSXm8ofHAXMIndcPHmd3JdK6QLE+p
eqMy64Ae2LYsu9H/+w8WevIA/nMhJcKsCX4pBNP/P6arkdkawwDDu4MtRKoO38cCKugtFSHRFjmT
jgYo6GksCRGgyNkN3sQgLRYTilA5PGN7qz+ZANy+3FIbKJ6XGn0pkUU1+OoBPJngp0lKogB3ybKI
OfldxGurhojA7vovYY5y9sIDuaYlTocme4bJT5nklW2K6OqozwqhMG3klO3GW/JoPimcAeAEjKoX
N8iLhQRne5cqb0EtvSzVcVdB3jAxO63f0YLgTqtZNQA6Ecbo/ewsuJ7pHuldaAJfQx8Ho3B8a2Oz
eQhkywyKFP3VOBPFJS+5+M1osRRr5eVYZNxT+5S1Cgu5Jj18TkE57lS/YG/AXk7SxeTSaPeeikoQ
yD4QM5YUEsfTjOEBkQzKchtEz3lQv00T/fijgFwiy8QFcu6jqhFD3PyEqUcM30XlLRSevfBrl/SR
0uIGQlcjW60vALetaDvep1hSFdOWJS2cnvs1QLUoORiGqV1EW5ord6qIlGgciVqm9UMaK1oEhDVw
Zv2cCUMxmQZdYv5l+/SDsR2cODppQmlIff7pYhe9708RIXjFqnfMTZ35MirakAwEiU/TRINk0dEN
JGm2ZbMVgTErn98431CbSSZcgzmDhSJlZnfnHZE0vS6ncdXbf6MIkY4os5WYKIAUCPrfr4kIgpwy
8jCIkcsZjJTyVmEYIm/2uJxU46VdoFKDhAezF7i8FFXpUR0WQGkuRQ3th3Pn8r4VPNW+TPTb+ISS
BdY/0JIoWVUF+i8dcrkEqPd/N9h7LGNEfaQKZnLWZ63k1f/UkUzCue/9s57MBM6/iuVWzyTSd48t
h+Zzqt6heXg+erbDPdQOQ/lxC14BVbEHWQxTqX4pAHnIDbknHK2FUJ04XDyAqHwekzXkWSoSpHv7
6x0gP2xSGCuBj7SIXKM+mwhuRRpWq/FZsj9a95l57kdda6IHC4QSrnfbZt/qK4p07HCIVh/1N+JK
haIYYdKd9sS1WfCATJ3OC6mjICe8VOfRp5Cye49WDIRqqV5kyUYqgYnz0jGWGaCo23WxUgm+uGZy
2P3PbHeQYtp5d/Lfbh/8hpiCh1+Ckg8mr9Pwg9zJrY7+DQC1JF41sp+ahzFxcE0qTCEgNmHDRsIc
Sgwb5lpAvAEsQAohhaHk6JGnWHdSQfOgAja9t3oQ9z9cMIR58ocjV2XwpAE9pipx11a7ci00AshD
Fz5Lg8QDKlgzbu3GHSbn1sO0rwHUSj0VWYxqb2hc2OSuEeYQSq1MnJxT5fyZBmCWhUC9F/hvZvoD
SaWZVljhs5vYXBx5VclpUf0ZuqoiTujDZoTIuqIP2acp/p/ScfW/ZTi6PDvYRCQ0LDQhikbWXyvE
7yBIkoRosL1SSVroGmEYOZdehIprdL7Q56WEL8cUxmWmAhRhskHJ+FIxYEtuAOWh3jxQckozKhEu
zHPreQpDSR7IImsqa1zReDSGBmWw7PKBdgvQPxM78blrjOCt4drnBTj5tda5D72pGpCfTJ9+UKEb
KOQxP9QFTIctcxiu2LfVnKYXp41D7qqoOR7yMDb4LaNWu4Rt4+wNJzeCvMrdXt4SDpT9pcqYBnW1
R2JeJdj5hGCzEWjmz57fZkSn4krpQorkcPZV1jwojXV6ulT+e2xEvKMQJGfIKxOvjPlyiW6DdzWu
9xezr9A6MvR81UU1NXbLCM3XtgZuxv8U51LcaYFxnBKXC8s2cLycTtv5b/MzT7SI2sQzXjvTtSUj
PSuWKjJYqhn2s5QW7oB+pujjdOn332IYzL5MakfeFw1MGLYcR3hTmpyt5xYiUS+Rt+DYqrE6H6fi
W8ZbdnKprf5NZSMBw96kgLTKPhGRTcbnJRmfFEFSUCQDlyq8f0OZNaa3N29nhH/gu8bGzqAxaJqP
EYye9Supmh+psk30tICsz6qwCa/PSKSaf9LQvVCspqCFa32RkYb3Nq2OpAPHc2je4OLVLwEh/YLw
hytFWxh8idnHJRMYx45V7o9L9fUIYmAQWVgVYdyXGCwPu3OiBbvcMMC9piIofaBlALNnsb3R+GW6
o+MeRKIIO3ghJRs53f2MBV1mgjXH1jADGp+ZZriFrmMdBFu+auD6piLdkyHelF3IXBolyxjLkeBX
oYmRW8XZOTyFWbOAdmETDNLQwH2owqFeZhCTZFzqPqbU0w59lvgAMAjpVswHcKB8oUZU69nGV0Xy
fMwu6hI24SnbD3ZWpIX2rLu8UO/S0gC74wojZWMDUWmcQyTC4yaEJrknmvdAux/c8b7B1BTVAr3+
YPdOfaSTi15ac5GVabqn2dyWmSF9dxoJ7O+Wh52eaQCKo0PW2Gii646G92cxAdj8wE+wxbPvYsyN
YINii5KOdSSzl2+UYjy3NWyVlFnT4Q0mRf/Xd81PlfqvKlznZ7fNm61hHpniEYz9h6uDvtF+Dox6
IINC0w1erB/gsaXZ9I78XTWWUZ42I1XSP2lYM7PCNrN57XEj33Y8gPdpZGu1piBoYCRRyTjxM7l7
EqfkEq3IGKK9ybODWfs5GyNlocJbgzWwh8UvvCWU0My4TESpYkWzxiOM2lMamkVPOrvJDEjFfGZg
OIUeJj6DoJeW8V2WV1sa7Wnxu/Ws/DV15YD9UrlMhK1mi+8XjTikbsjrmcs7xGCXeAO5erUruFtg
TDjKhd7XEs4Eeh0XVZr1py81bGgRdBtr4vePDP1tIsv0rQbY/Gb4KL2OxyaDZCm6kch/O/9E4qsV
kF4dX6E8qGBM3Y1zVqi/KDtSTmERxsfLxt3INOtAuScKhQgZtczUR2bUkxuYxmO7d+EpDVkQjl/v
aDQLOMz8r40Nrm2ClqYcUjtHBoyhkDVQQF7wa8wYECTE2Il1ZHVqaBpaY4qbzRYl6LkBAOWR4t4r
SpArfqqMc1Lhko/RyaEFrX4ZWW7e1sf5yAxEocbW5lqhQwGfBzQRlkfHNNR30/SXfVbtGIcvpp7J
FXeT4ZdaJ3aEQLQyEzFAF1fB8XjH0S9S4/IjyhosAv6GDLBmbBw3jp7SkGaZ+pKx471SSFHmSikt
BmbOiPUFpLNxD5znA31HMdnHkCN05OMx6o8khr9jusO+s4x+kOpa3OfA5TcaO3VSmYKPoRPnmTyY
SCWrkJPFxyZwvMa+3Sn0MJfxlGtpYz8KsXcz00jHBEGuhalg2Qu4EnvUMFhPwIkDKS0w08IDQwLV
SJYdfO20xmumD6HBSmEx+ItLXbFRIRDiZZbJsoqd41cxwWKtWFrqMC4zKMncfZ/QOslO0KyrPyiB
osY2yemWtd+kCqVJoEns1dNPiMORt7v9iVFvKjmaibgX8bRzXpoW+dgCkQUmqPuRixDk3aX8nQOL
ebl2vBTcn8o3h5b8Th7Xkuy7PoLzi3siDeI15KykTRySp2T+qfiHNEB9rrIVwzXtdcQvfQJAitb3
uy6cXLn6PbBZ3Wqr15kJvDF6lyTbxK6di6BsauzLYW/Er0Pqk6X8Wx6QpviQfQK41Ulk6Ii5U8NA
ZqRmjjWoy6/EfzNturMSEM8vPmanli2zt4Mq9fyzW+OdGwP4gjmPA8kRX9VnbuUG84VcQzeHHQd0
RDd0wfKDzrBGWypNFdOlBNAk+CmxNBoWVPOiPGjXFD6muhNdQFuWPwXzBOI3LOn2yVsJTm8o3bYd
PKnC69vtInuh5/cVoG0vF+ST1lH2Beohon5O0+9Qa+u46IGZSu+n4PDq2Yec4shKg3o0QFHpkmI2
4c/YXC4/JXaEvGICYV/6FR6l0b+IgGSg7KW3nVYVNpUNsEV9s3bINih5Gmcl03cK2OMGF16Z4s0P
Bx2yOT0JRPd1HGRvoYt8Ncp6G7mwSQ79Qgw4NZEKxzK0IKuarVqFDKNygbS+ExM43mxsX1w3jRu3
R63o/vZ1NfWg7r8YW8/IR4U1NUifQeTfkRkYrDlHDeeiqMuK6hU39k+T9TBUDWblMvk9oDaowMq5
DwVEvcAAOAyGrC8qncfjP/T6+Z+Jqy+IpfG44TJ1wOpGcsXBfBo6mASdWV9TllSYMWWia7k4IefK
zUuP8VvrD8grsw2bzfrrUGtsYxamSjkaEL4WhuePSuINqfuWqJL5PiOwR0Zl7uaDFrPJ0eA6R8Zq
TIWACGIOpvRvMGmDbLBW6vyqFFNXGNcvu1HQE16uMoOZ9KG2IV449NipiWWgVHGgZLqy6M+j8cA/
6vpVDsAd14rn7CXIdbrItWU1rWPrA81SXBU6JDr7U/u6FyOhOqc+WMKKZ0phEpFmssYp7sOdqTbt
P2LVwDSjze6fOeyzAZSJsvlukSqFn4YwblGZO8H+7BrAYTSGP4X+N9TlHpHbChypWHKZii0c2fOO
l883NosEwBHlEC02Qvwr4U6PTwkL7/kOmRaPJ9W4ICbylqKfOxXeP/Ju/WQTgz9tww6NuAxG8EhI
SiviXobZPItjX0nvzfFd3aNuM29kuUM8++OSk0H4ODQm+62GF5Yf8OudqyvDhN3j6UzfjzdeD3k6
YxvxhQQm3RG/1EUZkdaBh/lsFTUfDymhDH1lnGNKB93jBt8tHQa7FB2FOKlribCiKRaePQLPjxX9
d507Y4RoICf0ZCeyHkzUHj8v/VysML7UmpFSj+X4jVLM4VbShfVkfIzd6mAGuXnN+qZjnNqRytdn
1V019gY7NHhobDJo5qglfsN8OlC9edV9XT7jU4onfyfTRSXrO+kYjI5o0vtzcExLlZoaSQbVrU9O
fnjHJL5h6sCm2JveJ9k0H7hKIK5dW0e+q2W+GyiRCBK/EjYAesD0gd4eNUNZ9zJkjUUhITMxvkhu
RcQvrfHTgPmiG4vA2SuhE0opZkFmZyQxf45Y9XEx4XTD/JNPuhgOco/V+BE3yvtwRghOyrn2O2yE
gAlftg7aEaOVBGZdF4ETuRa64dYno8/jhdBN8n2cdqHrYui/hnixppRpQ2y34sekbrRdQOq0CCVk
uv0FTms9m3EQ5IBqlDeEiml9OdF+ZKSLd89AtTLLqY86gB0YvxbwwaBK9xHQYUFBmd3wJU56dUA8
R5NM7Sv6mheNFTGQNf5W4VRzyaebQl799uMDtqzPGPHpGZqB+0btPOXvGTzk2W9nERTuNcvEOI1v
oSMISuQbwgZfb2bH1B04FRKXjKS/Xbe/qdjp/Eai8OeLtDgzi0Ru7KtG4ZaYxYn6eXpeYXLO0wNr
cghNyonbZL1OUNwknSqOXiLi7xwcfy0ZaovfEnZucMqDoFZlBbiBcZBdV9uLGngfs/pRdFiA6NES
n25psYSBxYyMA1SNdNZYvivE29dRaMwWysXmWyEkfqWnT+2LmBzHiGFYHYv4yU3ggVGmH4fIjVx8
7Fw6RovQJOYkUvex5P3ejKnPYfIGamaUStmy8uAPMC6JTRK+lPH+O8xEQvO2XI9bTtAZObA5V6A9
yU2VUskTpKGj5tDPdcAWL2sDXYlHS2mWuJQGNdftr93Ld7xH3NB3AOoF91KddFxR+vOI8Q3h/KRa
ee1GFawgX4lRw+inqruQ7iV8dyi4yGAqwuI9w1leBXTRK2D3eKGAZ6/UPminJJdPw16+LMQQjAdh
22nV/fbQEGGXDJ7WHjOVV/OFo/F+HgYy9t6b1ZzoFVGAcOn5Sr7BA87cdzFGKCJ3JaC5o6Nw/KxQ
2bBe78hVl3yCR87yiLrMpElJYaIz/JTcxKgBnKxzJmXuYOuaF+6i5aEs4dM/YiV9cfL4EoErA8Sb
VxFOTQ9oAkYxIOwkgie2WbBbbw0daQpyaQ2FYgwPLcfLG7vNHMz9c+XPF6BwOo7fjtHy9N6bkEmB
rybqDY65gy8/HLLbq/exWdDZhqRxtYLYZdQg/N7+TLZMBR79tN4xK6fxY2fus03jnuv3MC2FceGJ
a5IyLfI9cgtBNKLuvsjTU1vvsj8WKFQRXqZ7urrgK3F/b/dorJkYPGPl3vSiNUhZzYBHAMBh2V2k
WaUC7AJuYyppc6Iyu8Gf7zodg4S+VKpgi3np3Tv6T7wnhPVSlMuWbqKz7+ORc2FSAVEn6xX//vDV
Ex7QrRRxDY+aKV7TslOC3aVhZpq5ETsZdI2Mt8WnosoWLbBGE0DOeVeoc33VocbwSa0eZkUndotR
DD2o8YCZLolEwB+lNp8vxWZkeUWtKu7Hl2kl1V3WYm7yV/dERYOfZaX5chPlaG24xigtywExCDR/
W5awNeVK14cxkMTiJpVMYWtJSJK6pd/SQyQc3apOvTRxFiNZ6zmrVxSUVowEeRHHWxn1+QH5MNMg
g/0os0uwNM0NiKTbf85RVt9UqDTTUZKV+6zAD4H8aSL83ldA/5KiR2w0YBTE5ROdM7PYBoBlImhi
TtMTeBrsoBPYHE7OxHpoyGK9Xhm8g1/nzcHaEDHQCoAglZ/kx0tBw96EmZFTFQszc27SokC4T5Uy
4qqXL8mtx9ZcrOhNtjeIqxTZT2D9ftChEUuyVuFRfCFHveORYma40KW2PmqvZIYfgqpP4WbQYNch
r1mTARYR03jelF5DkvYjmVu1HJOMDwiG3I5OIm2L8KzdiDLcwbbZYZXXYdS60ZUeKJNyo+P5fsCN
QTxj7/eVHXS0HREhhVa0KJjIUwsH7o00KOa40To6IUBIyC+3UxCHSry7gP7o0QO/oRoSNhGD6YWa
CijrpvyG9Fo8r9rTjk4Q1Mhh8c4TZIg2RBL4nCMnuPLDhZk3pnmusS8fgkFL/cWiLYBEbGseZry/
2mVL9MNPT6uiPDUuF8T7LcPZ6Ct+Ib9uuhYmX9joCISjAjhIY/irGYArgWfFVeQ6/2s0Kl4sze9U
X1N7F1juKbXJSxjIv/fLTcg/W6JFE1R6uLybU0vEoNweJENDWid86v/kSv3Z65O0G9KzylN3Li+p
IXe+6gVrwFWmWvE15qIL3Izq7uOCAGFO2DRFf5/D5Y1N1VVMkN5YCEuIbPS5lEQQw+LbBe7FA0RZ
GqwmtmK+8zg5iSYJlX6Q8nNljV0yWV5hVA5Of9GK+/Bqxt0thOL+OLASlxUHYIe3euZvhigo8QpC
U3Z1ILhN3Dd7oN6yUXoCj7U3+KKILNCOoctiIJ2MfK7+78+mQ+5E0PLDXSv7zpAS6CjDz3OSklRp
+/yIcIvK4AhEoZV9QTzSruE15jbT57FfVGP/6AEMWyRDX2pUdYzo4hWWROqMhB7DRjvFLvILLkCp
YofiRIoa/SlbyTX748fA0Pf8ykgVj2fIc7OMKg8lC5UCZ6OdsPUOeZERPcA2fB7XTR0UUAJw3mCV
Ou1m6FOK2Ztuh+toQGMcZBy/1KllbjMtxdc8BmrH/4kk4LEagsyqw8DjhnD1Zj/1RuMPGjfmINsY
fAP/+LKrqD5gXpftK2QGq8zf8XO2V2VPVBHlIu9BioikBVMHyuLOsCASRxTrjpIvXKTj/im6rGnZ
8+CiZD3FNIW4yrrzokpbHGWqnPr75iBtCxSxdwc8vqDQ5/e0DbS0EhlJVtMyK9CslYC8fiPbu/q9
74yV9VAdSq/HSGix0Ld7oL1jmY576Pifgbsk8fzTbZc3DszVzS0PITFFWFhgN0irIa2H54SogX3i
Va19DaqOG+B3J2ZjsUekLoeO9jx0uo8/qKl8SbZI0GuTXwZiUMHiiw4FNHVdBmneYpHi9ZZczlCD
JPT6nYx2wWYBF1jGe6CSENJWCuUegkcXIsbf0Av2/RqiMa/yv3/bYZBEe8mdquZvbGyRngIf8Uqt
CxrD/KypfGY+FXYqJLawNMP5zZq3+HfOV0BR2s3BpOSEb7FpMBNeO2xJdd6+evTas6YEjVnuBTpQ
dRHG7VdGYQQT3B3L+oknCn86oJikdEoyDy6c2Agay5EGdG6jEe40w+LuWtmeTBnZAvbtSIWgOuel
rOZWf4BPGePEU4uPbj5wKljN0H+HBwmJd9DJ3wLbgjSAb6izm1uarBNN78kdlPLR9rTsBJPfXmV0
Quvy15bXdDvaHGHs98YgbHnCTDIBP4yLKMraHwXD+pGKprOfkym035LOXMLD5b+9wL9HvdaqYf8E
8JoxVk1LMxlKfjzzeCNqbZQd9cvIxKv29jLjGaDQ92kW20t54zHljTXU5tbxUqDbwRtf0tZbaCb4
uQxdoUQrBleBr0vh5bV2kV2jsRBTtcyjwVpLv6FkQP79dU5aQSEblvIsddhxidCnLqFLoQtzogQK
Ip9HrUN874oVJsN2EqHbOffWGoVJMGIhnwqJPRmSenyzRDL7FdJ3aH+WoJUDwOG8Gpp4FwLObMWn
4eOea/naSuAnA7PoRCmk+y/1vWM2gTd4xRbJ9yZkEsd4N97I+WOWoVsMlRcsZcJxCCiYlg5qnZVz
TcdBQYe8+/MBxcK7jR9cyIW0XS7pvke5YLjvXdk43pMiW5rnlQFjLn8d6XqDHhxEVpzSYfvH+e4n
8Z9P2MSt2lBW9vhb8L7gnbSLz1i+chRQyvgx7kxExl4g2KsEsGe58/VKu+18wUzFBCMcI6wpCplS
WUukPD2W3nwnPXCgCmqIRipA/VgiANDpUWcTPOpJMe1Q+obwc6osnt6vohCg1gvSCmHazbeGPb3u
XyDIb1XFOPMlv90yJWnruGDkYsMpK8D0Ezb+8jyKCcMDWXDqbIgMZVyZQNrh5UiYtBqaFXs14idQ
I8PCB5UKOSX+aYZTc4IdJByV1nJ87nlAXihywFHOazOSEDFWv6kkPutLT9/wLCGbLOPKRkekckVB
hk8yNg0KeYIYzzHQ13cf+mLNer0iBvF9BmxG3aWkdllLKVx2EoowoatWwYAmuhwBsjJo4qPciXCt
mcjfIH9yQZuEPKmtlvHHVr/UlOLH/o3m09mO+1y2sXh21QPMGIlvTkWHyeAUXMX7xDBijqAp8amV
+0XBgOogkdzZ8YR5w3DUyqcXkwiEFue+7gaZxCHEpdOy2DeBYmUOB8BBk9ACAotPgmaqTYFozsSG
wx0wbaB4J1PbgvgZzP1eElHiIiKUt6P2aIz2LhhvOMcXAc0mjGVx+Vv0JBIyyENjYmckzwreBLFy
QHR6KaDMMW3m2szTyyr5RhYaDNnq3J4T8njLa7zYLKPKNXeWOgA8IQF+Up8/g6Wsu+PxbtQHUlL0
ugV4Vjl21oSSxTP5/o6sxFgHEit/WOSDTKtJ2jQ7khOSemmfn7n3BoTKP77p8WODL8+4tJ+jsf7i
sZ+OI/4IuwZQ4YFHghIzCyQoJC55IoFGJ5Za2b8S6tn+umxu8k08oUAHdPxiGBNIoWMbV9GUCnav
c8YxEwWjm1ht0qcoz6iIZP4E/Qxnblbq9zdVvihJmEEtbbtBdeBPDnVzzhRKu5Wu8sJU8XSAIZzh
UAUjH1eoxx2llVBBdcJq6DrwYTuqu57V7dsLlxUF6rCT6TPt2o6RSlktilKG84ZGBeuMoo5OJj/a
vKSwTjVYAXxFyyZbfLVEJoaJWrOSbIK2+Wh0jZm+Up3iHdy7wCipt2rV2mNdPzKW8oQGnRpboz+Z
0Do7hzKz5nc/8QmVc3xnzvGzbsdImWuIUlSnsTcrAP6qtGgGMJah274fTmezU/3O8H//GrfqA3/Y
kSoIlmixms5ipkXR3D3ZtFVqEQno2rSFNC1BgHYpEgWAM6zzxCnUsMoXTsTX7MW3lAZxXq2gWy9S
A7q8TOkcS4oqjQuCPO9HvfT3vVJP02ya0OuSqiwAbJoVnch6RZctYZ7jfu9AAKxV4VxRPsgLKD68
p9PvtJvfahVPfkpDOPkFJ6oY/jyRTIQ/SrMxZoaiDxR77kZDwwZ6ZANA54WrhfhqS12EhXyEUJxT
BYsOy1idgR4B2Ec4RloOQz5ybCRO+BNdeDD4VmdSqCa+HMYfcRvllC8+QVP5/fvPK608R5tWLTGY
+oFJmQU0IHMGZIy739GnE66c69C0ACRptIoIoKIjvHfVY2hR5f4hE14vYXmonnRgsifp6LFGjlME
cbh7Asl12GXda/MfSeIvwNfYwbKalZpd1DNhURtgkqobBZAcRGb2wHdtousdsLO75WpRLZH1ApG0
iSQuF9vHHJ3a2T0MRdymzIJ6R9YYDGbs51YOnVkAOTM8BzOP4XLm+xEHjvNsw9M+ZIOE2fDbx4Nk
7uRxA0V8nxLeDBKvfhyU4HBrlZ8INiIt0NaeGrgyELRMZApqtBK4swdZ7yXzYrlBVpbHF3ibwpoC
iecQiquQFrgLJFX5keYN6R7MF9ZEyGt3SEVH7zj43ZTksMZgz0nPqq3R8rmTgyFpZOEMMwZEyXNp
cct30pCFz1KjYwxfNClLHMjR87WotT+t4bDNQSG4Gm8r2l4LADbb0V4WSiKaUOyAT8nnJ6pYBOT1
Uz9FCOyZ+nq/4rX392rKdZW1s222XJG1YspKY5GigucQ2jMd8wTKmrbYIM8aUeJ49s+00otgEsdr
cRWllQPeyEn9EL5xRepSRIw+9cNIB9/FrN+fhpj+DKoXBGO3kmyWPyiNVkUB3F2wkNncX4rtDPXA
N6313pYmzz8Dnw8prqCCC1UBpCiBrlbAIOTtJwko8fSOQ7Ewt4BiLpCfIkkyg0bTh7hTDtmkol8X
dZuvljsAMuhNr2p/8ptcvpf2pO5bScxt+jvwHaKFmqC3aE9Rb9hCXJGhnEJBc6DBwlMY38fLqstf
NMWPxoOPQ9G2V9I/AL+Qs+1bSDg+85NbZdyrcEfmLOwWXWMBID1Nn2FwWtEy/HYF5GpfHOuBrNdd
+P4bmEiyGaO3iJGLyJSxW8UCt+tO1lS7PoYzRGKkmS78lA9BVzod1ir5urFayM9CHxDwmn1S/VsO
yIIWmbpiht46W9n+JtIQ/buRu/Ms9X+PpUEHWFxqTZzrB5JRnz9ZQhb6IF3nkpMmzNwPjtp3P3yx
c2SdKlq1wplf8PJ4gmoJlE6nEbVKR2/RaCMf2MyuNTdTcwKPbTrxXxBLBnT7Zywod+D2H8B+pD4o
paNBq9anDoy20+N6mHthwLxfwGATrJHFGWPXXkjU8s4ySJBUTJ5VEY7NmB8uxGDbylEk0dx0irb6
T/9kGzmAKvgBKVKwNYpGknY4yUu44TslKUub51h/0w02um+PULfTNduuWWg4tNTZc1QE44BGZ5zU
QR5ItgPUXRZDkQLS4/teCPGQv7W+qE6gRdJ+VWCtLmd3VuyDtfwODpW6GQG2tJtO9GdUFhOtLHrv
BFOXYHaBLxPS5ElZTuicXC8gN1PjwQGCki+mIqqU7ZbVqtVUNJNoCzB/arEKK3DLq3dNUXZ33T45
mxRsggnz4ohStubS6+lgyAu6WgHtF92miPVWhJyG2pI7QevfZMcdkjVT/NmelomQJD3zMd4ppYpb
RGsjDWLL1pDzDFaR4Exsvv8sWJrLNSOzaUq5iB5x2zz5TP72/bwPCVtzsu946TKViRYMjpwGrtK/
vJ6PnM6Nn5sXxbkmOHkLf8mNk//QNvQ5TzZWZd9fhVvAs5iibA2w14UGgR4m3zOCSIcuWZ5QTDlT
B6e9wNSJ/+hQpeeEaBBtNNJs8H29pYBMv4mGn7apqNt0GNxKTIBxR55SY6yKN6XpySKdRhjCdcGd
HJd3N/FneYhRbwmBQaYEAqcySTGVKSyvF4Ns4ytbPGUa2ekj9YqwfGmoeA10RYyNWOMMyRbdoWfn
YAb9IwTMK3D9vV/nDEj+dFNHjGb4YHf2RMQGMRjPE3oSeEcAX87jVRCoeaAW47rAGrs6h3RuOfyz
lBI7R/yjJOVeZeq1qWzreQuRMeUc3tBxoWJcM6BGY6baEPi0e/JPZ7UgR8hFIovzaEPE/B8VFeN4
Cr9YNcV1JLKw388lf3At0J2o24m6X5qf2LDXqwj1EKVMTTPV6Au9SOynhf15IApuV129yUVCrfif
fOAR88k1DuhGvZS1YePqMuJchlu2/wK6nZ/MUTvCCqADJGcPPUz5yB4tBZuRWzWEddLWL6VhIQrK
1UPnKHrDPtbDH0FeGRESW9NeXheEK8LwlxQeY9LJvYs1qmzE0JCDR6VueYOCYmc74hE4HJjSsW0h
9nOIT+PirGFYWJZzKj7HIL6vZb0lcy/AiRnampsVcX1lgKo/CGeYhj7dVGhf/XL3ZD6QbTxN0a51
EqcIf/21irjj8uO/v10eEfI7rPRg8cMccF23UzFxbaMTtDwPFvA300mFa7rPYWgMH22gKkn8Hv2F
XS9uvS3MYrvOYe58sq5EdhuYD64tl1uVabtfxLEC3nBAAdKlzBQt51KjmteeCAdqEwhDj7ty3ira
+pFCn1xxcrWsR0BWfD7JaCPTe0EyxqAUiRuYh5+yy55lrHmAlnlWiof3pfqefMspyRtkp1dl/HKY
lPsFytfPPu/WPFpfaGIJiUUB/scFf3oxqol/rMRHGNBkJdYj460+N3dM7NFM7x6t+THAs7VZ3Os4
owyXbSJDJhqnTCeCCWgFJhC6xq4YW8Jl6Mz3awo/ysqiyeQTMqzLahAEta24n2TjO8zofbg2zTTW
V/tn5AwGRI3xWQvY8CN0vLeQ3lOadU5IWMFJCVFo3OjHrh+H0Vl+8AYWBNNZssy2oS+93HEhVhmp
kRQxghAS87+epDhhIZ+QqycfXJ5L1HZbkSxU7FS+2DdlRe6I4ogzeN2XQpJoj05n+aYgg7Lyb3dp
iRX/hhIfLLdV0LNx4GVPqCtYqe1srqbeSoY7BbHHqRV8rgrP0VSpydzQ3rFQyQb0Mf/jQ6tMQZGM
PMVQkpEje0Cz/B3zPdvE/qEJkoj69ZVMLjnls7wwyrB7ZnGAajzL7Eajq5rBR60qJWWsWvL5lVZY
P+X9ilEdZdZ8CfXihwmwxht1waxo30qCFfSkAiyn96+WVRh/3tekIqaQAVW89V1rBE/Ptu3PoifY
sOjChaonm0kIo3U0EKM/ij/X49biN5bZTA1aa7NJm0QkFYHrNKU48tO49BMAlyWAUkVLLOvDntf7
R5NLZHWpk9XAltPIJnyIpvT2LwcWSAYwUcoLjkf9mnd5j/rih/OBw1KJctBtVW3cSRoLIXt3k37Y
8qYconluqdnzVlPasqRS7YyFQwyFUCgeMRm/VXThhlTa1UBzf9LiH2YU8aBwvAgADzbbRUDWd5RJ
VivAJjG6kUMlY1aENc5MZmjWodGbvj8k1SgHujMWnQzmUsJ18LTg78pN31KkDDD7+CEX5JT2PXmC
UCWU9KGDjzgp3mWBi5AeeLpd3I2930QI1shJoz5qJnKLb6Rb38QQRzWtWT1VL5GJM9VKYTmGmWXg
fO9Q+VIiuUtM3n7fHjmWkIZHk3aD8TqjvYmNWiOrMTs1Z86NsGFAd8kJ3vF1zroAheNE4EIjALiL
rpYrjeJTTL8rw5KTCNX73z9SbftWm00B30xnCuqT3A2Ri4n1xC9RfhovQQUvKxsJyku4xxjJFUP6
5XfZKNT9awAPMTyu0UCUg127j1JPvEH4hPtEn5J1dkqG8UrXM7ybCTF1AZQ0+vei1pjZ0FtwF3gW
khzD2dn6kDg48YpQ8D5W8h29kWAUlm9r0uV1Ic0u5lVvjLBAlscJOdGxL2PrDDXLww1t/zlydCH+
PwPL4gCJt/KjkepL9NQ40EyGCKoYbwmUbP+p4VJsawoTdLI5iGkZIRrRXMTi0aBHuDkgIYxHsgn5
u/EwjbZs+JnvoXJs1jj6YXLvoTlT1EPxBuf/jZPJyvS45rB39XFx7GA11K1nPZzZYCrLFrYiAbzc
TCgGvuNk23YxS13/udU4DPfv6gWXmTBBri1AOCNwBpHwbn7JHB8kTsNns9DiNbhw2e1JrMsAG9Fe
Lz1jKKAc7C6AgQDYu71RnvC7cAJ5M95LHAR/OFB0nrFnwOHK41LnBWaWAg/2uWGikTlY3rjz1Asb
pxNrOFt5Ema3ghcQqe4I//zIufcX47WjB5UmllUgjTrPyjxpzfqhOWxfHnBMY8NRu3zYokmuX6ey
6rJZ4AxdVnR2yZM8Bl59x9T6HNjFrXTpV0MpXiVERjL8Gk4S5OfI4wXkoL5NjW3J/3Ot2WFFcuCN
7FMECEXPYfB95CcaipyT1feq+1y6yyv1nP+rHywySbvf/BPQbN0GYIVslr3higEDDrmOLJoN0NrB
sKlozt2CxYEnYGBWgYkN4oMH6+zRFM2D5AzNpe1JJXjbinXvWb8X/LLFhXvJBSfI8aRNrkR70wMM
KnxcpchhAAQp2dtxqhq/9Llm7c/LPcEYewoZwC4pCUklsu1BuNM1Gs50vBhxbEx9kUkFBz4y2R8z
6jloR7OrvNwCqf/UUVImD3udE9LrzFa9zN8KnOohJ2zhvJqHo3OW1RYDYg/X4zQe0gvHWRCBECD6
mPjRf6qMRVyiXitrmjycVvOpIoJ9sl2qRaXRwDjuQ4q7VLI8xBNZyZIUOioaQMXBMzEAEtB1rBf6
uWASTEd9fkWcZ3JmTyLRrrR/1JwNWfikWj+012FcQachFTyejyVzh4kyqYDSx9qqPCqWpwAMG7vR
YNJ0SmEAe2IEK23vbCnMXiSs+BtOp+jMqBYlrgHGPoe32qD7s2FvoDexK5aVXrpBSYV+bvPGqpdU
3UekUtBUt7TeuX3rVDzfc+4SjDFv1k5tw0R9Qw1OyV62QEe9K9q1o19NUhW8SCBaZ+y+Nj3qvM2o
Ok9THOoW/5ycyqGz8GpaITDAIDWUygTzVLQgEwYjmNkfVwD6eCMon3+ZhjyFqy4ZcduCMv65tzjl
Ge0QDyRQ+pzRecWd/6InIJqsvSd1zwUp7U9O3y8i6ShJpD7hpR7VD8pvIvz287aYXr+5c4GFZ3nz
t6D1R4axIBSLkh5UcWsuw7caB2sMjjBfPnWJ2hNRyoIEOwrH80AZrQDqKFNOYkxMOz/8MHTKMggi
Jx0FyxLcJNOaQ/vFKxEttYmYZd3YXIFvDhTrTCPUI+xIDTJeZpcd5x1Bb9kCO1MVKFQHTblEpDPP
uiwfz5/SHF16dZK/PIXQZLnMTWBhDoEkyc25nFWiJ5D7XAfcGdE2raamcUMdok/KtO3pxjzcj7ZQ
kAwlBv6S4sQwxFsaFhbN5eHMrKQYil0EfG/zhOOLDG9XaEoe86NqclXmQdxR07KD7h5rjfq0NceE
NPu2ATLUGpfKicKJAc+naIRF2+NJZiqJ32OpbeGdrZAficIQQ+YqErEL2HVmBsXT8TiH7bFSmGOm
0uagSCCO7mzodPDbd66qPix22ISPlTivpnu4ISL0O7xSsdPn4mPNMMLaPTk3YBadk6++SBtsEapW
Dp1+dGWUTA0CX1UQAWcwOJlyFhGiS/35KcmOgtJMXS7tet90WNPdP/tuawzI79BRzvO+yevCvi4n
SpqG0y6CiPwD6X61DriovMFMZ9QAtjFLfgTiPD6hAMvDdWbzCYaGuo1WI7FG1Pw1rqx/8Ano8igY
loeDlh7YdBtjniOJRlMPNcXyOfTDb/vJi4EB5VlhM2jdD8MLHI367Coz8ppFK7fg3eIxUgkGF/OF
xehZ5JhbhNBCFtibtp1Om4rP2B7N+mng9tqhswjVMRq42J6WP+tKI3/SI9MGmAjNw5l3vowb7Yp7
EHXGX6m2OPpw/XBxIf2iVoE1KW4K2ZCsN4Fz0B8/sTC5ta8wFG2TCu0GmoCkb5k5ygcuI0VBWzar
IiT/z5pzXaNzXqMx+B5GuRz1h22orPxhW86LI+vm+Eudx8xQJtD4U13As60FV2vZPnQq2Q6aF9fV
LE1z/pq2B+8cCFGvPRUlefb4LsQsvZa6I5HOYOeswLDUgGq7SsZC0u5Dtq683Mhi+EwdPEMpXR1C
Aly6Ql0X4YmH8XdkbshNhv+J3/FAMB0KoaHi0TsjKbe9fX2p3yJT3dIH49era+jiOHtEYF+J+DWZ
s9Hahc+4IdwF9rKwzvzQ6ZxORUu38Zl5Xbov1TN/kzmVga1zICv+if2/EjKAx3rhte725QVF++Dh
RAJcH0N8hjw9pXuyjzck10+V4G4P/OBj2RgKWpQSI99XPTMCVgF2Y3Xh4i8qsJV9LLPFzIRUVLao
30VETiFNuQl9ttftLxTQ6iaQOOdy66c2nSAP41g8JspE1+l3kpNMg8sm6uYKzfheJikkaTjbCU79
wf0L2eKiMF5bMpcz5llYTNtglCspYFr8CHBKJT/idO/vutWPulRV2nRQ5t4DItv9hv3ViW9Mn9Kv
Tq8mZex0p5zZuO5vxavyfxLRzL2YLpPmHmmakxufNjVMgOSpGgks4RYOEPig+e5zu6rJVHlQkUht
l9GE3J0c3OX8Npxmi+gqek3/aqGKAa3gbRePdCs5awpMLN/2Ta5T5yLZTVXkFW3W90rPYP5pibwq
z2ERaGRNuC+7pqTBvNuP3HUJLFVnJdeGbwRuZRP6w4NbstG3n0QC9wZ9iLlYQ74LcD2n5pMju7Ea
hEAsM16DDenb59BigQQ8Vu7hPiQzE1QTQXjqRRtzqpQZYZpxV/sNUzgXwAiGzhD9F16Tm732HEIt
zVe5bHgVs8q8vFfjNPaaH/jWDaO6Dogm6fKwXLF1KhLESrxv79GutalJVCkl40EWFlrxgIHAuCCF
7t01EIww1lyOPmVKqDjYJT2uAPgY/g9/yBB7AMljkHWUmAo11fqi8Z82zRqTTOGXPknUGc0SbAHB
vS9vLElHp6/QY0cUkjGS9IhpKVwFDF40h6ooKykawSgkYht3wC7mcOTy5YCpfMZHjIBYFQgQJYxc
P4iu0RKmvx23hKeGrM+iYbZTXGhvKNeS3Cxeaw0UwMcBL3wZszOWsdKoFMzOZ27cAE1WbLY4IPtU
nb6YI6zoD8+whui30j9sz/xdLqCn0p7YA7ZhqMcdZgbkatluIr/f3PZ85LyMcnP4Y0dSC9Gzjky7
IGhLoWUP6VGr+b/PU6mb3UR/OWg+9zwxXTZXjl4YCZenbDEiWMXk7C/ZLS2U7nUKx3Qvi9EA+FQ0
R/hJERMk3oGdVdCebfRh7OebBMS8ns5Vwm4FbN6CQRt6SMescLaEOfEIXyVnV0/70LCASbUnj4Ij
1Ujl3CqGxY4J7nnP3R2nOQ4c7GZNcKzsdD47xJVs99lgNdcHdy8cKR6F2u0m+6m491Uyp0FXWDBx
D/sK9lLqxTdTzb2k6RH2NiIANuyjPWdipRdnPbki6UYlf/TgIXkhRPJRcyisj8xXnVkua1SW2vd/
RgZXbB9t7FHvSkUPvsqObfr+UjZa3oTXtDfVa4X/LMi+G7ZCPHOZRBpZl/LYXFxSoQVKaQD/p9kt
SPst+dGwc5MFKqCvO5yR8TbJ5sriFrPmKFZNlSY/5TSek87EJJteJPkYIT+/VyLoKOdY7DUAacvJ
4cVIuullvMP/D3NNiGgb5BEKgzLe9xcGjQMSgf1dufG8wuc+PHqRMBeNW8d2CMsc3Nts7qW4zXOb
5ecAqEPt5wGIITJ3fLeZHi2c5x6lxwmmgQzYszIveEUGL4BtB/L3CT2SQW/JNy0twNVodJtP9+Nx
xotrxD+FRbPU6Gp98HSgAaLE0C2m5fytfUbPiXOP+QSXxE7RjZlWxxyC51bcxvg6BKmSdFxZ+K8x
A6WABnkIq0rCmgwdlFUx7rAl1KeJ9lGjXBq3Rd+iq+Z7Cf2dlMYv9wXqigktLlUuud2d2nO8bPpH
JjFIf835M//boSHY6DgdiBBiA8mLvI7Rw/yMQjVmU/Volvy/1e2G6Um4It+5NHK5KZ/tc1A5enUc
Zm3rGYXvsqkOHlv+TP/GtF6Afdz1G9mr9gaoQfiyzgN6HlZ9SXGNyr9V7+QlxFvrnBT8wCVvr1wy
ace5XPFEoljPq8WoazfCNoxAGQuNK1f3pzYImWn82pWvV+H+J0FFNJc+ZEVjCKX61En12IGPTjpG
QnJeeGlGpheCabQDw+ICbHWqX1gDpA11vfvzHBlQAQdgg8I4Cw4SssUh8k6Ned7wOO3lAJB0afxX
tDGbUQ7f06nwm2nxXxK0QyBzEeQThkHUj2oB1nP4nP9FHdAFUgD13Ak316Ob6F6Mrp+Wype2Kcpr
RKXsNITvL3szFYCamV/xTtZN8yk18L7wXszGR4UBNHCr7cqXQgAzkl6qENu1Ie2gYrZZ5XyO3dx7
LriUHB6FFXOk4wWTwewKOJE9aalOt7s09AjdYNh804GvQ28wCt3dht+pjXhZZBYjWFIy+Zgiuor1
/NRrh/5piEQoo6e7izixGQdodQAwZb9MC2v11MmhTq+96HzMuss+Y1tPFfxTiKU811hCcB+bXMdl
MqKzTyYDSEnRYSEfCFKZUjkHbhTfWh7nhBubbkNEVZr6jTHyYmnhu89tzZpyompXwhXf3GBGHvwA
NhWFQYlqROqQ9qMX8ufgYDFf3vsf0pTytamg1kjSKX7NjUIAm9H7kL84/G3IJfinhLs5mzE2SV4o
Zh4RCifqdoOBSmUm0RTf7zfn9PlRYdxkTCdi8Zky7xq1cbA9y95jHjwujIzWY6aAsmLTqZG3zePb
mNUTkio6DScPTxGNrCFStGkZkrn5VhOgTx31EccbVrlKbtvu1q7Y/NKCd6+6GpxEeHMK97wicJ5s
7oOxBGVWZUo9px25RDkpIV8XWMYLSSpV95BU6b7FGOfVTwBFHK6n++3KW7RaiH1O+vcxCa35pL0x
sPNCHT5nartZ9rEts5lSX3hbJeMiNd2tbKEiMfWLMbb75KJyDbceKmperwPo57Gizz666KvvVauq
19KQg0mY5eoes5ayXb7IA/8pDARw+NPIKFxSt4rZeXmw5X7vu2Rcvdn0q0apI4qIxIPhB1gmA6BG
b27devo3Fr6Ze+SwszEE05SQHEiYRUIQJ+WRDMCsIXEh32DswJ5m5GYSszeBinD3f3p82RBbrlKn
D+mUOmZTvIdxcnC/1W18u5Nml13m3EcHCtYMD9u6/kovL+nqWe9xhUCVle1URj+hpbuAVuFMsbjP
p3Lshj67KNX7q0j6LrfRlt5enhWHM7b+SXFyf+O+StJjqDN5zUc1eqgMNtCzeBjPO1uMU7ERHrr0
VzmiikzI0pyIIWmSf8DjVuRq4DM6Q0T+3zi4hRIB+Uks3scROLsG2VE509EOzQM1pVru5+k2LEP0
Zxb9UGIoDtzofN22FVScIl9zxopAzffwEQgsxz20ZXXf/ZX0EHGb412zDYqvEqSnduSoIv5RXQaY
xIbwWeEyK3XYE7JQUpiI56ox6QUfVI2Ao9IBytzJ2aomqUFNteJVb6IND8xTLWndsL0C8y+UYCgA
CmjT7slR1+fcXWlzN4f8NJ5qcokytH2M9jLPoHBAx3PKPjMW2uJR/AdWF2LyYj0PRTzujj0IsfMQ
BQlgxDq543rqjK42A3EwcVh0zC1fPPYNMyeyTWgCylwBJT0R6asix/TbjZGSQ9Hndn+6aaOYxueK
XbPuQ5RoeqJfJapTH/TVvEyAaIbvnEa9Qoru3nj2MxW1ZHA6b8kpEL7SxcYn3Gf9eGd7Sg1I0/oV
t+uZyWuwqTYFRsWW068ZuzyUgjni6/e93Vnd61ZGqYNUV90aOD/eOP93XE6fgWAA0emDfU+OPknu
tWtjnWg522wNaP2RTAZy7bVGPFJ1Q+KPgT9cHTFr70KG/C3y/YUHUv+fbf4vvtzxNopJNIsDq9of
dBxv41Dc02AboDu/fob8wrum4rRDVLlEO99lKRYm3GEQwni8bTCaR/SpFZBgBGOiY6WYltzlU7JA
UIn4AkwoLxLByVk7xF/bktiGQhobpKyOWe+fadOmCCBWZbjIyjxSxpMw6pK+0JHSgVrCH677HGQ1
2uaRfX3KwNYyo6WF2E7oReA38LWIHgssLFMzLUxl2Pz9OMmKulmPDQwZTvMuz/tHhGdB06AtoMnT
VYb7E5rl4P7pdgCXCPowTiULYqI489jXiFa12F5DEGvQ7XH6XVTlpzbOmCHBArFXahQDj6knNNpD
xrCca+NErmKOdREyNmz6mLgxwuUH20JtNZFx1/AZSrBQyQMxvKhSxKF39xn7Y9T8T9oDJ3dTVb+B
znDzyxSFLqeUQZMfZSeev1t2OqX8mpRTejaxdxDxCcpJyj+OMlEO6AcyNxJHXhLRst2BZlhSph3q
FI8OHScuOR2eucmfoZVAd67HZ0Ue3fWeLNxuk79eVcGi/qldiDszXYMHQBbY9PWv1bXY+gn+zR6f
4jhmclrqB7CkwAxH0T8i2aLecMI7lmdB3PRHu+DjJAts6gIgx24NkUCRzYjVobwRw35nWps8Bo66
LHp7laQDI/bn7uf07xqb/nAsKWOMdd0IVpkwd/i8Biqyoj6dJgYXYba/YoE3F33TJYpyCIgtFBLM
yecHDC0glPsvQggoBEMl8dEiaqJjyKMvI0u9xAchXVwdxgfLhUuidFgVqukMJctnMdtWU3Xei9vI
AMBg3RpvzLtm3iOZEHJyS32/1ycAwcTkebMxdo/y6PtXJM7qnl4olOUWpCNLtkws4k6Ko4PYe7Zy
EqKxAterjzrpBHHSwJ208gOR6e6IrB670V+Jl6yubVrEA7SFdxiMjJlHs3LOX8JmmApZrAHfJHj0
HgkvOvcIudGaJoSGz6rocmMEIWDDxqKkzOKJA4sZS+U4yHCvtPK2iKbB2ri4fimwE6mpWRB2Vo6y
OqTNhV41HBT7Oc+noKQYfou/ZrILddoZHLYF27JdzV/10Ae77Z+J8Hdd/z7rQKi8VuEPZH3PoGJC
Xq2iSdJnfMwH0sesQ11WeMsepY9PyR3NHoGgHbvmjD8PnwOA1qpe58GcIdrIpopHm5oSqRQD/fSP
EVOl5w9CBG1uBZWNe/YQRsaqp4S2l+bVxwkuLkhJUP7yB9BawnfeHBXiWbxjogHnPQ0PBeE6rMGV
TEGo0qKBtUQ+3NjzvSfLUxT6JXrj+UijaafoFb2IIIACC9VDSda3p6JIhU0YFsADGBz9YtRRo21g
DG092vkVgT1uT9eF0GzmBvk4Xi19+tlXaDwaKvKm7Jdt2uXNo+pms6KqjwveHcriyY6yQM6W6syC
GdpB03yU+MPJKHml/4fuWeNI0HozRqsBihg9DripPpMf6xNZuNrAfWwAGoQTjQ++ZsSn70wwiWKw
HtoY3CQ7wv7mDaXtrAPHGyxGF2cJMLxvDbWwaTeyqSVELPHTOHy1sCrmkuvpdwshSVd1VrErlJSv
rm/pnTWds/zKwEhsxn4/6cp93PLkLEnHjPEkXnzkBMDT9UwUKthymeQnutTaLy7gcZKyspou1HBm
RP4KFDr50vXldGEvUhtFawZx4ijjOOI7neVqV3o2TE/vC9ePXlJWlVTUZeNuLcBcJ7gYoW0zHQBh
rzXxrh8ayULwsUnX2lDJ2O1HcGXZdffV3WxL2EqJgMiJYVNyNzjZZ/BnhJADGfwJ0xSYbyDl3qFO
gH6QtlCkQFJiJGPK+ypeDzUkscyv8LasU0UXdBdp3HExiIz6scypjGla2SkEx2VYchFsweTXt0ca
vzDOuwB54JrRbJi7w7x/3bIY8yeDd15C+Lp8VMYj8yaP4yEexkxTDRMkXXw4EMidFadwqdeq9Jaq
aURz/pt105jA/zRsxiBVYEromK+IxiSSmLRiVgXIb0OybWW43WwmEIk+K6Cng/CaCJhY8Y30vBBS
BNEVUd4RqshYBUwz6xyeODNtQGbww1UbSkA9m7b0Mj+cEEquut/fH4oibyU3lgvlgS8/WafklE5g
K8PIlWI0shj8Akeq9U+ud9G1yPI3IW/F+6qPrkso8EgnvF1Pt1zWK20Br2R+5eVsNucBccNpDtgO
usfgC0CfJ9q2REkHoNIWvCxFxjv5FgaS1TWV1pzuNTQ0e0nUh5vEc9F155tN3TJfmTtDva8gCyd/
F1EQcyQM6V7a1YTpzXAD/G0dpVD/Js7ImsU62A5DSViGMxi17B87oENZVvZldc4kgzoDRKgbrUPD
NWIhwKShFSzbt2ilFu0pgLW2pER6id8Vdyg+xuZfl5fsPBlMQNSGmrc9jnknRzE3j9nJwWtX/jxM
xlnhyu1250zkb3K4TMWAfz9sNLMb7afxed/o3zRVchU7jRh0sSoAEtYedKZrDJJih7EXiRDUO4ZP
REehUFzc56DwJAkzQo/r3JOEOVtvm2tUh+RXTIf5TSZP8ExVnkbWuf2m30ku9Oy9ap/EOr3LuPCe
NxCCpY0D9ESZIbxFPR6rPeVJml3S7LHuZ5bwdoukmbX2v+AgC9NzYxrSk4fwn5omfjoCHFsXd5cg
/v1BjBLnnEJfOc0sE9ojhcD2o9Bxr7E8sbbUUlNrfzcAUyufEilX372GufPmhR7Rsfpj3PZT9iHK
M3uRVufVBkq5u3l2fjFJmm/YaFrMerfgd9MOT8vcjEuc3C7Tw7XIqLSyVgpYWVTv8Oj2HgUYd1GW
sryBKmK4L1/PPvvy5whJIcvOhqzZRwYX3T3jPWWqzpnFVB1K+VKWUDMpdy7CP3QxemKjKac6qlvH
epBosdUzw+XKTqFVoaEJVmsoKj17dn6t07Dy22EFxuF5czWE6bedi4snNvI6n2gjf1RqbIIT7pDL
nHzn4o8fSOKuID0GE1vu+ORNeruCh1Pe3uzgv4n23I7LPGmWr3o1JQmI5C6DfK69t/iPNOXimRGj
WxDPvjNaS9mECf9C55bTNkpPOcC2I/NwbQkizLjq+l+sjRXN5kw4l4+PPXtssX5bc5+XtLIMqSpI
56eik+e9LfQ2oDSFvLIuzPSUKVH/ao18eA6lQE9+cyHGcd9sZIAzsOUQXJHdtbEPHYR5Hgbp4wBS
Hy89oF1WP+Z5YQ/tPwOoa6kyDyuLtZFkZHxsJyM0tGODzK1Pv31TLlAgUAIGVWUBhiiWcXEFw9K2
D22wX1UmCpMx953cXxVNtm2B+yHpPb1ypGmpymXx4bMnm/vLPNx1BEszQcT6pGQDlQ3xmvO55Kmw
Yt09cpIz+I4f6goYe80zg/B36WAGgxucwcBUm4tMTcP4dgh16Z33WeGj+VHJYls78uNujaiCLye4
b+VAv8/EpFFRQfi8CEhl2BPqUs5pu081CcidlvylfOaAaurTY7cbGzXpk/R8IE8iJ0elxP5kqQ77
oguLcFDQkIZ5P1cnhLGIN/GTOB+IyZ2fCtb/7irab4oc6bDtW8bRcc3GR4K/5HGSUcRLjPIcxlix
HERzFhbEq25mY9OXqhZzNHxVcyLuf2ANg1dGoAYpIiYbqZEIZryvRGbkDSm2/+GvM2CJlOKojMqq
wWKXdMLMtmpMmkWLcCJ1HoeOLteMWIUt9hTqsOwY+YrQP/qHysuPkYmi6maTR2m+HaR+6ifqfhNX
2IpFjIlfYdaNH7OqLh6Fx2txHDTT/Ef1y3W/6104oWiCP1yCymqsj6zut3Az94oZrwN6IXon/4KC
8vrnGS1mIgGvmXSP3mzZgp7urYDj+XsUlQ9jJhMD6Qg+7U05epGVPZMtVVh6aYRZFPjeVg3nbOYJ
wtNu5ZdZwlMnLVBFSvjoQj3Yqsk27Zh8/eETw3/K1zCHvAr2RsKx9iyh4Gm3GYVre1JsYEWd1NQD
BkmUM2pgOpHUzMeo553dAesEiGpThb5tY4TD33auHy84TDjRzLex7S/Og+7CS8ZKWXzNNWzZBnBe
tgGBShkV+qiUsAqpvj1G7kh+UeISYBPz4e7YFNGg1k2GgvL95rGv9j85DxwQcOJQ7wwYvOW2hX7Q
JGcqo6GWniKiBIsHijBkHce+ppke0hQFQnqOtsFyOXr/sQIjg/4WFMXnwF7gHB3HD2E14SM2Ti9J
7zyRqZ6uOtrWdg8Ux5TVR1IdsNdKAacLtJbdY5KHt54w5MQe/+mJST0/xiuraeELeeLsiTXeLQjt
53vFaob0gNNFa2BM0jwqxLZd3IKxEbIm9OUw8l/7wrnRtYaW5nH6FxbBgdaP8bTwD5uyLhpveI/M
Sfqc3p+duNaTEbBohbrE/0iSxE45ILNEGfnLEYo67cnaSnUj05sPA/hFwgOlkY7h66rSO1X+1ghQ
AeKBbVokP0KzuNVb5iE4HPgIaJZpz8AdSVk70mtnQH3G3z41OtOM4NjikyiU+O++cwwnZoENS3F0
S+8lqCUgJBrbre08W7zPe98PBVYHeZdvHAIMNKKqlyGie49+BXMoNrGlZ9VSFglxvi9+FaJhqouk
OpApV+pcg2381hiaiabF3/O+Y9WkbLCKlvSTJdx+n3ELNlFGEK6wWn9Bzf8pazWtzXpKwIGzrHsc
ISLxkCM1JvGXKf1qF0+qb5kfAU1FOTjaZbB/bBYHMWLqWe5iaRtrEM4UaaOMVQEsZ7xy701q0Z65
4AOcfMedciwcaxO3aBWDQ8DS2wloONxkbiMP9Dz9zNHVLEaej3RB4CUXXTA1KyAheYUoJvBEAvFf
HBRcQg81ITrOSlqrcJAkn05rPtayCJE/8T3w/EyNlh3QLdCl6wE0j2wNY+6K8kKRfivnUAScfTAo
r3tXBW7Xbj/5mgG+HnlSp0VS6yHWqkZQanSWXaH3hswPiQgDds5Ozm10YEegZoMm2VadV5v9enss
e5jOi58+cJ89D2BYDPkjDtxnBNA4McQk4kn/Y+ERCjJIHBxIzQEkQaymC+xeXxxc6ZSZVuesd0qM
GBkDDrrapyuhGbYqE3lFhM2Z3ff4JDreIbWcP/osuSNzumqWCdlxk2EzDgPohoUVK/tbd706Dw1p
MixOyA5LNp+CBP8YsEd4C+mceS2O/W6pV+FIP7JAPiBGDFLxnopw6WOb4lXTycEZGakormR6kjI9
vh86EYtXb1V480kUQoOE+TODyIlUkDFebuYERfb9ojAhJkTFzuTwRBJlKFX+rOer9iLRaWwJnJ48
23y4Z/KYzzuPWRY90W46hBIlJKQ0iZrjBdOaxuuks14XlzZJxmrMRY/aR0NNXynAXFEFGYyV7/0X
QyskxcIdzKb9cUGiYcMizjWywF2EhU3A59aeuO5sYQQQ+hl64/csfjP0X7uSIKBBc7Hs1TKXcw5H
8p2DgzgZ50kAmRozeArDXyH1u2scGh5jh1zvI6c5ACGhxaH8orVaeEgMkbrPBw0+G1gQf8B/PaMt
0ds0to6iVTD02vdFU/QLiWva/cv/kXz1GvEtCjbYkTnFcowvak+wpfucirLBUlxOl3F3I9B/5ED2
5/EFWgU5aqBJ+BEnfMa8+jhwqpiE89mqsp0rE4bjk31gjXEpB2RriNYO7AOM65jJLQzTzesq1EDw
0dyOumk+WEJM+wXGL0nUz0JdS+dRivOiIs0ig5JYqIzfbyyNXffDtAX4/ON+bAfCVtwROf167joL
watEHGRNhbxhT5XIuCfw7dWdWnDIWP5rYPOxDNN64J60F6OlXM79P9dilcrBbt5CoSyiTJPykAC3
kieWcGLPZi8zdJKIRa61HlknHWeLG2/2CnPbgb0/6SWe3vZvqKuZgonhYqbSxeFIhpceHewftPkA
IgHsBEJHsFLqLcl3todtgib9uOFuPVnfYUh99gxsiI2MBbkEtnHuX42lnJqYN800dLgbnIaze/2a
10rNBN5sw/rkp1ATU3NUGR8Swv8Q8Z5TCpUocN0D56swq5IMP7jEE8oCERaXYDxzzhd5ITvCUjqo
6Hg5dAu8WHZ8l/GMoOEl06/7KEDHb+f3PoacHbDIwNNFDbasqDCLH+bC7TzD0wZRNaP2F46UPzgv
SYLKyaxytDRqO0gGL80saS2EDq0XhoxY558GhImkTWOaNYZ2BN1ljZZT/LaXdk3eToUfvj6LVmJD
Go8tBkY7jOWjNFJeWi3whcJpRPIM5dgdiFQ1eA+IRHIxffaiKO2ndlba8Sla/JoVyqd1jFMtnzi2
tyCLiBf9XNZwcpJytuqRkvPFf7cEQNHQsj5e/e/cc6u2boKnKldCnaGiH7dQ1rG5WkVFiFXKaY1p
363g0iUqbX7kXhPHaVJW1u8UQUfeozae+IuZw11Y7ywSCQBXL38zPn1HOAeItZWwzoIdOgCWkCD+
sQn3aDhxwQWtYR4IDGJG6H4axNUWSLjlUDEy+/g3m6vVRuqQIAvcGD98Zry5B9AueaykVHRXLP1i
H3A8PPsRIZsdQXjPA7lx0ZfMX0ShUljqSIfPfkBQQOisCoLAvo3JiamM02CegDi7bRzphQFAoMen
ju9mEwRq5R8LD2H6Sf3DyUb4Wq/9v35f16HnAv31TbLzEezyQimOQVK/4Pf68kx+vn5WnbiF4gWd
9DqZZNLY/PgUjaD002BWqPbKvHpop659NDojxoGiBLuD4Khj2Wi8jhZ54dBKeZYkC2A1TtWU32yt
vdZbZzLP86cSIUMBiclnu2mfL9ZaVar4a6tYNBm7OAtg7BG/2yTXafjuf5P9mhbdHhJT8CCLORIE
1cdmZLfI+K95r/FDaRxUhHQ6Rg5PcAKgX5Q8wO21W0ap+KIqcLf2yHYT5rTA4zhYzLlZiAVCMXyA
5Sf5uBdDIyJPq3zP/CsHFsAHuloJ/P1B0c1TYqaKJAdGQBv2Gn0CqbhMap90l5/I1ha/1wDru5kB
09GsvAlG6QpA3gTdq1qYE6oPXRgL8e/TI8AxnQ3Xsq400YR29M6eP6TI1xJl/5f0CZ8ngosC1J29
q6cNJCjdTtRCM3BFWXWl0KIkHkIa32i+HGrKNUKjvISmISiwonwlfNNddczYkPx7dur5vlRp/QmS
ovJa/wKPwsJo/po+f4j+JwYHSmAz0SKh7sLnO8graAq5jMLh7mEqsxyCevvfHD33pyR/AaK7zU1T
NQ1pbaE25BWBmulyLFkUgCC5KCoZi6QpUobv61txcskIeRfwhAt1P32ISMWlWU7ckw+oj8nbTDRq
tPUqp/N7enTlowKrBy1IAnjNKT9+nxfAWNFmxYniLbI3N5tVgXVcM5NzV9pZIihN2x0QA5hE6KWn
Q09k3Nr/f8XS+/2PxOwBmiUiQ9UAZMIzX+It40SLGJPBFGEo6/nBuncCx06ea9lRitwKyeVBqpJj
KnJgZsx0sO08N4Z9b56ZJsXunUslOL23S/lyv3TaEzPbG7PwebKGONfVrWrD349UC2nnI40wSMDz
5RjAhv1ykSL+KU9S7KUN5nOxYbiA5nCSmSZZ2Amz6zjf263/5e5xzDcJQLvizbluxymhvq6ZubRw
s+HWR61uF7Kxr1f3GUx3JmBLaBdIRN5+jNVbJ/qvDNCyy2HmKXxjq9cLqG9S7yKj62Mu9Ll+pd6I
qFNZAoGodUdLTcHXOjTLTcpDZzqEcB6/RLqCEWV7ho2EYv9D/AuhlkjHPzyY9pbQsaYfSj7PWx6h
qCX6Rb962p16vS0Krw11YFD1AiNfQNc7G+k6auQ8UEDqVaYlFR1/o+0CXwKFSDpjGGiA8qepdPEO
53QI1ZfJk9mpoZ0vgdLDDCljoiSlq+j/DX62jH7OxjacHo3UyZ+SAIsMvbfUmcFuJANF828cz8WE
BQTjQbxPVTdnWx/PINkP/i3LcXUbAdG4whunvhlg5S0qBMI2xuA83JejmYyuU0MrI8mw+8ACffPw
dvWt5AIrTXTJJi6wh4wuLYTLMRrLxU1HSJqxuTaQILNjvRPBcSF1APpjpR679IMXRVT7m3E7IgC4
YQAo/oqH7EAWF6567b0CrCd/KDAItVdWVjxsrJ3Ww7yecAvhrSKMTWuGjmw6P0wMDBeu+L6db3Lz
UplnYFMWKuOz8FtIdRVJLBmt0vv5wuMg5PGd0gYYax5CriMG0XdEpfRTjI6yOR2F1gvqvjtUrA3P
eUoxNQrVlbIveILOlaIwltQwoBA01OhU+d6ODjcGpMXA78MAEKxjyPSTZEsU9JLxlGjvGfsnEHUG
IsLHolbKxp+bFM/I8k9e/FC52v/9DCGvzCPQ3TugFB+rhzQ/zyf5BYTOs3i70WG86Tr3q0L+lgzY
RyU7UNbRC4FpL8g9I3NF62dmLapI1gngR7Hrd8zDTImbVG+yJ2XzGyOyl8qVNjA40FmaQjGhTF4H
MvhpW+rZdM6EyC7Iu2QtzxFq2rxGUlUkEWgJFDmaOPM467d/5wW3QllMmbPEWU8EUKfIl8+CJd8Q
9isfnEE4ksCDZvSY5gmBSj+BmHD2fX/xkm28fHysCvDVY+enMQIn4sXB36F/FV0jGTAvKhYysx3v
uvKkdTifD+AZDmDYIs34yld1xtINcta47yEGkPQRk0cDk2pHOJ5kGesU7wzFnYhL3JC0AZHxm4Yl
j07gvQ/3GM6eOdi2TCp4TqtQF+JPNcTXXjXfCltTeTs0fZdEFYZx0VOzwi6arTep3ZjP5B0LzjcN
sf4/gFmp/cjvTAxnp4TGG+MHIYz56sPGoOxLDYjJlWBmvwFvMugUQxCNbRZ1LzgoTFD693ZWO/L4
99ICG+qsIpquNngJHx98F4spG/oWpI637j8XEJuXNep6tB+GKhWClAOrJaaqTc3Qnw3YobFdtZOg
SY9D5sVgopohzTmsonPX5dSPIK262Tr+MgfEdeuH5PxApxrcgAhAhniMKLIEPo+Chjqxtepby3CS
fHljoIBiJVk/u0NwFxP3e63+0fHmokp8ZgFgvRyYsUvv5jOdVkX9AUWOdiad5DCLoP6H49/wf6o1
PYo3fS/9VNkTkG6wkCEUx65J+mcS8DDRvBEHcbFAyKWUarXu74YMZrJPkdmPNz1d+A+x8f4bO/EK
XB49pDVbCuch3LSHNPTcdPQD701I7BQH+/VOUwIpPHOHnV80Tf1yKxooF+tnDFp0z4LU275epPfH
3tJpw/TFTfv85Xy1hs2K4hQydouA5CM+93O5e4sRsHNb8Sduor4W10Gr0g/XTaWdB3595JBUDw6d
mZxC3Ix1EcqanOnj303L/8ti1hExm/khEgOglx6KLn38BOxxb2TvFVXbyor22iWqqmuNgO3KAIUd
5RjjIRf1nSGb44/kazvJVM+QuoT9VyTA1WqjgczwqeE5uedI0RhacalOkWe5eug5H9pTktWfZpxK
Onq85LcFNX/Q0y+vHZhe89nIka6J3F/ffSho/l18MCf7gjHKLBUzHniESHvoAipsAKVMFPsbZSpe
e+unE72gBV8ON08sbldA1dTOs92W/aEptMQHqi/CYAz/HkDmTw45HsfbjptY6+R0bGrMqHcCvxAS
fsv53jRhC1z9EKxIcNdmHx73cxOqb53HrREgEfDIrT9X7/W7rcHHpcPlVRj0jBtXC0U5tpC5LgYc
qOzLYR/4VZMBTUF8HxY8bLABMriwV/WmpQfLobYhyXOm5QQdGTTaa9V+kEwJBIyO6BIzRsTjVOtt
bS5yyqiZTe4s0eRRdIu2Xl2LV0FSiIhdtNS+l0kBvN3riHh91tMh/WlHo6TdypjHO+3iTtdKtJ8G
4ambuJ3rXjRnMuW6SI5Yd3JbPX3kv/Ro07jRdfSlyLNZnqjxZaLzBeYLbGTv5UlIZ8a2FcV4UPZQ
kHwqzarDp9DDptb4+M6oHktJS9clDSqf+317nTVVIdMpM+XyBe5PCm60urSv+QefJ+mx6Oh1eD+J
ZH9Phpvl6HjCmBthKQa1LIMyH/sfsn+9e8kZ7r6IuxJO/hAsW7/ElQML3Y2t8sa22Gy0474dlNlk
PfQunjKlFCFxI9kNpcce+w5ySqKyz++cQ9SmaEoAhAjoDLWAyJE4GvuY4FDKmzrV8StATokFesc5
70y3frLNoxg/wy30MPAyGnKLPYz8y18Qpma6gaAKw8Ybb14bJIhoRipW3hkZJS06u20MkatKzIwq
VSNVJaibH9bjIbXEYIpCndW8+nmqGeTdhgHNRiCaFI2MejcTj2MmAUyBgvxZYwB32elVoPZ552Ac
A7SnqnO6AkJ1jfiSt/uclYbgqq6FZ6y6hGaibALiDH5qwK5kOshcLYYjtWMZK51KU6v0YEtqoWaQ
PLb3Kjb9kpf3WSz24dORSW6qkhFIHELZJqdZV32+xLZwLg0Bhm7sBXghDAMFptbI1G9uRF2gJuxr
3e5abRukj3KxveEz0xLW6gGW3SfARXsFibvj/ENaAxYLBZoULKdWrVdGJuIcfqQimMdGWtazLDxt
gpqPXg/dzAULKauDnjSQi9bWUSXF+A7TobaFqawAd2MihlJ1Zq6/TEqDsqpXXkIDJGnObAolc955
NPcLnqw/2EUY6hc42+f0QSUQeTWFdlPjN5SFVKOIhMzMECHzTs/3FhJmPvw2Owqdb15rMKAyO4xw
hGkr3gQilvsFgnpaCj38I32wJK1RPZYoK+A1nKvSXlBcuqSplrpLJpdNNEjJyPfb1+7g+VOlUpaG
lQZ+K80cUV+ftg+FFhwvHLdQQab3Zp1bl0uQZEboYy6BilR7jtdfcmQT/yZnCWqEIqZt5KluOn4l
iypC2s/eMYoxYR5avU7Gj13seon/odtj6Ae+uv0w49o6Mq9MG+ZLjIOAbNDZW4JkYaNolkN3Tifh
le+EqnGpNcTt3waH/LUnq90oN/mP6SMwu/JqQ18X5ACJiwX3/DfpKqNMG1EZD8z0Yjgd3pew65Uv
rDzVZq6Hd3iy3pr5KsbVoNyQ9tYt9JZxxbLvuCbxp20FN11hKl0wjyxHmni8+57YckLGg/nieFxT
xCO+FZr9GhhqYDgIs3z+4aO44Y+BkA30wT7nhPjnnCBJCo+66a1Ium559LI+ojZZUwGiRq5ds6NQ
FuUxoSDhWq2U1O24v3oM3ssAa+OkQyQcSK/tI1oGqD1ycoE07+mzyFrr1CycMUUY42MGs/vcLViw
yhdVo1Y5deRWE7E9g8h6trosEMmrobd1W4Duf5uwQjnskbZKrnSkVPgO/6jsjMkxbr9sOFBAhwV7
idi9BFLN/HPynjmgmlSPDkqevhJdsdT81AtdwawXMveZnp/PKmzLuHwMZon+GN1NJ+otrUsWFRY5
8y9D2ewhpJB3hNqYC63uVcKTQ4GOnzOw/ZoWDV/4CTiKd0umP29Fp955GUA1XbK5gTSrUdTSaYbK
onkisXYloSmtTU+3ITGEz0zaPaLho3Cha4hoebRnL4TXH4ZR7ebfwJL0Vo8WUzI4064TJ26wUIzJ
pbyhDR/cuSTtKVVtJI2U/+K784OM0eFgMkgmoFrSNGoPzi9TqDXz3Aau9R+H2axWoIsmfnLaYuV+
TRFaJP4HrULL05LHOrNxojPXphQprGZxW5PMyz0m0zHSvB7DRTKASDtw1ecVptx4cEQIomF/sAwM
j+2e5rentktQGgMZw/BNO6WI39MJNq7QAEHdIdNTar6RMjAFVT4wrrU+8u7/Xy0cJgIcVYTdFkYM
vCV2RGLqRbtQ65xnz9dS+7yps8DfpeML5JFo1rjJWRQgP1y4EubyLblRrDRIie1dlwvws9kvOIQt
nVGQPR8GK82+BtpnF8MfdbTQ50JUJlznrhlFW77N/kun0JIDNFV93dDmr3peJaERQj5qCVBa9GeV
PY4W+rECyhFoJdNkXJY0o0LjUNkDbkPAeupIn52UI/GibrT7Mr4cLB8vakzZx3AUP9GhaNAxp13i
jKDa80YgvarlIqPD5/PEKzEV3C2VysYD6BFnEanCfsGb1NqI1GlTnhQequE2VV0OX3KH/SIotc/I
P0WbvGcZldncfz8FLieioPr993TA1hWqA5RYGdziCPnhOjWIEo0QELWwmR698pbXSjS4vQ1dbi8r
p/+k9J3cQtby+nk8w9AJtL0wD8RG9tHoNp3smbvd54MUFTMDsm8xU9fAt9z6Ao2FT6XM/WDoiwiD
0qRq7/RVpGfCcIX0epfVtb30uXwYE8E+x0ul5C1UeplnP4ovhghpwRf5D4EoCqgAWJ0Kv5X8zUd5
Wa0zoPoOnFEuBmHbX8rr3q0p7zvKQnKgvYOR2ISW9mxEIFSmzca5dF7FT7mudNqsipmKwaQw3Y3R
Pp6RxrWAI9PZhA7jawtOVsyItluLo8cnG18FoB5AubItNvIsNl3EMa2KjjsBk4lvKwxEnLksNz2A
+VEHrldPKTBMQoHdzu9Eltsp/bIqPuRuGC912HBAIhw5f7GsqtpONsPGw05pgLsyI5u8I3ygOrWs
VLEfpAwqmyQaQ4CW0Tt8tXA4tZ51EJpOLugL+z3HqFVmyVpZl3c5uWiaL0ucTFpWvqUSEzsb7FIq
+eXE2vRk3/vkQgLStL8Lmw6SmYuR9Y8vPWu5hwA2aAOtNMFyvmXDXgu3jMFvkqxG0926QtWUyn0r
Dh3SCpl2/LR1HSDLVg8FVmd3unfd5Y0bIbhdeAF+xgMAgdXpuyC9NYhiXO8gyUEMaT8t0dW6o+I2
Tf5SuZUanw22SCtTbgLP+cLOs23GN/wBO0j8s6N8WT+6qCfFFDtCPCjEDR25SCKcEcNkkXuXw1Nz
jgsy70FykIyCLZQkYGNteHjaYb7/XuhorYxdDHzIJrmwtap71bzOkYgi+/81pomqYdUoz763yksY
Rj7KhXZiPl7bLt3kWQDQk1aJzSGt/4bZoH2vRwf/PS9siSlJd/ZKLuaDBIKZBq01R67/El8lMQ5O
3MlEEJSe85uZdiHDkV1AFvTM9ujWyDaxiWWPSKtttlQqoS2i0fPBjJM9T92T9uiZrNDw5AQiKS7z
ZKBBs+8glzO/v8Gc0NIdS72DYMhCYfxhhWaeAricg/uCKDqOJeE+XhYyGk/6xga4oHcSu3vzkMN+
xJ8ZpW4lGTzrSe0ApVT6h6gZgBBqDNkkLJjOYsrDUmoM0+siNZYnFyNp4seuGIueSkIPqygXqMIy
WTRNcTWQ4Xyi9+hOyiRdpoN0CPHBeMzTFvSXYPk99vlbJkeR7Vohd4wSA3o8a3WVYmUswFvbqILe
BX4xonBrKSTfaXQXn2/VN1A9TKbmkF4cN6TNfRTC4/OstCD0HxgxTgQ00N+Xn4l9O21ijayKHVC2
YRNsYkrafvZH9d1N4lYYSvIK5frwvX074VdLI6CfMSLgvEpwX/Db9Pb25SP9/zy4MeKjVVMbtQl3
t3c2rDU1Y60aUF6+jVJyePxrhp1nP0/DfkwFQvrYeqD2fInWbEG+7Ssk04EvYXka1p9OE9yOd2Ru
sSx95SwexnX8YwrLcxx5YvnbQNVnknH98liFvYVl5Z9ewNQFbHKp/BiuhBhaStpfZRa5koAn6+Nn
8VS3uWiwKkcbo9dncRwmbLXFJi5LI0vFo5vBNd/CySy65/HR4s3nYcBfyA34s8Ulc9+ad+mkPVk5
TNN44kBig6zyNmPpL/78WNC1KN9aUqjZZGJjKApsBeSQGWdtPX5uHxU7GQYhLzjn+k/i54VDRDFy
nYLCQRd8a94VAyLNPQTraI6hRddXKWLMQHMrjTQJMugptTw7j5GfgRg2h7ut5AUs8F1iw0v0DjUu
4yC8/rfA2ovh9sunztwSriULyh/tOwHHP+IOVTAkLp2MnS6aPprvVXHAeYujPmoSX+wrBGgETkzy
64K2Hvm22KnLobFyVT28KlgF3wIazx632K9bmEFt2J3W44r+gkZUjueWnmzdvdHdzeO3X4sC/eMG
dYmAHNY864U2JOcb5ZkspwjJRAG95n4B7fYZbQ6ni+/SfSaZyr1sUV3mradZuem0SHAcTA+pgo0v
8bXFKQBNEQ5KU5acfD8BqviJQmyL/onKDJ4F96xJQbP2dXpBF7fCOtMC/GD7tpnEbgg1pNt11n/N
HDIlLkcb9U8+6kHajjJp7VDdwMp0rLc0kEFgAEVjssm3lCbCMrtzbsh11nyFfC3TcS5hTJU+J47x
ktSvFj6KuHKC19qtavhnmt8QMYVWwYmiqYs69WdpvxEK7pOaqYulZi20SnLtwfcS2YMzrAeVXNcS
l8+/YXWipfq3fwtICEsYVWlC/yFskRsE22WSodaXCIuXAo+wV/RvlYNB/TEESQBPnUjQEjqQJ1gM
pwiDIRwJAqo7nPxaGIzchwgnrCk5/21YpKV0Ab0N1ldM4SZN1YdxFJecMP8bzceR0UVhKMlOEZ/q
JPmWxDj/SM8orS/f3NFUxDc2U7AC3HmJQBNAujw8s/5+aVWPkVllnQKsZm84Gp3aC9S284/gHQ8k
7jz8sbpndP6oGKSxOShcdcXbJMP6jH43xPILN3swu0W40bBG61ok8moD53IWfx0p9pvN/l91QMMA
gkL/lmKI3URRCzZVN+Ac0ZRodbWWwl1q/e9hR7ERaAlfxu6kKHSVjTmF/yRKOWeRIhUFgd1e5r8Y
mapp8s8K23XmyThZe9flMVbucPRErp/BZpJ7E+JsVnR45DJmvqAWHUEMilc7cj8Sc7sxRmQxDwMx
ASOmpP3AM8kUuDANeSiqfLO+OXo/5mKxIjU6eaaPjnz5ESWFQG6Ue1TbIKqcUk/JiEklSz1fLfco
CUz37145C8+jy1JeFob+UR8VbBH85wKZSGFBspOLeHATcukWWspYCWH1hHHp5/8XuowS//KmUFE9
/OsXR20A4sbDwG/2jybGhDhrk1kJCSmeKpHMFgiHqO5WPfrsaNd5/j+FNiASGij6K7COXnMXfR2n
gpQRlD/qnp2+7/4Hpnr8ppKk33QQopWw0VU0BiW7NwqwTbU6YnvZF776GPSXT2HiCXcif4768xdR
Onscf/91jPXCgnb02QrL4VBEAwiGyPFPIoo5bNFj5V1Jj60Byp2MDTfueZy5ejg7TzfAiKmLjk5E
58mmrR0PZ3IJxHe6MDPiFTQ1vpbOlocBB0mKl+kJL++YFCzngfL8ZLTyHgmtA6/jQadLBokc+3Ga
sUtB91ihaGY46Sy6vt+VaTSAgBtJyUfdi9xpPKqT1k10xEUQLgI/EfQ5Ia/iZEMX/SXso2xywQw6
cuilQlWbgZqr1JrWHQ+E/JhAC/zbXgMbtin5KHbsvx7+Gp4OSBdgcMC5A8YQaVvtyVueQZsIWT5m
iTl4M0esb9ZXbWulYTbfqVt8ECk2pEHisPdt2lvpRhSXyfSuM+0mrI3C7llCroPLTY5qgPE5Uo9p
zaMJ3WFIsMRqPsamIIYS0oB4VWOv88ZO6uQIq39V+mLeOpNEv1XLaOKcvjo7VlfUsNCcwiTxNBmL
yq0j6pArsyzX3C9zedO0UMqsHiiw9Ok6ajg5z/KrF3HXpqttLFeLjQlIPze2Pu6ZzvTrjmc5TiM9
fKP1Oi6RLaKlOT+km5OdyYJ/cEuM/jWKl6VPgbEqCV6Ypiq0K034MP7chYCLIqKs/HEcJCW2D6Vk
g1ivUqUFGcuwFjzFlO9GJmduF/R59o/7LSTtZt8wyZALixHAlkMni3pl8rsQmxbuQ16Oix+XwLHK
nQ1KAxNQ9G2LqLvBAZNd0IRYeGZGwYvjsECaKx4AB+ne5jqblfogumY36YmB6nj9lkxMs8Y/+ycf
q52P0eI2pHIn2w8B9nWAWe7ZU2q7meWIBC3UUMTvffv0wfwoMfew0mCEMxxd44pUgZ/vKCfGeeSq
OFksaw5sg2KJrz5BW0vFuVkxGI4vHFnSJ/cXR5Pm24lafCTn1yImb1P6L45z1vRu+hoMaOSwEYxT
TXFQuPjRVHgAWirEOwDGYBCCrZVN94Yxalu80hDZomFxAjXZh5OCAXPhYUAXzpeHFZq/dpJd32fV
WSVI9NJL16i5BAvytpAmGWwb7OpraxpxQGlDOWFBn4WIiAid83oaWJYAW8plybzF4vKpkbchomEf
vU1IyOejW3VxddzCsJuK5bBze/6EXFrHGm/dpdgaKuGchK7nzGbN2/Z/lfey4lvKS5uQ0tTfhYHD
ESMNrnOr2SpmAOQ67B8WitvWyZ/w0awwIaXcps5rZHSJ5GnKYXvf7WbQBzHEHRefnZ//wsMhqmqP
RjggYBUCvB9h1lAIMmPCyikbATHDvyRoJg270WVJiL2T68KtmYT4vSkMphpjcxjJNGqdHdJ1U+PE
FEfDbj0xaJEVzJfKLRO4gLpBadTepGjfOdwZ8u65S2xVPZDMdRCoGYvDxm1oISSGRQVb6M1P9aK6
yYhLmW3j09OmGulkpdPdXruu+i5QyfG06VkkVUQ884L5CdiDUGIX9RHXYEJF6YAoPmWMCGiPIkUz
rlnNr29PfBJ0kvbOPm8zEBdW+KX0USDJuHM+AgwqhB8IG/1i4qG9pzkQtEVDHGJEBBA9WwQJF9GF
OnhSUFg3hW/VrSkPHWhXNxBv9NyOY3RIW9ESgr6xAj8tV7TovNWKUBxS6+voffObjj0Og49EqlOH
V85TyIOyL9O9nFKITZxrKBGhdh0W+/GfX+jnZxVclSHtQP72neGk9Mpk8Uxr3Y6aMNKcb7gY+cwv
e3GxaZyWbeYfYP09/MDQ6dgnlz/oIBUFmk0i3/bNeAS6pbLjh0rIl5Gf0tEqt36fEBNILpi8pxsp
q21NBUYqvjBOhwQbLmvT9XPC/TEwZCJcf6rhlnCJ25X/1QkK8USuJHEoJaogcFn7Mjn6+eirbFfR
sNUvxSQOMzQ2q4cmCfTd+kOlOsgUQqS7W5jLOG2zYarh/c1ZvSSvHgqclCqpxCe2tYz2nwogzY4j
vJTwhYvD2zc4teM4cGCM+tC0M3zP+mGlW5r2sKApgkIRr/LfvCEVxEL84EdFBKlGfQBGTSbT75JU
jucpTvDDdbuMjk/rnrudHcsKNN5m4Eqe8YO56+L0AIi9s2Y3XWn0NBtxh7z2Su8RbeYUMIRbV/02
BM589f7hB4VWjKFeTW0ZXvAx7NzC8C6dwmv+FBF4N8ykUqlTovpfwtnnl2fUHda+V+CKtGFs2o/9
J7i3aszJGAOlqJsov/VRTcgHxai6YxB3L73pONvMFEMZrtZT57ayY8wVHY2Yzx8iViAenu/4D6OV
E7YcydouMW/xmgoKrUEyQSmnXBxTDKzZOdvvnE6C7AhAzq9/3j8e4Ov62sdDI6BTypBLUaAjg67Q
MyonsiSIWJWTknIQXLv9hazBSiR1cO/iq2APTGS3Oy3YuMoCRTagd2RDaUJvnV2doH0fbMdZbPPj
lpb1bLq37wsSfRgiYU1E0gvfjUI3GeHMtA/NnTB/JHjd4khFxMRJXOS0PJj6pB20h/R1CKY0JkIS
8zCfp1Ba78YmpmATQQQA9GQPfoJEDZTnf6GwFkxsbSBy3//3WLXlCaHwO/ssZC5oNJeRSIUdmc1f
QsPl0qCCpnTDLVA9oL0fqnmxAZ4pvoRAeHWATqTkgwrCcCFd76nbvHT/2IRXlY1gP3BSurGbJPWT
dHDmS/AjjbXuxU6A1uXy5Ld2WK6nlzcNH5euW1iPl3fWtneKXOajDZwWVkxZzAbZKEjw3o1AD61P
Ev6uKACUI5IEa4hkuuhl1zydXbRk3YnHNag4NPMm79NfDUSr4ZFlTdU1jSLh/MiNdqZrmn4daAY5
6UJ1npCSpk/z2GkM5uGHhT1Q5DbSPXBSvgqPIR9fbTu+x7elYW09oYpQKluDGUPuCblTSG7dFE2E
pSaw/6kILV/nGyugupZAufaBvDXzW2yP2ibQtpiPF4/6Q8irQmPqmYlPOHET8XmRtIRFiSIq5JEI
Z+p4fkhtTCRhPQ98KKPZZUDnC3ZP9EXWSojusNqcTFJJMDJrhfFC2A7rl9oQqj2WFpNuBS46Yj15
J3v+D4rQx2jtafm6Dk+i02mFG3wEGKTEobpOThitujHGn4EK+aHruWq0X+dCcnupYtedmd45fDRY
In/CB0e/Fw/RJYeGREWmggKId8Pa9yPkXx/a9baZoxhBOp7QRLOxeSvlck9KWOZ2Lh3YSgaY+8u8
sx/K1jbUR3rF0UH3juoKcaJ/mOIPKai4XHG5VlM9w8RUBeqmqjjZjXpmh2YPGC3AuyybbdGbyJ5S
Zqwol3ts0eu3ZYH9Uq+7bubLZSIhvrFG/Wb2MRd4IqJr3Wj6ocNI9bO9bxSqqthMqSrV5jYG50qL
IzY8gXGvahR44c2crEL/rj3ALwweuSZr5P8SIUnv5JlfiwjwdDkeRvu74BN07+Xe/pSxqH5rgig6
eRfRTRhCdwA9KREnFQQhQqnY+rAhvWTzOrYexSSlL1XY5and80lDIlag5tzmuClQCs83EXseJUOA
y2bhj4jw05lmmUkVZkZFcL1w9IGS7n9vxf/lkjuyx3AkHE4Jue+0Zvz5QzIp2/tARJd2qacCafvm
ctsQ5Weog7kEHhHe+Lt5PslxuUQvA63qzwuOkH6l/KH37FEBUM4WfGfcvC+D0zVkutlOyzhcutKU
gYqCx1GUadDm6ulW+KLvgGGeIwX2BQjQdAOj0S0htPg3pgU48TumttujO7UaT0Mxd3AGTqVxnuPw
tmDOKKr1dkotsNnQW6Fi4+9kuBYDhIJyOCQk14hUdYbqjfgS/eevICx8YE2fYMl17KduZ+VT8hJD
wAXbbMzTryC8/jSujLKBgIdIaDMpA/jv6pnpcJapaBNw1/VKYgdB1QgiYWrNWbtzCIR7dahgTmA1
HV069SHNZKDgv1POLKgHFOtkp0EwIttcGnSJApKrFkbON+JZatIKByN0Q1p8yPUtsjhA82/9/bn6
mcN8K9qqFjoV0YOH+j7ru7g0FO0lQTnRujAUUf+yVHzrmGjoGepc2JeC9ZTrE6Jt2Z5/HF1gpuNn
mUkUkI4/MP2D0wCETgizAHOE3Jaus0oxDxReg0KnnSTl81CrXwQFgq2ubudSkftiHJIPElgzRFt/
Maese5XpaRNzXOkF5wTFfXFpzn++lrWTGTch1BV/c0o0eaexnkoORaAi/IjCLA799BBfano/gKP8
ArHhQ1zHF66CFtOQ/oRMzXgdTJJsaFi0/jqmxxRovFEkPPgbdJR8VbkvrrjumhzK7V6HJJO9/lDP
l2NFwoxD4lSmsSwBk0L3ixprZadoV6Hh8+NXf1UR6SaCHfCAQ4Yx6+6Iv/IJ3o0hTnrItxW6uoE9
LgjuRJSWngJT49W2SEMoO6HL4yADSurJQfCcyawlWKUCylefH7q34jABleuKRlKLCuUifSXEhdKC
JFh071VdU5mZqQCeElmIocA7vg+Bz5+KEJX78ZESs1Fwns0+f2ouUWalEgGjnHtK8t9fyScFBhf1
I8adlVxmWrRVpg2YeH/A2WGo8j32wcwO1J1QXDdsJ+k3E1ZPxMfz6IB5cYkmHZ2bvpmckw5spwEi
HEcWeVb7X0OC7wb2SS99k7PwXw6rjCiVHYzKSLIV1u8nenAfRb5FYnhOl2SJFTu+6vYwVfjU1UrD
hMgSeQm9sserd31Ai4263IhgUhzkAeWXdG7J/6bVDREaW9d9vPOdWOBK4zb7PQrIaThNPDiQJV3l
J5wrlcmlbsv5n9MFdzahYQgWqL6izjgGKbn5R2IcXeZMa4TTeKDYvB9v9moLiAU7ALT3paHVPD5C
cjRMD7vQ7UxY6o3HMZngyek97DvsstCldqMpRRdnnhD+prNIxn3tZR6HU+cZzT8A7ec/QlXNjK/t
aNEcObMvgIluZD2yS3DbSSyjHjwbt10tjg0NQeNCHF3SluMsd9Cm29Qr6xr3ao31JCyeeD9gUlGV
CFa3HUkCnQVYR++Ht54R5LaMPLziPaRy+lwgzamBTEQNTe6TlQzWlDondVXgjk9b1ggMbX6cPPOm
A+BmDh0Gr/PnazcJOp6BQdsFNnyrC/WmmY02qeYV/lAE524KDzJItVotGBQ1jdh542s03p+GTtqI
tMZx1YsKDAGDPJHW9hd8lQPj7DfRub9jr1ujT6GfslDrtYfx2scIzakib80Hnr9Qdm10oVVuZwYB
khEUjsKxFaV5Bk+pP9hjl8YpWjoKldjtBRX47PDuYTqvc3m2X/J0MuWSVw+fIXcoi00WH0r4XLcW
rchJBrTYeJlKLsJYrcnj2O/Bkb9IwduHjuaxpKjmh4PlMWyCtYEgcRjTdRJj6ww7dli1k3MX2m5O
WpzNYJCCImFOjqdAsNzk1RtKTJ/HxEFvoY8YExFzxT0hFlA/VI9BMUAwQNb6N8uOVDJ67PvmPvSK
GA/AICV1kgVi6E3AioSV/aavcLen7NW1/bMhbHVoIzDZzTiWsoN5ktXeck7gftd0WGJt2cJAaj+q
PTyqZibTYzR5EoKuu+7Ajo/D6iJkhXQF9/gB6qlRHchEBRjlBdvc5c/DIv9PaQUIDIrLl+D73dos
byATgo4RI1Q3yvoWQWlTagQcVb2U74RrtADgj/kk/4H6yhrN8ie8aTsegazTiW2FSMfB441/lWj9
CU1AF0mre2HGQ6GJ/0+WU8X8EmT807qWv/Gb5fxP5D3ZeG0fRL9pJKABuAsf9mLWWx60gueg6gBi
rbZv9rpP4JoS35SgQE/L8n7gXbdCCSFAZXR3AMxRCE4p/Wd17Vd7sZjvExGeQ1pm3AV/G5KAKcJC
x8p8NKRRR0WFP4pg22NhUffrlK6jjPHmfLHAZA28h6BSVzwEhiko7Gonibc5b9p5zhdWtBVsKlmf
6AFAdsZEiebwE5/NaF4hXSSQoBEa8aolNW71Kd7UVH1qugjsL0ZIQ4TN+YYOx8dHUdtAOgt+kRaq
ZSEzGrxP38hf4d9UZDsERZcBarh66+HQB5cGoTYglqyMpV8wty7gr5tjdeEyhajRiN/DUYaaQShJ
hluS+F1XdJ+oY11YrL7OQ933PYW+2TB252Uv6iGRpc8VY3QCOb1UuENZcQxc8t3MDZaDgN4+sBm6
9AF81OWWE+gi74Gi7RLZk0akQl88rGqgzEWkJUws4Vs3Oyeb4iPIhtZnNwAwZC3jFDY2O+FioTS9
ZSCDgnFA92rJZh5XqLMMlvwy1Mx2YfdrQ08oepgBImXojm0V46xA4rn2kKz2T8ML7vPd58g19zk3
Mf0vUTtOAiXfakVmJkK0oyKOnbM+EHiTPNVrtBq3SDjBs41sWLhhQyZDl169t5tVpEjpbv3/GzY8
Oc8leA76JaFcG6cNNm0oFeMY/Nn3RS9HUCYzhaRMSaNDR+wqV083+xUTUCC2ENWsvZvI23jyiXVq
Xr5dsNoqNpQ4PehXw4PU8flNvf5gmoyfH08oChuahmiMjmw282krn6Hs26GyQwoG14VKwCa1jH3W
0AKHVzihQwh4i/aFr6Bb6mxEd0RLQJuwnYI3RQsODORiDZx7Wo30mkjuyq/0dS1wtSaUSNpxWAiI
uM/2rFV8aEV/WQR2ps3rr78tS6SKZ4/RGW2WdW6pKhAC9t+txIOCl2ZS8Jp3jLQT5yvAvL65eYUc
n/U3LYWGr6dApGcXueQiqS9EMTOXveDOM5tBj0JL8OFsZ0hjdkpYSQNs5HIVyRZsRheQWnejifox
5AqBr9l3jIcSOpkOUMPmuom4zBGafDYJChh39xk62vf8MHmv3NW+IHV18/NZ71AmxmXsZQ4emJYY
OFJvzeb2h4uXNdwTHnj2kWigO4wjc5Cpakasmil3W0dJOYlJrMmZ0KdB+SFa2Rw8AFhM8VNidIx1
WBHJVQPR6L3XJAmT+U156o/CSac+9xS23T2dw52CiJArUaaQN9pKsxtPYjtT5R4/5HDlAuF4jrnH
o7Epkq5psxhRT0uuUCc+NF9ZRQHUXcuxNgVYnICFDBohbVkU46Q0BbIeX5TOxczae8qJL7W4aath
ysax1Ub3t2pMicpffLrNXtgU2i09rrFHuA+cFizB2HgUiBCBrbCJMs27OMzBA1wQVbsCa9iPY5NF
0ud/KtIKJenjuZqfQG1hvo+RSpuhoJ0vWgHhQRL3UrxDziAwST9pcg98bur5H43BLrWgGDN01Yze
t/rRFo2qgN683373F9oDBMnRbebpABfdPA/44Js5EjcyHPJApllf5msYb8erGSa+1Co95sK72gbv
aURboKA+xsy364mWJOjC1XycHGq/NAa9QHo21oi8bKGKFGhuwF4aGMH4w1iv9lqO4hjx83yV6E0c
2hnclKzl7yoyPemZugS4jkMfHGEZ2vR4OVgfmC7p6p9DDO3zdeWSKMkdNqrKZoGDsoPYWd0yLaD5
vcOTW9CkWxtBQNyR5iILmv5EUEOFzVm2lR90VImcpIpYlYDD/COLVQHu3/z5WO+ODDV2JLnu/4g2
A/n2bYEYXI3MacnwzkL+kaIqymIT7Csx8/imOilAJ37c6Jb0Qh5C1w4uUsNvhBFi2J4sR+CupprS
nPtK7wL6UQWoE+3EEVhHeuWg51xY2TBOTPyOwf+Xvs+je4aLblKTcKKAVKCVpLUgAusq+m4DsUKm
OvQsVHfowP5MDITvGCoYdMSG6cmYZS5KX9t90yTSBl5ACYXu8yrowWIjop+p5HjfyedmbrrfdsR6
N73/2CqO4PdwHvnlQRr6lgq+UwY7pOTa58BZqHHVFFGjtckdj57wSNq87PO+30YbaCibs/nO3l+n
6C9smxrTr1g4JeTnNqIs4Re1m8FchLnw56UwI68N8zWlNVlZLQkyhnYaaLtxKJCuVCzLUeLVct7E
CqQa9Kcq8ydDcHRw5DfQHru8TroWOy1CD4nHRLnry5ZPhrCsG8+pjm3QPVEpF/IXILO6lk2OLkoF
/KqGvMer8epfYnylaz9Nwt3f5+DfqD4aqO6UhYly6ZZavrCpMT6iBcsyodgys7BYkYlz25AGRu6I
NgXbaQ+dn3CQx+lf+YE7+9JyHegoaw/hmpjYMZj89BSUD+5s7gqPKqj21KaFoKACF/Xt+TxXezNv
o22m8WA3+BTCCBX+Z6twh4MBRWqIEuKY2rlxJSycBBikNKEVu1ilDaC0ZBRLugJbQyeHZIFCJNU8
PxpEChfWrWYdq5AlVeYp0b4mUhJ5pNfa+lciZjaDzM+r7+GZJ99DqQ2bJKXNEDxI2ngQJJSxLuIs
jirtwhyg7Nr/kSHZkTJVyQWzuWlrXn5/StcRls1XMFk5XQegBUMDlJfGrV4ubxCcVh5W6oeqv3Pw
gMnXGKp00GdRt2u3p3oUI5OvnIp19up2ocEsVugMqByHNkqoCzVQOxaKygQRe8Z4GJ0dnwstcG0w
qnulWlzA7she+gF5hZv/3xw2bMHX5Yuv2gLDMjpGs5DWe3kOKlqcnlimzi06pIMl5UxPLbXFftjl
VBkILRHlStGVgaEFc4iaFYQklya7LGhKiED+M9f2kydH6K5GwkeC+/CIqeQinUi8qJun0N5YRvtV
K+jnHqE+MdkrzJs16KnVLCDgJ07zhJCZaMS6Gz2c1j+qhhtKEOjJ2q8Y3gkBIGgyeFdmeQwWHPUp
0/QE6QOpifhO0eHf3joyUWWnCMlPiRnK4g482s1U9lcSZ8aKb6CqfApuAmi2NDEfnQ2YzppGrjVa
XiA62lVO3RrnwQQCRiRht4tbtKPAehb3731jIC/ffdcULizK+NC6UTSSjxMqyTW4FbPymJSt7ppD
+SrmABzdKQJyQsuGxZBzww7D/zEnEfX7AVgUD/p1VZX6aJyPjxckWf17p0Kk0dRdU8SA9NXwlIRL
+gj8pusJ+GEAklDIHVxiKuPtfgJaDnehvAwKn8eWZ6UWx3UNQDNZ/dkUEa4huhtqWASCduaKGVKE
Boijz2jPJJaKe2fg9ErBiWbLWrZpn6wUmlizbXWLPcbn9qMmKrcB7nLEnq1X1KpBcquy8r0TQ9Uv
LxX6LeqvK7eKNPeM/2I8MlRVXKp5MYi4cbdt/+FBIMSFRgq4CG9MYA7G+tOi1UjHVoAc8n3285yT
MLPVuhuia/illPL+N41wui2TwFYQjan98Onx4qtxLfiiODmaTDEyWIVGucPc8FnEfnDimWVcJf+5
hAT1LLy65zL5jvJJ0XWyHz8F4o3/zxU5gCuHMIGEjxY0b3h+y0utx8t6w1aEQVEkTgc7qOTVnQb3
6AOmvfw2xdX7MKU5U7NYnA79hT894Aw+i9mwXO7eV/mMn5sTPbOEX8IheicTLMSM13tWjhGvxwB/
KWV9ZC0r8cRaVwHr1R6wS6jC/CDtsrTzihaQ1RRhJIw8kuiFlMh/yurDZVdh3LP4FLvR/IplqKY1
ZFXbzP8XjEAAHqQCdE54VTiwV2vtIH75wc4/MGpnlTotVODXfzLB+vHrKoUyTNBFJFS7Y4J3pSy/
SG5UTUSKUZWb7pmRmlKqs01wTH2c0pzBwMmYWORTxczGQmTfZ04aJbMdn+aBLpLf+kZ3L0+nYRnf
UeadqXDSw5crpxCRkwpq7Ga4PRHZd/w0LYb9SsD7TOIKQPJswOb4mfmk9YQTOgSWzOrEB+4COGq3
ZQKHpdDWmk96EXxH4DvVyV1C1wNd5LhxwJ8mo9sKnyvfY0F2SfLAbRgYRsM1rg4QD1DOtT4UQGvl
XyHJEYpmfJ++69mqUeJQFLieoOmymzu8jJlbZonQ9uOgnOxyuK6Yf4FpH8IByxesJek3/Ge8kK0y
Hy5BU0/1ty3MDQA463j+2MTw/DJyCiaCTp6cEnlzhMgVPAGMTkSFkX00bgE61y0oP5gTZPy6QOLD
kzFinGZCO3nD+e9AfP10KF/C9kj6M1XGM8M7Cu/ychmgoiVesj31C0WTIbHEUbyjtT4cKIlNBaXr
oyrX671/I5jKunVg13RbwoX0TmCGPfHulta1nv9UQRKZDSDkkXLvbAEiT9c4HVO7IU5iBggQoq1j
kuaksd2xqb2723FXVsWcq6G/bMVr00ow8K5rtyZe314qqt3meD1STtQ6I+Fhcvfr6RhzOmOUhUhb
6xi94/5uLuOKLPj6EmirqS6k7pxY9ejHtgp9sZyuI03AQdcm3I0jKAjsTukHiKb/W2gF3SfZYx/s
9SYuJIlwxOQHGXqqrVB+QRlJ2gGQ9hfc7tPoCW90UsUa0tf5FsQdINSNgRZZlrC6ho1GJ/bo7R38
oF/JWcypACcnPo8sWt2VmIyXaJlpY6Xn5R1UDdlsNxXcyjOih3aThLqoCuPVCfGiD0lwuDtoF42j
cSKSwZmGWrx8E6cp+In/bj0vmCyh41PhDwgrSfJM6iZr58PAM+EzQ/LyCv7XjpKMVbMpVolqKbd2
IpmBu7Te3NRN8P07svO4zoFufdROTfh5DsNix0b7vInPHrHuSi7eSu7liVaKgc8vhJ+9ncGowiTb
EkDSIOmvrlbK9oTjIpA0U9uqZL7cbEbYZxTeN/WMfAN6kKrPo8mW552F96X6m0R9NfQGHmE6eaQa
eEWTRhHEajxGfcbZb8CJOGer1iDjujMfg3q+sBvrd7dLTaVnUD7klQP/Mfst/VgsAow3/iD/5Oob
HS/2y5lVXLh/IJ/3XqXdx87LQAlg2igJIpc51qF8TUuNhpW+vXW2dhQqSrvPSebc7ElisJUyzfjk
0FvsPc7VALHDmdSXkwR1Tew1zgJMqYlURAWJSCaLO2dMVm5vvxk6OObYJNPeYElstPlRiCADFDQM
7S0socQJI392sfTvYr7cW1djFfi71xXDSEPjWlkb52TSATudEXxEhE1XisBhhzuV7zTT5xvjh7NI
vWLSlqTG+XnRFdKVcxe5kcZsBMUhlJyCAq8hqSwn8PAEU84OhhjiCwaRPInrQAEi0TcrqxADxEmQ
9vJVzfIv1KRgjv8rDMoA5RN26+p3wojJMXXGhbXIE5VZXEk4g5sgzx6Wr4S1GMIlG9rguxgQAq2j
/25+tBo125mKwFhxXyZnGAII4ZScG3WqmjqHyWWJTEs65BvdssOfiqsFniJAWOpNANevHNBtb5rZ
eXf9zBJ9UBtGuB1rHexqvUhvqm1gFvzbI5YjrgPKrVB3hdNDwl1jq4bRXgJI7REcpb+z5vVkeI2/
C6HTIc451gLLP+XBn+cFBLihgKbZ3ZsqEOXVanyGB+A2GmQW6tAi4Gtt+b8mG1f5xs6omorVZG/b
BAt759aqvtpURk04YyftAWV7tYf+11lie+Y2CTo62SJN2Lg/7ULRFl4KQggZQDh1yCWJYaR2soDw
IJaMyGGeWmNY3zgqQfQZO9Mz0nuARXbesEbZuirQXYWLcZD74hV6eUOaFnqBcLEu5G8XpkAgXBNf
O1zhg2qHRzV8WcQuNWbGatdrI6qRYjFRR96psT5XXFCZr88F4ylSHSlP9jzTJnvvHDYl9GAv647i
sGaXo77VtH9DCuQ9zTmjDx7Z+TLsVHPvMD5T8uEBAGvmVbbnCgL0V8vyazvyQhpYU9Zk9jJc0N5M
4kgn+MtLUU3KNJner1v7LWYGd/Zjj0ErN1EL1/2auZyZwO4Xw83l2u6YZUS5HGsVPJ9tBYhXyeVe
wRY2DERBmtZWRVGOhqvxw7xI+12877ZKcOsHb39VUv+1+bOanDSAI9NeET1cBDkRAGmiAjXYSkN2
DPHLhtY/SRicebgofPka6r00+sxyunWAC2jgC5zvLPOfDUNHe3c8r0gt5FQJcpOeLPkOUfRwKhX+
60U5Hy+3661y23gX64MKhCUikSRTU1Vp6yYVtBKAAXrNk6I4MQWQd3d3WsrwVw/F1aeSqYDyC007
ueMSAsr0eZuChYPX+U28wRTSjfNfMBET5jsBOyr2SIqzdoFdLHZ8atnNH9Jn4u3WIu6ICzrz4mkI
6dfKZ3aio+69WLZA6xN4q41Gwo/PfnzGiBm/JQVYOkwzHtk4Pc/VvKmmbJIl7z0qCH35ZuBVWc8l
7Rs2E1aab/jOuXbYbSaJrRgkfnvfeOTwcIgOcWIyrxwNQ0xV5qTGPhNcrh1aI3203GIfOPL6HCyz
WIuNIrqSOEhBcom/Pb8aXLCCGllGzLh7GNnb0MwOnZaAo2NKFisUTbbxHYh/0odp8zuIkCamupcS
+CPmHT+SDiYElEi17SbdWENU4xSEHJwrmlblltm6jOENUd228V2Al7Z5H09v1wd1dCR2AqtYWaZZ
otAn3N8cuv5P9cmt+myLih8mjol0tF/32ISUpmRkPULP++wcGAUSs/DW+cE1TbZFNC1iNGCyOOz1
N22XXNkB9E3/XVSeEJL69J5lR550pybsG6bRgsZe6kkwzByzfxjJ7QYXE8ltwq4jMODqxWqvDDRr
3bDQYH2uexk+/ma/ww3grSN6n5nDIOiC6wkOQ8jl8tsjXv4tmhoSRvJS2FV8xDscRNGcQgQmromx
2fXBGcRJU0M4INX83IYk2IBDCSj5a0EVmZWTyrrfov83FShliaLT84oqn97AWiujwATHRfCsfSsn
KcKixbtQqoJQIaiC6VOP0N6NIB7eYb549Ag2lfKDbkj9/jcDTdvucKPj/liq8Qqn8k3AFdqwow3p
kEvxzbEhgojOw+17DgKsPUWkAdKnYz5UoSeGPkopUmvgFOPjJC2pXbUjtDso12U00y33W3MUzaKI
FQj0lAfiw4DoZaO+luGLpL43pRnjMFvXhCmP1ipW8ptgSk267g/vKx2LNvb7zZtOuJ9a2PiDbjQt
H/JBAKJYpIrzZZR9y5Hpc9lgIkNpQDxGLGL/49ulZRROM+rxvu06xVlNE7+1Am0gYkVqhYnivzI4
ACc7xhAF2qLqscX+BTkcA2IAUJfA27/d/LLG0GFrUN+e5TwIor9gunPAtHyLRUnS50JujalPuY0j
byqeJjDbymP4pyINgIhT2Bw2Ap0aERq1W27LszX+LiEkJeTJJUFzpsZW+ff9Ra2gTSu2Y6gaHrQL
iCZ8dkuSW4p3rJpaxk18Icklhz3seMbi+IOvOkGxL8U3RFZu5y+EahLy2gpp/o7vQiK8p1PApADs
xyL5aPBZajKCnGIF++qWevTKcMmxYXoK25AyW9kWzzPiHlJEgS4+Af4SfEAfSZnWw7JkQnKArBxJ
hSxDlr6ErOKG5vrodGum2HjpD5nCaNusYE1K9S9AdeWWBYNpdQgvZxWOvIJDSUt+0BSBsBDA9Qj7
f7uBnpypwxlQ0+W4ilSv8J4W4B/np4/DuDno+cpixr6tNF7pKqZpWXtBzSypaDYF7eKKi+U6FVbX
zC67InQqvupjJpVyBiBgmnHIS5YaS+LCLuFtyZ3ElQq3UvkA07TMYZ5Phpv1Dp8hZzpEXVJxgMPr
or/nes5q3OynA/vt1N80NQ14+tVhrP9JyFJH1u2vViqbp574w+PKb64u3g7Onv1XiVUvC8+MNISG
ISmVC1wIazEszisE1kcz84HzzkUWHMG7vh3L5Mn2cm9c+xNNdQM+Z+iOpG+hoNVkVQ03heRUpyyQ
PMg+PxScGSukgYgeqQo4Vr7bI5cvwLVOEfXBkTu5BsAogQy7NEmaBBppXtmyY/d7pITaQBEx5gzX
MO2b3ldjvAy1kCFo2jlP/6Xzbto5PEVHAdVHEJ8P1MUQL/fIU34AvJ1zfeyObYYOQAFGGa7mhwku
73zp00LchR+QQUUiRNK4qJIl3oS7z0h0zd2xBVq0puMauFp5Wvu165m3ckR08/hS7H/LmKOj72C3
P9+p+WE/muywrVy4LBDXEp3Ns6mGxyMfTvNKGewNTWc/HrBvEh0wx18x344h/v+0QvJHd3Hj2sx5
CjKrulsGtaordn3pe/1Fr7vHIs3CcrwigLdCOMB9nrv+7kugPx4PNySX0FLsTz0qJuZqJZMyNzYU
ZjEqiLweuLbE+/kvTll3dW7htjCM7Bb24Lqnrby7a9NmS0Bdrjw4z6YSstSYWgYDs/W1oyqXyAxF
JQ/GPjfJcqbwXUvYtvN83N+d31hJM1z5DuNINI8aKL+YrEZdiYnmeF3xln/whWmHQkDlVsCACcu2
bzfbySIQ5C6SoQWovzO3UsicrQFyUHwymlSAgpdNMsY3jC2Q/vlHYU6IIm3ZKQpaotpoUVHXYq0b
yX7uGwfYAEdxMtufRtAuN7pwt+INzyJ+6u+/z5QewyePc4qQ6w/YUYx3tZug32fFanhaft+d1eon
Cl6F5R0g1IFY+7+w9MdHinE3O+hTctKYtnWOgBzNfchTS1qTKwHTc8XcTXoLWV7QYT4Wm1TLifVv
vpoanYJ8HG1FuisUmP5TWUrbgCKse9l+BVVWDuw144pWDO+4sh6WF4YVlFJrzQOgWNLCC5KSWogn
mQjX5r/em27XemEl0m+5mVUr3edNhcRdDpFzeOD+29MIHtsAsQk7NDSVksotA05Gr3sAyV08vwG8
gcwQBXOcT9Aw+j64gG2dfPZ+S4uRGnzCz8A4u82635aB++tlFE4WHX31fRo0ByilkFblIKuf7WFb
atd7J6DWHQWdb6vHOUZBNcZutRo4/eiNjSG2qoUXJgFqrPc2h0iXNG2UfG2lkKO/z/MfLgEJk4zj
gGd9E1Ayz75RPGoLC0jNBbLtorgZoMg/ArB+0bqdxMEMlzsuoxS4HIY6bjv0yapEdlIl067lOyUh
L0QeZN+wmyTDFrvyBvD2DFyIeJnzw5MiL61Bd5WbXVZEtWtQ/iLC2BPNTNzAmfYq6vWXn7vsUfSK
hgArcw/BRFDVO0ndoRUWct+XkozmQULnizoVwLjrRLmUSVtJ3fuoQV4wzgAO3gX2SQYFh+GLGFRu
qjdfAdNJ6F0rr7ijv3RTH2fFZUn12+Wsr2yC6GMychaq9M9vxBLshsjFw6C/a2MsA2+xUixw0rzB
KA80VM77Vm2zvM6JTojdDbytW10svyqxeLYo2FDAr9f0fyw6HcxmeX1pJqTxkmIXikaN+Gvgs2bA
vCD30kh16lherQX+HqYunyS2lJz9hW7BdECb9+QpBk8bKoebmZQ98V/wUVvU+3zK4bBM8XJtOBdd
gO7dFEeVmuKjNnj8dwaofLH3MeMZPKZ56xH5ovY6UskZOjuHb2NaA44pu2dfZtk79tDPu8saHlE7
o+n+HJO2l35x95Kenwv5HXEbiVIuf1XpwtdGFAjce+xhTlvQcol8f1eSKYLoZDX75QVX08iLHlHo
Py4S3aE8m5OUH8/fWnerZXkGZpT6OXYpJXCaOr+LFjuwlAw73ciHoxPmGaX5I/Vwq++PJ9ZjPw4k
8VS2Ow0BVKSLVpWPeGg+D18zzqFix1hiMwVJkSkARsawQfLr4QzhkTXC4rOqbnshzI0kuKJMTosQ
GViBGHdjXCYLhjOtRSHrbIJkpR2ZTbjsl7d/GjgUpUjrFpe3lKsUr54FBFLJYo75w4X6r5S8sSNk
wLxGtDuGWWcSXTijOyqHcP0sL0ANl53xPhbfS7zyrAUm+LqsAtIATslx4gT+7i0DtgjuEaTH1yvH
PYHLToylaTydINjhDOBJCqNqcu+AKtiZfohN+Tn9MQnQhX7K3Hb7cAa5mHzlBjx5P2YtSyf0Hoi4
HMx4hZ2UXDZhW+Yv6nO60wUB4OpGRsYvZnz1oCE2hgmvQoJYPwgxBwARM9lotpmtDDE80G4Wn3bu
5P9ibcB9Vz4in1cJLeGK36PJJaAvcOQYbIo+JruyohlBHjABL8EUgJ4FG0KOLNeCu0XzdwPL13qK
hEfSl8eMWc0Yek3EdG2vxcLqsXDSAHNmIjJyq3GJqJH8f7bawjZgliHVqtvOzzxkl75YyvQgAMen
jD0V5Rxo25TmUVBVwQ7aYtgN10ksm/r9K9ZXz/f8VHbyIASS2p5btZ5nhkpLFKWvMZMQ/lBLKZTp
Bm0aMwLR5VWcQw6GVtJLij307eGC8b0RsXb7+EPW6tcmeb8KP4JVqGBMy+u18QtzrZx15dLG9oYP
X20cc7x3C3A99SNtNdoadnn6So442zkldxwfB7xx/p69AdO7zYmeGERYKAgxaFfhjHMyQv6ZGMOq
QS6ykWbBL4qD6t4yMboYis43gfNJMz9MlW5t30jsaJ2WEawUB1HVx/N1ecA3F4uxz9IgscvYlQlR
bnj9aY1RPBIuIEBOWN8UmBMfiwn988eILiyjVdw9L6DZZvWE43rbHNi+VzEcTL3Rn/5XdYzSTDqn
aksU/FjbIHEmLAXzQ0UFWdg51WdLJH2VwnCFiGj60jSn2kS9l9bIBhsY9opX1MxWocgbSNkPF2AZ
WtWZPoLIxWV3PKoZh7RlGfSWxdXNv+bJV98RyiT1VId+r4alS2VQtYrUL8414Hxpi+W+bXMm/95E
NGbcs9eF/UlCXj97dUfPgXg0OGCG5FHqbj0Kw9QbeiwZenLgXXnsyO4K5y4hPPc93YcXgGGWzOWo
Eg0hmITBDn5Eg0GanGWgizW+d2CczNTeC1NP9V/IY7V2Td46QEcF3wm2lsxwb7QlBWs0FIPj3mcp
ASLeHnNLBXD/yhi2SWJdMdszpT5qzzo0za8yxL2HY0CK2tGhXRzzJVz30seNgnonVe+ijxfvpvH6
O7SJxmy/4VNmmDxFN/8j6I18RSF9JN/QvS6/um6Wn9k1vZKR7h+L2rPqGa7atArbWFzOoMgdWfr9
pGQjoIlts8aIYEUMuS1NvzE6c6wy/O+VNjtbIQvPTiDJDkypcrHctREOtblELEJ3LjvEqOofYp/L
J/sPxLkOqDGH47xG57l6RVH1AtnAakUX/yLPhEfzLrGrOdy8eZ6UaJn6UocrdjliSHjbR8iMfyX1
sUvusltuxz0NVV098STthBUDUbbnfvDGf6lM+ZreSMkjvYcf0ZzNxWDdW2RT0CTJDTTiqjHZPZtW
vV48ogCDJ0fk9+v1Ta1s/4bN2XPlp2bWPoLHBSMnvlc5kSfaAWYgrv5LtvmAudj2MN3P4fC2/key
S2mztP8b4rsFdg4pjGVZ9dnJiqjUGdCT+mZ+CYrVg+6EzX9oEtAU39jmFklBG2LPpfIPIkEd0LxH
/KWY6mIaqD+DhRm6DhmdVvC9aT5rc8fA8XPHVkRdGXDdb8K+MP6YCmJzCOKfx/JkgplITx8ohRpJ
WyuJrCWP2u+8iwIB5uQtiek7Fepml4ReH8Sr/mEHdFISu2CG9h/vCc3SvXQo396Wmh1Dy9+wosIt
RpKtPm9mDv1OQk2EtHntsR7TJLQOCdXWqtylerqadMEwMiD4+vprEyz5f7dXa9v78Tte0UHEc6VI
xFMaljbp0Uigpq2YjxxIDR7dWln9fr6QuCYhQTfHAWH8R9+k7Wiht2qxmd1d4z6dZ/EA90ftXP3e
n323RdclHJS9a8GiPQdCUaj73BZ8puVjt1Lbtn5dMomdKGGNqzraoYJ/eVKqDOJYdC9g9PQWbUVt
Pn5DKepAx+QXcWUxON8AE6Kn2X7oqzysUTml/lPz1VJJrIRgw/ioIZgVBIemr9jsZccMb7x1IwLL
SKj1HgCrQIrAO9VahcJ7hTpYkMr5v61OLs7aeeO5vnDpJbsQsu138W7f70CRhtUsh0S2UiUTe3ow
XnqaYJpWExEpZFEDNRcJ5MKaNTXq5B7b9/f0oEMWllLCiA0208CEai0wzg2OG6Zi8gEtR309OAnH
5xf6/GrCKJCHk911hYG3cn0sjQLcVaI7pJmAr1fRxGrehNQJok5sDjRI46ZnhveaRtZEUwSzSMRM
9GiDdT6rbwqSnZo3gkm5AmFj7E2k3e4fxwRrNMWzTCOoFkXGg1bqOt5efY0gVtBUPK8pFCyeNRnr
5bPixGbVivSFfKjgjYLBqakNRkCo9wUg9uvUvLrewieeDI5pTn00sbjGFYgP4LKhGF25IMW2PVSC
2V29JmG8iKbitVfImlKC1PRNTfQNIacC8NyX2T6ybUAaFRfVTMXhQb+fLJh0fNX1lgcjeWeBg4uW
5epxCqxld4Cp7/4qDdmJ5DAXU9NfqqTb8UESv0W9HcH4HVGsSa+HNZFCc5eNejYQLlaBNQ2cNhpu
bhTPs3O0zhjpYVFN9DaDZ3G+bNWI7q3gMSoU5tr9umXvAUFEBKQ/C9wDJwblqlYuaWjkDgtriFja
yJ2mBOiYcp9wwp7OsxuE3GGzi6fXLflR36MB5aF4DVzUw5FegZ3uhpqxu2O0qTKALITQSF4Kz6ip
sxcxpioJmycN4wRFXbyVFsXG2NDAje2vrYx6GqMMRB00V3hU8X/96TKPafmnz2lhWStOCrkTzWZg
I58UOprC1TM7GfOlwDypvZzxroy2oHe1Q7yyb1WPt6foe0kGIXqZFmx9WhhfV460CAftuuN+lbUs
grRNCi9kaHH7anyukNAnIbUSMcqIQl4B9OmF5De8vn9BRR6wDSp/1ses010ATEsvvpu484AIEmgJ
+OpW0RHRCbcRgzBFOiulg2PFogI5PDc//357+d88IWtBChe4CeKQJgEzl9NrPXmjGS+jB+igsZSd
0VyXenyxtpcuIg2vfJ+DaCpm3CWoAYW68uGCaKqsLBuNqllwjUUwtjqw0u7l7w7+kweiFxFYue/L
VmhmTdG14xa5Jdors+Z1ZsonLWjXo4qH9uV2XjnbrLoMzWf0nHhPEa/aXJz/viXFV0OUmJQFGfb2
UKXVuCZRkXh2z7aeJyDzis2HFHfQmRH4HBxAB8H3pbXH29lQgTOQWJCpE99aWwvO/q2XPWdQgFmX
RVDzmSKSRpbTt/yo3me/xXsyqyWV2K/ADxMdyJz63yLgUTyZafLoE7kEAn7JBKleOSaF5S7AnsCk
iOIYNuV7b8dqpzvIaHHXSC6yVPBqueFt7IpoJYbMfuyzMlcC4UEyJoX9CBEUTg8lejDOr6wRrqpq
67Koeg89nCRlAvj4MgyuKDlnrYmPHbsgvXOmBkP+Gt9EU1x+5oN3pM5e83nFctlWEIw1Gfy6acZR
eGN/IQcrLECyjfAp/h+Xd0sUPcr1eKLhFgkqcSlmJ8DFp55TzZsR/AlBvcBU9apvMP/n40lKFJnc
nrfEJHGUm1mOmQt4LcsWA2C2z52n8ZF5AExuLsPBZRwqH0crKFOR7IFE4ya3p4xhyztO3VDXXfAu
asopw+WZ0ucAI4HMluTuDa/dnotCv5QFwh4l7Neghsl7LtBctYrhASOksK4yQ2FZHu6pAYRblHLN
6QcC8SEpGoVHnTETKfBYIs3zbjp0Evvzx5o1lRuqBVxMpv1BHbegRDf6uUYc+KQB3UH5SkJDAGYW
VYP6MFH9jfeiRNbo/jXlwPENlAfd92p7hNzSnqVOXElFaWsWaOUdtzRA+Z5bioBuHmL2vQnnytW2
oDzZYqP3eqrZ8cZoLTijqx2mq6fBEh55SA6zYk7MU165x3Yn1xdoIziICk1/uyUXPCUbHxkweCpH
rdwcOGSr8t/e0JBd5qxOT9ibzq1Sc0NuKrpOujLDdw8mFLRoe9K2vaJNroFfHMD+XJWG+f5pwl7u
l5W2XYMHj3daSCu6psRnGb+6IUZFhP4wP0E9j0cLY5P4RggUc3BIAmSWXAY6uigd7oQRD3CMOP43
wFUesVa9JOzJHfsh+GMjjvOT1REAshi0YrCdMKuF59+dyqzMDpg0yr9IACUuSCyWuH4JDuYVB33n
qE+uMn0FQqJqNreTwKIVyzl2Kd4tHx61MHgGbA9qxbOuy0K4xVF3VA5P94hmj0siOn9M9F/hI49k
+wWSlrI4R3wQWCeIv6onihZ2YM6/KthZtz8apP7l5Eoco8Ndxbf0uygJrhuoWnr3bXWWmk9yHErK
84mKaefcJR7tXGMcGxEHm04yCaVGpvmW+eO58kuqUFjOOWnX342JhG5uqlEJtWIU8IN7X1rXLcol
s7WPUfB4F1ySMMDaCL7IQ3DCl5HzL+vs+ikzbNcA4I9K/A6dh534cqIhIR64t3/Cse8OVE1FbPNB
Xa1cTCkRC6rhnCqenGGW4prrjZKD1hBvnfif0lOAOzZDCjCcN9jutcPTWuvEceNPuFAYIv+nVHLg
lRn1KbK8Ir3/OQIaB2OHDvhx6/ynvFURya+ffCspkD5RR/Lm2ohVMpCUwhamL6whiuLMoBlllzP9
pTkz9CVpQE39K9RBEl/skoagfK418udd39MgUTBEJuB+T5MHykLqxtJKYwFeYh+pnM8COnteYDCj
vLhs94I2DvNRiQ4vGTdmyg0lKn32eKd6C3y7mvdyCiHUiisGOnPQUVltYBTyVQwsEllDQUKPYXiX
LE6vLuxqRHGHk8y09iXOodzOZ5ZT3WDCo9D4rVKylq8uXL9jYN1jES5AMFIoWtP7cwgY4niuw5DK
uMfjNdsz8W4uaxthHoFe5K6V4lA0ThGXyPeMLVNQ3nHOiHQfhYguJyEGAuEKGzQ+lK+c/VxXIDh7
Q8by/NqyrdS7OHd9N+Y7gzCwRA8sfNR/XwqHqXuZhZKGBy7D47yOLvAfU4IxUK1oMiOqV49ARCpr
Rr9eup1voNr3CoExDWq5XjjAn6l2Bd3sGSWlwaRBWXPfH6Ao9VAlBySrbQKSnJZBHyDCSyOe6/N2
0oyWCDGbMEXfrDQuueKX9HxaRsLNObjHZ6V3BHMkexB66HgVlvIxfzt5aifn3TpJ4zA730Lue8Jf
vfEbty7A4abaVeTeY7sX/HbKnC1WwKh62B6yWoH+bWoXW3sVyPuCjQQWVOiLpnE16k47maQEUbr6
RXyiZvqeNBtmyuE7Pbb0y9hWwzKrcxuNtWLM0ah7ZSCTN/gOqwo1RpPDNsVoPHAyu9F1Y+4eABou
326gZXRWbOtlofSPybvPMSUMPmRQ0zqPn64bWsf4qUFT4GJGxxt9FPV8z1W1uRJGwDp35n7Q0CZn
DC9zCnPXJUqgTxjrJ4Ld/L/cJKPmeFr3zKXF/tAazGeUZ2nW7022syrQd3UL49epXInZI7b4Z3hF
4iuBk8vBIetbJEaxAZhPcYpIMVsiq8q9FZIhptCpWqiyeAg7kUhN5h6X/oMFr26Q0FrBLicer5+d
vMIf/xEMGR1RLfD5Fcf2hrpMcRs8NUEvi6N1g+vutX2jfHcL05ZOcrNXyzpA3gpvpsQqR9jWajaD
cLA1qCYTjVDU4ngh/jRVusVkl0vpbSE0Qcdt71b+vaI4x12KkBypfiN34MK7Zrl5atnFGTwlhM3h
pf5fQCs3j925TfPiVOYyNyhfgFv4eoBelztrO/KTHy7vLDGQKqgHdWRVl5qkP52a/SYOK/0yJ0Y3
jafLaNuaCnY4Tzd31FMz0f2favI7ZPs2nBMiiXFhntcWC77A30bgTRBxCZd/vTm2ZHcmEW1XRpAR
TgW3GDkWp/VjGNng6syvA2E39Zg0778Bvkuju63XH2PRg1qKJ4WnUsvSkJ1qO+IWYhxX5KBFuwBJ
MUT+RtKRNg/dlw1SDQ/Ac7p6RIyXGztiJEjNwNF3HhOM1C2LiCUgm3Mh9YJRPmF5mX0Snc5wnFlV
TAnkpzN0/tKwRRxeNf8SadMaHEpYh+cNcLjKrRYVQwcFBjOHAewpxDWOXsMZuj10iij6bbdwDR3O
AVrk4U4ap18XiRAfBMTDghhviPEnHjyGIbKinG6TmmUGjEGIn/fve/Rb+mstFzXHZ6V0Ni+EleNE
eDe+cPhwQsSLm2g2nzN+IJhCEan/lNBk6rzSWJl9jRVwXVlmUGIdnfC0P3S0JZA6Qfz7SfwLr8j/
r94uh3PAdCctDbl2JgC/YUS0nwZYdGVwuWBBOt6D18k38dkQRQn7+E0YNZa5VOTH4/X/UlsBYGPE
J7zSNqRtwYg7MBFTUDq3KoSZ76XcATZlX4FKQHeGnYlyiAKmDFngkNIVCODJ1RwXdGejV33eI5tZ
BNxX7ZNVlAlaCUkWBzHg+I/RuqsOq5KCuOpel7xcq/tJrE12aKXlVzMn7DnEHk7ebLsgQdXx4pIo
XhL22Sshu+CMuFiHRwnl47xCk9ec/TPyJBsl7U0b3YBXvCH/MEt7W7yk+k3wWNlXiH5o7/bGdSD1
ZQrJpwmD0EBfoz7EBkvSXdGbGAqKCPAgZyepj/KNq7RJ6l9W6Lqg+E+K11W4sn8MNGYEAckUz912
TVr++S+pJa/AGWTKz6tMpDvvrfGF3YcdVdaHBy8aYY6KaZXVlj+9Y1+/d65D/Hc5iA2QZSwhyIOm
goOVgtU6d8NyFeHWJHSHtnHPgh+VbBDjo1WYVfBHuq82pggBQVrdpYDGzUfbRLPT2F5gsm0jkAuH
ThsmXHm9Q98sHft102lUZWBenBpMhKVGxsFzACCS/Q18kWjef91ktetJUVcpvYxBj1ampcCSGKIh
HJ1M6q8yZ8Ohm9WITRjMq4Gf2KSV6IOp763gPidiESx5kh+dix6tPWZZWudxNEj3D7V+6jDFk3rM
RtDfMQe1feFrlDsopLRkuwkSIm4NZIt/v+SCeQy6JWHFAEYxU5XRgrcA8wfa3HsngpuMDsYozmfS
f+6MMkDkb5NDih4CJ9oc88NUmb4wf9Q/9eyntOnEodYkrAJEqArZ/VnPDlDvDz3G3iWRLrpnnPbx
9ZviTix7PQ1mJ5EIcWIY8Vu6DITzs+1is2GKemMjy0BR/DS63c/VMKlmVTbWvNTgwuWe2yzwSNIc
RIAZL9QFt4s3CqdANuoMJA2rxZsY1XyScY3mALAiNJinqGgvMEItvr/Z5i8SqQE54B21408bOemQ
IV3jDQNO+QELWw4l4QvDRBIl7MHm9iVntq52QVjL9ND7MEHGLWq4WmpDjnH2Ec0Yty9isfcSAB5p
roZNNgIb4NyU5tqwbuH93BY96/yGwZDvRREyciJZTRCWBHdnlkvNeketSd4jZwYf/+hjpC/etofe
24XRxqY3X4M99J7g/6boQk1BLz4MtSH2+XaAu1Gxnik7BXKcNHDfmB6eHpuh/WOIHovwlqY/B/4w
LlYVJBC8QGA6CZl2IUZX8HFN3PrpiITl5+x5joVl+Sx60SoxXlwZQlWkWy9vCZVdOHIpf1giBoPJ
u56vz/xrrgR0f4Evdw/RnLGL7dX3/zngPMQM5+c9E6uzDOvRIoh1RirnYwpj9WlYKeg63Eda9leD
UWb2MVc/bwAeQXmLzwoiqoARF4oopAncAeNmrDPlEiXm+8lwBfiMnDCapdchO7XvOW1ADiIAfY47
ySArqGcp1Etjhy8UFWvYD1HVfE7b7mWaVhHQvc7Hwhn150vsTziulSleXBbXLxOm7/+B+V9RjECU
IdYqqxMkxIH8AxaFcOshdfEF3s5t+XE+ixU5lPtXPYGDONBVpadjGHzLjoOYv88SRWNBIzMsH83q
46e4YK44N8YzTYwva+USJMB8+yO8KYNq0DEKxzC9cW+BEVjgmgnYql4ahYWnXUiTiZAehnqkwQKF
TEp2XwiprlSMJ2uu1RhDc7E7wPEF+kxsi+VuRYkov/dYoa/uTdyn8spBDMGEeB+y8fIyhCGJjOZ1
s59musLZ0LDaVZP6zFGrgvvlYS+fXRWFP2S3QgD17GQ5l301sLGw22I4xB6gSoZpH582euet40YK
Veue/S1iihJR2LCNjAYwGOPuzf+vgyKQ1VdmuQBc6OnFWptuECMIUlZG8qCEhhEf2Kd/UHPL0Be1
74wtye67uSGRG/gfIG2jm5Mz36SsrI4ndXbOQ4yl5wrctQEdHRIuaSUb1hJlnkGYZnSuVLmh7DWN
giQaljO2atgBPDRSb9SG+a//h2btDX2Tl7PuancH9iJeUTIowqCUeasXPXyqdMXzCdBWamgPeyKy
t2m/xmWqKHGQDJIhoxmLZovboZXvN8IEjli7DKJzkVfQjkEvxEEMvNsymRy7o5aP29wZ894Qe5+w
np3s6vK9r2NSiyGDa0anM1N/QCzPOQBQ7svhhfBV6uO/Z9XPhW0E9XGrJ/LZbea2Oi5N7CYDXRC4
/UU/sgVdOqGtoJa/Ft/9aF5qvojLWSj8yY2ezG9o77I13MrV/65pnz10d72So+/Ft70zqxDw5hrv
JKHzeaGR5EWbYCA3PXgvQdtemfA6fb708V85+PNExrKrT2xj1oINl8gScCIMvnS6H1YPu4/m7OK4
mL/Kwh2Q/xKRLJpM6Ga9DckWutVXf3h4ZIv0ROxHsVuXRJ2B5wzePz+iNGZ7zmwEEA339D3b4E9G
RDEDWTxEegaAKU09xNSOEhEuX/ubOYbWB9Z5lPp2OGz0PXsbxqEREv8/r1MsYdXF6GrloDRpNVFY
x19zr4g0BmDDJFrNU3CiMon+wsaqZgHrQUKqitUFg5vi3fwgd1K4NJxS9TzZBm6yw50c+f+p0nd0
FzGvSbT5i1EKy6JjfQi45PU8u/Nfgx/Giq5eoA3YzJX4WupHy9hOn+ySXVmhb1h161y2ObBfwlqy
+mUB/Inyu2iPbZOML6ntrYUzQTvDk3lBBtghHVVPvB8laJidh8o8oV51JxKf8HLBTBP2iiCx5KyB
9Odk3qWPOlp1CrOm+V4fBW8yly4zFvArd+k97/240h03Pe77g+O4iCZyFpt0kuT6l2k2tnx+Drpg
z5+2oo66qJfUknz/W9QhJoFNKtPTisrZkDsVd6q0WNOOfZaFlpy0cjA1Tv9zzZTAZrRrQomj2a6g
KNGsC7NjDviJM4ngyXdBCcMmAwXn30FW7vABB+cHjHRoxw1wx0ROqAtPj5+IaEbGqupewG5DblZe
pASh3qJSFtLYMNR3KxOf4pn5mL2mM+Lb7TJ9bz3/tNZv4oORLqIpZwZI6Qdpj1IdAdW/oAMdBRI6
mbUlwNBEqxoqbDA0HmLchn6jZAQR5XsGk6PTOMYr/et32gBVmdCa+CtycAge4neO3tJsgpfbmW0x
PWLNfMSMQKaBbidQz7SOkqWBaBCtrMXLrwsDSKaPRX/hTHILueWJFhgnNrXpbpNWXOPOgQ6G6vH/
QLEDQSxmOYeMvsA1HqoDiA5Hg9FzggJb0+dG7Lepp6o25BnVjsDQ7KLfI2rd6i2VzeRLySfXs91B
5mBS9HhxNm00KM5TxAscYbZ7h1dySClAIk6buJ6TDuDm9fyGkaaOSozebFZAhAB9SfmBz0e6FPGn
ylz8jXEvGUgEoZODF2SFeh2W8JcwKxb9nx/LtB5dShQzirYyELiBdf/rVSRh4YkYZJArAamH6dJZ
ri7i2+vWk2/awhsKlNXATX9gZDSXEZUM5Fm8lA9rISdYb3ZldKeJMz6wg9xTtzbZUL5uZnTkfJxP
lRsKEy6wtvTuqrV1QiE85veHBrf/Gm3Kq2O2u1Si2PO6O3YOJ5yG+LalyUaduvE5XyMqKkpQ2MOT
j2N81GpXZ8knmxr5TD46wO5k5IjvNJPc1+RPuB4z+siMYmvf/fajfvirlIzFYqPc2mpSZhEuNcCL
Q5TE9/N5bQURVD3WrV6akbS0ZaGkjaZ929mb2STvfGrTI3MriW32w3Fnt241ct3dW6BLd8hWG3Y/
68feO9jjbL+81ZY7VBFMxTuFASAbxkAJhEH5K39THslHxB+qKm/lKssZWmWpnyjGLJck/JSunY7s
WRncdsZgOnNj3PmFoDGvolHwSA+EDx36d2ZnAnEO9lMtzj2DT0taz5CJQPEmYII+bOM6/j2HOQ3F
bHmOxz/9SsEzmPgByCJlp+8Bo+K2MqgtWghMTyDq76WwebT+/JojW4BXCnQN1An8fMc+TefISofg
vrWv3NycWgfrOOZYJPokNmWRfQ6mCXArTrGlcGmCTyIhlH6mlmhjDogxS/Y9ASPn7yJyNt0ReEJa
rokxLrZqJSn0Krk/39Z/A82xQg68uL0PqiD8ZzT+viXYmHKNrEyJ9MoPxhHzclKurLPXa4sFvUp9
TEVVaRHijH3qNDdfbPduFt5sqz8vRrkcs3+bqfsQ/q1OqHlALo5X/pz12UqMMGFJQdko4Svs2x9J
HipIM+YyIw3xPPJv5v/estR/9x2b4U/Hy8/LXnnpAPIgUNPdR0o1Ed8CNZUhUgrhX5H9w+9/xbQp
g5u+t8M1s0JSg4xZnvZ4q+kK89J0reXpnYiI9BtWYyOxHbRtcIHfMn797MwMHOt+QXoL451E6yhC
t5DqyKMMJiyYEpl3Qu/4uWX1VOzjpCpMQHMZQrBIQo5sg7hLhoztVWa/13Tw0m+L1Bwk1lGXQ/Fh
hz1lSVe1XKHeRrIj1mRc6u836oxsK8/L2OFtoGotHNW3gEUijoHJsAdtW0Fp00fPSfWCDOQhxXdw
qbE4YiV6EpmdWbKX7+jZMkxdHoPwOwc6v/5bDFZOXyrt0IbCS3KcjlUSj/gmgBF967AEkCmwzfGQ
VSGPKdbuqjEjvCzxIwav3UkKGy5c9sUs1qg1QVf9zUgaqCne11IKKRDjEKeYxMiYGTVb+530IztO
oi+1eT0sqHGRjnenqghMxCWmJjZ+mkHJGDfSr7Nx+d//hoXbfopkCl14pWnQTioNEHcs6PCHLecu
yHlI5UC6ec0x2U0Fnjryu75AHvoeqTBZ97dGLfwrvX8Afe1yyrSruFUaUyJKSRNrvGQU/f84DOhh
zRJH4XFsiQ5mGjEXvOw4kAGhbIKQGSxZSdtwynv2l+e6yzQPCTfMb4HITiCKXoa8QR90vcOw+CCg
2NIh7aD7jzJ1PZtJ2anTYdCyVqD14B++CvYUyTuUDMXnBRhsHE/S6x+oIGon5WCLs4dJSxYz6JQN
h3IidZNXhB66jOcNyMYHc7rIj9wQuap8W7nzZCOJdH4O9HA71WPObtT8xkI4bnUkyKR+4QFfWpDA
DqqSt4XXd0yC8hIeCDTEsVamMJADxGYHabss2MgPZxvxqY12vFB26z2rF+oHoJo8beiw2l7pKJZK
WRNcoVuv5Iz8QMmuYphAT7fxJYBbSDLfEULYXvsHOPD4GH/P6EEcElumLj6GQXtIlr135iuTLiIw
k2fA2Xu4APenOTsD/mH7kKKJszUDQdXQjGdUyPKpbW5tdOaMcgJJ7zbbq4WW7O6mlA7lH2VJgh/x
YDfMFVpJpc+vY08TKD+/D5mhU+Nd20g14O9o1o3RDJZMD6ZuxR1yCVzADtLXJ8giVF73fgjGP5tp
xI7pwC7P75s8OdXAUAvhkEvUCOGF3bTnp3ZlP34fbTuTWxktL9C/itplHbngZj95eZBj7NS+U9lj
MGQQEoYtNqgX/QTVwBoF8c+T14WT7aSQOzDXwAiriTMIFEhaw+zJ5uH8iAVq3RP3oIWyIbL0TwYT
4lEVC9RXf4dupAI63HFosz8BJq69ITqJnbH8vuNOqpo9FOimxdT3gGZAQz24JcuEOgo/BbQn9aN+
maGZ9XwwJR398Yv85IW8UHevUh/sa4UqKvkOdRCRA1evW36b1UBUH8w80cwMpSiFonfaNN1J8ST9
LySbQFO3iAGwOyWd10U7pnU+UDFm2u3j4IxouQDcTe0TU7XS81lxV1zd0hnuG3Y6rIgP5QEarOit
4+c8d5F0CDf3PRfRnE5dBcIgZEBkBtqb3MY6kWgH6/haTt9yYeTSrVXWCcPZfPktpASr9UE/2kx7
Hh0usw3Hed7exWb3pdzjU7mbehYbCz5hOHf0v94ky5WEVgl079TzYPMWeVmFdLcj8XHYz/xyJIAt
7i9Vni3aHwGh2AoGCf/ewG6qW/YiGyw0u8JERZFvvdlGehup7ygSw+dyp2Nh62KddaC7157awP6Y
ZbTE6c1E1fkPIfwBvv1+pp02aI8R2wPJi9vbwUzp6edb/jsTb7xtHCc+KJpWaCLxdyWn07JS3ujN
BbO6LjAv4Fr8dPSzAwkKMSEAHcXgufKrnjtxmcFKj33FpEncvy5ycb5q/IpCtuMAgx3d7jSnhdKF
vf0qeBOetIk9d7+PH5rbiH8KP3xrh1T624udNfm0JJ720Vflc3pJChzuYiKqDrP2dyVIRjGOLkh/
98A6SvtdxAdDsCEIE3MAZZWSnndedIV0UdJO5PD/YAgolTjkbQ3mZciVFFj6L7jvFLByF+3IRAxR
xhN1cx2QT/tg23ZI8ZSg2DipICuAqewqoaBuFhG4Q601oNzKrssYWSeEf3iThVTvloI6d5mt/YEd
AdXS/9M2yoxHfynLIVO8JtwoH4C3tGNHO2tYIMW32hK42tt6IsZieslwCLUuYsD5zBWOI7CRkwLS
OKlhYZFC0VQK9j8aKGAswb2OkCocizXokf7GxtxZyxM9/0UoeunZUciC1juMZ4x/6GJhMWp3Zf+F
+JuYYq0u27NQQlptkoNgsbK7/H2P9NbcOM2E8GDSv+zEGBQCb7P+IQY10m92BB5TIb1cnWzHVNac
spoBkuBFofluroaR8nzWEYQWS60qA8SIXptKu8kD9dEJsjUOC8pRfAxymD86iCuqBVkG9yUUW6dA
W/Dzno33rHoblmmj8EX5IHMRV351+JWnsgOHBE9XRLMAsp0kYUCKDgXgzmiwzjBaGeoRk9HkVA8v
XANtAgncztwpoSLoJ9E4Fiwb44x11ojtTE5t3Mc3dglxumGmRF3fIPI+GI7JwSliykEgwRrnZJrN
ANixKxvOk/BcN9tzr0kaMDfgcJNZVR92JQU+XGZRptuQxb3tLapE9APfugqt0VTGyh/+9+l5VxAE
WPOKv0qVxCDpNytxHeprUQhnoeJKFp7SAgjUvOalcpsxSq+4w9NOUUka7y7KX5iB56ML/tV2k8kx
SKpCQI51WHv45yqyYrHZu+udrD9W0/n41AvwTIQuMWcEGzWTxP5xef/N32Ul83mbPuGsmtxkeRYG
T+uTqfiqYdDP9gVBfpDteRrCigcBLgEQaT3uZUJlr59/n5fIR+wgNiXPBdywTbcVnzXCzyx6IPth
160QmUWdkgAAeIizYdAahZRZH0gg0MaTg7krPwpXJC2gfiRWHQ7tavrAvzPegUJoTFNqwdmwzjfh
4LO07XihJK4EgENeeiSceL/ERYJMF9epUMybQ9BNffsCUoRKf5EOj6PCxmEvcEhg+E9pUaahx/Fe
tDW0wSAEJUTP1gIuEoVH9kWKKm2VJHXJSVI/HmJTqrK2uHE6lcoOtXeO+QmdMyYB0E7mvjVisofz
c9/soqMlIkZgGUo2g/YaTsWsS+d2jnBxESdK0w14PN5VDRC1YaxuED9ONK+YGbzwIqYr4WdbEUBn
27IXBMBl32AAn72kG90Vxj6+60I8s4zt2HoqsJz6gYjCaZVdSEFJkvf/uZ/S8KnuoC8Uq4dxa06Z
Vx7b+NCMS4mC+xyNBhBXimBVJHiP98jIwYFH+fGlWZwxumxFOLcLQTalB4su7JAp1V2TVcjkCAWI
oFiXCZ6NHUCDUPzkKAiKjH8BVI9vrqYP/Pg/poqCzOo5gmZMQ7gETDrGTe9sxmveUMjTvxwUJaP9
7+ldBMzD+woW3vx6b7HdQSkDzvtxmFXUztPFlPQYOVaym2bh9Bb4qDhCKeGcgcdu+XFaIab/tbXV
tp+68CDQ+loOvQHlSHs3HOsWqI0nMklzZr/tQfXTm99lleua/A62s8VtQZSLiZ+X9SVjdXVLQh8Z
0LmDh6bijMjm/WotRfvIql2OsM9SwKS8yMTyU4C+5OT98DqVrCFh0OlHYFauiSHiD9YyOqz8/NwQ
vgUPxJaU6g8SL6ptoyCo+608rIu1btE6Zm9vm3sA4eKLEB/27+2mN2B/OxE51dlxr4hVKYceeoAc
NYgZbHZBsOTApSi6J6SGWITRFYdLM0AAyP4Vv6lKjqtds5CQytC2rzaJ2GRLOPQsZKMNcDampZDF
Gk9yIU/IEj1ykgY59BAIHBajggvqBRP5eoAG8nVGjTtfrSSB0ZcAGiyWT3N3/D0lrPDkXtLFKURb
x4iOrFTIQ1v3PBsDX80ARnIGemmW83dIiRcFLUp7omZprwcTKInNMs6pdfmDYvf+lDuDhj1C09DF
/AS//UMLLAqSFJ8MMLRmQUH3R5L6duPX74OVq152Rk0U2jckg4i9Ekoo0lbf2qh1Sj6ECGXXNnTg
t0nWdZj9OB0PtjSEQcEXZ+Qq3dvSc/EjNiBmRVww+C8J2rKhGxpkbpI2NjyHIZK+/OckuIsg7k1h
XLgriS+MpBWxEnmQwltCwM1ztvJBNTCwdC20EEl9M/2mKpA8nMIPOIGYcvEMQjWHkIUQNTWrnOqi
BYkEsBGqC8QxlcrPYA703dwaAbC7DTIkqyxtRQvevjeU6rzWsISxILVbNWaFsS5Ho8NmQIZNX0rT
dVtbkW4lt1GAZraiBYXkFDiBTYzeGdONGmobUxsw4TNyW1YDpFdjJMCslJ98R5RzXDC5XxUD5F/Y
gcGg42rD73Kuch6fjtHYYvYJr0ymON9RyhUvWC++K8119jtohca8824VHj39iD/BAV/4jDvHlbw8
M2doWYl5Kkf/HCA+1lJ9ryDhcBbo/3GrSlME4LGyBwVZATbjXtEPUhmcV5xYF7e8FIyGzaPo+XL7
8Ay8qst/kPk3+TbHqR9LKJSMaU9k5qIk8d78XfSAI+HdVgjVzMvC6V6PKGbKR8wVejqYMP52rsOw
iFrdSjy7aauwfnpkVUGvbRYBhFMFh19A2adgAeOm3nA/oPtv2+jqehftl2Ec6Of6fEZ2pRJZj9se
+S28feJZ9ST17hTjxptB7cimfCv95rb55Dey8wYx4/l44q6sse9VGxvlQsRG4QaH3bsbXO1QruC7
IdBGIc+VAWKM1NriqsU8lrSvClkHpIrtoxIo6C6BQ3nJa6YrhOpUF9KZBu62f2dFOKn39EsqRLSq
BFISFPIVSF5Qu+9riCnuIL4AwmNL0DWYFSsHYQFr3Z1aJruSaNnaavFSsOX9MI1NaEWqhgUqRIa2
aHAkRqaBnV7D96l3kpuf3jg7WAHYprSbRMSIUH0IQOuZyNrLwxx7q/F/5aSAYCk1G2P6TqWqKlRj
8tqJK/pxbhXsUmslIYrtCshdcJNHGXEROS/SQp+b5oN8FTc46WbhWs5kdNJhD8hV1FPv/mzO4dk7
KU/t1Eh92Ekcjrta/GYEjj66o+UePdjL1Q5RkhcFVp+eX6dOzGY+KY7B6b6u+hXyn9HM/cTkmIzM
W7t+/sci1Z9ub+teBtuf6EmANR9mPukJoKphBFii36hYNmIv/WqJvNTkQBNvxAVvsiyPyu2g/7+m
vy3h4+jKJmvgpt2VwuAOaaX26+3ALmau7KXPUJxf1Y4Gnpu8reKBmgB5DM5swCThFcjcD79oh5n4
e5QfmeV1oX75qKoLR4ce65pfPr76kDmyvo5OcZqNu6qOzyhNiZWh9bsHu9tlhWqJWauOuWPNTKkd
0tHHYyav/PMsENjh949EE9+a+tmMjw54gtnTMY5pWuxTqKK+t6vzNX+mGBIRxYGs+sMXfn3yvb/5
ii+MW0k48H1vK1TypMtUFb9q9eJ3e9O35EaI+Wxmb1n1sau25PiG9Csp7pzXwILKF67ha5bfm6z0
QKTr1VS1+OB9u+Vgfnn1MKPRR+WzJzx4ztuS3CmfYJiZgPNf/IQcmYkKdTx+7AowFzOB7Ez/PxFV
J70RjOfNn4OfDLI27ypGqzOKvyZtfaWIdBUO7gOC0nAlElxiebgIW5b99Q1K+ZsMz9u0BiNQrD9V
KmOXtBDRPUSLbPcqk+sK/lH/+OGAz2tHDeNDPHx0dCfB9iRe7I4z9C190fyX8TV6bX7DWLQEF3fL
VxMkeo3wVoLEFcm/b8OGibQOqi5UzSkPNhoCdCminW6dBAXRMjGOOIQwwi63+UETiQFqmXjoY8sQ
P+ab/WI0ZdNY7Gze9+GyzeU6GG1Ak8eNxuagNPQ0Q4rPykQftMiw9iI4VQ3eCRvQIGenXEpEutRw
bS21UE5TkH8WATLWIG1yIV7YNv0Nn/bpYWv11PCoUj3lXOwFnjN+zPQ8pgN5PLJ+OX3aNysGtrH+
TaZvQOtUXwbIOgEgiJnb8WBfg3G2VytZ+7LZ6/cOAWQvtuveuHAqslwfS7pk516FvE9euSm4kDbX
k6Q29KjseLPzJoV5nxNFOOpW5us8CiNGbmAn4hAT93YtuRTCfvDgpluMSxKhVPcT+TMSHu/Wt9ri
okZr6InfAc/dp41C8cMd9oII+bthU8k5BnQZv5gEKpn2tGEJMHkdCHoNH+s4NuiHeHvc84uVhlIC
/1l/Ni4uGdBFIlXhuC697Q4CRT6PJcV5JLUrXwobXCEgz4NSUX8PyI1Ogj7+MQMaWzFw8XG+lj6N
x3bxzQ5JOusCMuqvnrBxlsYznOWj9HZsBsooxNchCsLLW2UAqlvCff6Vp7h7qAONSjW6P+c4cmb7
JPDPjJw7tWGznk39v/xACiKPdBKIfUYblK+rOfIJ1ErlIfQbSbzn127hG4QuZIQcSi4xj4z5JM7E
ss/9Gsf+Vlf8+tHmu++ZlAUYmnXtEtflmS1/49TpXM/XG/kAypFhT3JpnE8oMbwYTvYuXo2OsTer
R+PHE5Ca/LZfpieiTdSXiemyXasUPVzjp9/o0jb72cOgAMv8uR0nFfsrdZpJu3n8RfYJ9Q8t03/E
1VS11lo5CxmDfXnv0MoH3tTjFFuaLC3lz9cQ5Clj0UIilPkhFoxGq9GsZmrF6mDjLvgeEVTaZqZX
znFsTab45V+HUbM3NzS3nGxH7LW3CzKCS/WFd7myZZD5UDOZGMmeFgn7z41vC0UZnAwma3HP6b9h
gikaGWRqe1zmGnRLbUe86Ydkkw7Zv9gl3IMSU0+1m8zvz1FIKVwGguKrL2WucjIAxaFuSZVcqkNz
8wA1JFDqXkTVTNDldtOtz7uSiasSyjaFK5XdEXNJX7Yj5bro0DdtkCfrwvfq/QSKU1NvTLI0ZAOX
LOqW91vQaUzu7mU8x0nFzRJ/IL5wyMLxmbKoLpVu8iM42603zSS1C4UJRgML1ojfzr+pwKT6vgli
13bNnUl65MoDRaXvAceOICSvsriiiqZKkBw4tQkd66lAHX0pYmBmwQzWxOAUjQygw2mKYSQ9gY1L
Cu7+16T/8orrjsmlBR+nmeyiIJPiPyuJvs++6RIKS2q8Rcbk2PFLdNng9R0UsY1bjWFZ0f0YVzfX
ygY8X3o4suHs3GowcJF1eoFuF3VKIUbUxK00gK+KHP+CLj/e2zjVAgG+PTBzb6CbQnqHHlbe8S3o
4lFFu6Nxtgd+Zx2upzQ/uoX92QL//+ZhGKn7moumRguzGgNp1r7Ara0fKZ/086EIi1wZEvF8GqE1
m8o21j//CuVoQB24Qf8V1DTb2sLPFaXQsRowfLKJjb4irlbfv1hxdPkNvKkzSH1u/H6w2LtPMhn2
+5CXYtnu9JEM9WvLqrj1T3QTl+RCsEGDJDCdnlXE18nPI/JDZUnK1uvqkfc/CKDg1A1Ds1Uf4+s9
wG2Nr1bW2i1c9VfSApYQAkbl/tQ7tCEBRvFiZ7mCc6twHTnDqod1PQgFpFgwGoWbCE2iq+xx/tCi
+1Pxn0A6H/B3Ga5fPBKGCHyl3NGKyYvmf0r97zFqHfH5lSoDOJGjfXP3HqdpWtO7HJDFuQRKY+G5
gvoVcqUmdoxbHtiXNQfIg2cDHgR5ai43jNZfJ7Pw0ioOsivRMMFzbiPpFr437QynbqHQpkLP3jF5
Q1JUvMHev7iuiXtJvgRbz/qPaRSrrqLU4WRxzfvvDQyWQ73iBVdl3sE+dywVaubY9T6IJsWEuoys
3ShpWVNrEd17g/XKoUZb2jw8wXKwomn2vcY3EM5A5HWVbNurGl7SUwnnDE43kowSAh847D0G3OSb
z0Jie4grb9BSOH2+4MUEmDrg2Z/xfR3fqlJnQmaog+1gJMjP6ZJO1FkhlxM9wgd4Rl1sz37f0xSc
LD/xIdaCNE8PTPNdEal2yN03dCUVA5strRxIe4zADQg1jrKTLlhGCHBt+u41/uv5+3g7Af/ILbU5
WGsvxMuK1oQHtNDKs8Y4bqapQIcpeqlwzWY+edk4Qp+pc8IEKfd7LK45BwQoEChdym72/d+y7A8D
VAI/fg1BhWyu2N9JzAtNnVA9KE24k1obAuGCsiABY5S+iveOS2sLXFisfg69+cw3xXiXtd5ZBJRN
r/DZIAG9A4Qe6426UFgI3OQa+XMo3fdqNdM/TUfUAIKjF6f4Ve/hGBrgLzDQ37eOPiXJ0AZA3ueh
SPL0hG2/38lzDaYjGqgF78Gy5ta05Oygs/DXvo/NMunPs8LzOyMVxmvrFE8kdJ5jMsmTzeIbfE1q
JkAcD6jVue20TX9gJpdOFXMHpFf2wYpf57oUT2GNT3anXmkWGKd690wJ26CGoveqXn7ixNaLCYls
voYul9K3rfECWhwjokKUxF1FkldCmEBdTVin8SmW2s0q06W44H3mJ2FRwwaOJhlsgorPY5fpR7jW
GFmZ7Athqv+UUQFM1Qru+pHPqciSNmKk4KXm8Rkh0t+HRyOChFLw77CFwxmXzeKPkRKVtEf+/VUh
FNTnN06iLRYtHAnfkXmZX1wGXCQg3t0qGE2/+QhNhM78G/KYr/3DwxmmIHo7B1/xUWOZzbcQL3hO
AeMfWsebcBZI/nQCaDxC1rcnRvb428fVBMd7hmUMr/u9pGIXVGQgyDmJJwHAZPv5XtwAVaQfrGUw
MfuCz3DbDKByvZMeMu+BdrKCa6lh7od4kWEh0+Aq2gASlgHU9xjDUhyaFbsem1VG5uACjWSFGxtg
UrW+CI1+ybjGoa8jO0ou4IDtmjYWqgvrkP9C4uMGcvi60vC8SLeyjcv9eEhJ/KfUs6Q4JihN4498
6+/ek/Jen4r/zvbFWQYpQDdw9Ed2Z8k/WcTIyak2iVCxar4iKF8RIyHOgRhHKn+DfbKpZYHWhEVU
vsmt8ZNdmC5zCNQHSWgUzQuPK40sKyt4J735nEeoPmqtDaEtruTpmYxIgwO1rlsahuVG5oUZLn6d
1FTt/4kMAhXSWUy2WlJNXYiUZt3mT5XLwTpjl//SyuzpBrBeP+D8Dyd0dJVu0Fdp9YagF3Whnmoi
D8h0qGskVI7f3oI83P9cz+4HBT/+L9kO+XCEYVfCARMr68LS2nnrE3MzrrdwVwXR4GUvv+3JTOvU
fj4+jk4qJFufSgAgKg/ZgGJXncVZ63ortHHfjNXnqxcTk8YPRo5SycYJIo9hszH1JzQnUy5GRgxp
Y2O3XtT79dR7Q1POhXi1IlW/uOkoLIcLu+hrtbrMd8P9OB8vO04C6baTy4VpnLuVjq2cL7443Zyy
5qlu+UmYSxNOZmrz3gG6fNA5Uhyn3X8aEw655dBZx+SUQSNaH7LArTcz2jBnmi1TSMZ24JPkhvu3
sPSp+8rkD/P39k1p+krnvsSQhYP1S+M33du7Yg6hWHxdWHToOIiO55cOMjAgPhn955O0muC7Gx88
MR4Y4/YTNx74ib0L8VhYYhQquHdS7AC8oPf+loorPt5CYXjNYE9FgDC4GAP25+M5CxvvTO3vl9a2
h0Hxhwn/9qPqWc8l6sTnQAhb45on3pf9uuR+22xJGTDQQDDdHp1OKC2+yQdp4dJIqvY8SPzCVZ7L
6DR6KkP9rAfm9iHoTGqBb9FPl9YejkUkAIAfhB0pvsdbW/ncKzh7bXCvs49HhP0UOQQjxasx9ac1
7t5A5DhegiAMPoGfc4ZXGmmiHd6QCxPMh4xT0hatkndZW/ONF5Lu4BSq3jtPpN0GQl1Dv3zPP8/D
9mRwBLsmFDx68srO6+2UOll/7mF0isE48eWrD9rB2+LonD3ZOkYF9BYXbCbusbxPykAriRw6BE21
3h4Ua1ojT7bMANxMMolc6goYiqPOk4O+6DLS3dj7iklK+JmR0QW2Mih/8U3JztLzpnbFCS9YPXIC
+cM5KTLSfU59U0GtAROaNsIiAsPthlCc1KD73a/RgE1C5jDx5ErX9dBxJpjjRf8VHpnLJNDrMnib
qQQrkngdTa0tLkGaR/239BQZ8b+KgclnksVHXSIQ6ASY/MPIM2mlHWkX7atDAClHAkxYOsGDcRDD
+rATozfOb0rwsugscCmkp93UozVKhhxqGxWtDxLSHfqI7aw2qUyz7KoCWTWAsQ4enDP6z2m7mUqp
RUGSKPSJ0P3qIKk8HM7ulVCPhoeclJV4883GrM8hUaBnkPK1EaVzrXT+ioU6ik5QMC8Y1PPhGA4I
Wxi6hJeiMs65PDVGpQ5aODFlsrmDRnmSRJQsWGObR2ArATbMQEAwehIyEmnGB5r5DpIse966MKVB
RV3zTgCnzb33FAY/dLynzoqgCPp1Siein6tkojy4LyteVDSoji1RLnuqXuNAu56gwwAcNapiwQvq
ZMlkmyO6x7KaHKcBc9MCksekXodxTRDWF2P4oJ58RmbjqF3de9/zKanj0/Q59t4Ujj3ysu7yYPrZ
qcbm7voqZoLTGOPuUZFTSQ8YdrDfi9SdCfipv0o/3vhpQuWX4m1y/aaF4odXYDrasTiu/ejjUaiz
SR+ljspRHKt/Dyp/cNIH0WvruQUv5nEAIv2bdWGSz6E8+bM8BwTXBwyXqCdFJW2pbFvPXE/WGv8C
ST+PWDbXeqPMVpKw2MU7YPXHjeofMdzFyGi0NzW6O0wZRAKa2aNa79Z68uw0GYhpeJeK/890LRNg
uSQyPzigaryc7GZvUh6CNi/k7jViufyvlK/4LP7NRJCZS+5WDsq4iMdmTSyiHF1uiwEgE4M1qJLO
fVMYTSy6TGFIKxPvlxYDFiIs4Zpl6PE5Y/Yi4FEM1ZmMenvOb9wdL1s64cOe8bnDbSgQSM8uxX76
hVv7e5UbdbCePzuN3mFmFJ9fxWxJww+FgmmMgB0OsQnh8dOSVtgXSyZdOxcu6aSmxIDgpn9DbP5/
BWJes2x0KlM+smigE/fS+twsrFF3hIPNF/pk+sjrH7jIspoWBpuMoJV6U7App6qZx1ZQBhr6Ich0
zqMR8YWWlalLNPYXSzuzxM4z9oAjmDNX8tiMMh2EFsC24RvxVieL1tAyHwJakHTiFPviMN01/X78
rBpYOR0nVy53luofxJuLE4f1QAtrLbRe1eO4/UK9f0uJtg5DCSBuX3wGH0USuvijXH3hf4hsxmZ9
FIZ0xXBDTqW4QtzlYSY9pIjPiu22ICEyF7l6vPiETAAEoXYByECdrsMz2NC2wEOaaulL+S4Iy9g+
KPAM/o96110F4ZVhNy4Oe87MsVQCLWe7haS1Am/0Z3LEN2nAE5Z+swlfdfpPixDAqbK5CwtZmjwn
iP18Usq6mpomKa5ZW4AXbU1JWoY/gYHXZLb2PzROIpwBdoUSdq60rcHHFHZOe7e7mkhjftfFhBvG
34BE6URfgxcfvrGU0C+G5grSinPJoxWo3SI7RcsGS87d/ovz81/iOxqWADROBuX2H/Vtc3686BmA
th04jcAf1gNNK596RsgpgmOKiRj12398nM8Sw47kl1RY/AxCkkkzk/lgJgysCK4GSOjyH2cmX1p/
fNgUyxkZkbNOSaXUXeCe1HOzcKg3Lj1n1IQ/JTCV0ayZAsN8CKTqsnCa9vOzJUGL8Ezv/YgjzNso
0DSmtu56q9X5kp9L0nIn/7yEUQu5oNdE2FR3EOoBGcjW0SEEWqB0PBv9Z5PCGpnMxP0HitZ25VMM
6IsgOjEzruOl/gD1JwVUfrDMuoSE57LrrmBK5UmlXIpfsyn28VeCzeN/rQMs/WcrilnTsT/j2+Om
rfV42/o5uyFjGs87XW1WtOIBB6LuVLdEw6sbwhBpy2S2wmiUovGcNWFHrvg7nAIUUkt5cJm2HNVN
I8yVjFjHDnF3/b/mbCamNYjbXUKldGtgkt78R3E4FGxez+Q7pFqO81lTdW+/Yupem2tuAMj5xBYH
PveG2yXqwU6bgctmt7qaDGFo2RbKRnZjGcNUXRJBiEmj9jwQcpamhMkuJ80VbxbBw3CjSuF38t+p
+N4JdBx4g4eoM00156OdL69jcDDthGF3okL72IJ8NeXifDBdpbZuAosXAMdRCPPMKzhn7gFdUGzM
HIGmIeO3XYj0ib/lvqZ7mzVZeuZB96SO4rY7K05gQDKYn4o5k/qoAUHW2JVI8x9I6BgKkXxZz1aY
/sm1GmAXaShll+6+DsT4+vbJ1KnnoBZml9gRinbFnAxN7zZOidOws5ZB6FR6gyegQaI0G/qTtYKv
vGpeeRTA/tlfWoJX/cU5b0GhZYMC1BaZLoNRaVhx82w0uh8RM8lF4bpp74lbR80xwi73EgLNJqp2
I2heTMtRfyNzgkEGj/uRHHWTN7M72SlEVIZSS+ZHWSx2pcrTpiERRCZyo90DzNVtbUGX9Ga/ASaQ
UGCmUJIB1mbdOSuEvDDSHHpaenNWadus1eo46IbY2hQKdtBon5MxZQElB3N+becNPb8yt22icXHV
uUCmePY+MI8y4ze+6q98m43CamA4vHaX33e1b4lwZHsISk3Wru2OGl97KBxiDx6JPb6ES1DZO3B7
Znccpg6kO3HDEEJqXLMWL0USXZvBxa1Jh6+W18vvoap2740NgqnPhJqLjpI+KLYgepR9fW+tojts
Ovxpy50chNHEiKEU5yMRxOD1AjoXqGEasrvJ1vGYQgLtVzc2v5N33z1et5jMz4vIqvYv8/oVfqAF
ULn3OjnCwnO1KJpck2CQudJG7oGQPeG0cAkXVwEonOusEHF8YPU8mOPXjQXYsbjxAeWuLwB6t9YQ
+ZrMMXbBPYIUYxWHn/uqAt92OCBhSnMkFCJ4witn2GNFNsrK3e4rRzZDOqoR2FBNg9UMPJA/Li9Y
jE71NXv2ql4Wtd+BzyDh4QiJRcwhb6iLuQCd4TnAi7HbVbgn87XrmhZDa2dSjFQyWDvfaba+TXyr
HFTMpPzsLVCnoiuE4Ro9fLC/AGkI0q/FH3da8jquaLQc7VLnT0PigqzrVu4KiLayH3mr5eZKtk6C
uKskGGDTOx+C1/pTheYZHEb0b48bUG+2thzoNhJjHSTLB6T04LzD4gsnpDJAYq1+7pX/yWADcSdy
8MzS0LGo00dn7tD6zEtTTajWYl11FirnkQHsQTQ7jG+Xf8betHmU3z3ZshmWXZ7kTlxiQJeEfgOx
ZN0zitE/kfWi0L9CbID3Xpdfzcvnq77gngbqScWvieRBZufmKSo5FZ7OUWubVpL5QicgkhwYgz1p
Zjr/uLKFT831sFlMxDFd+BFIeAKwfdf6z2stYBsS/3MRoTU8VRqWCerkbrd7GQ65piZT3xC2/mkP
QAWOgipPF7QwWvoBLW4pncXecyXjd3tNjOWtnoc8CSlXFSJMfMFr7FtWQo6gU77FsZ/dO02cpe8h
XQbwCsONQPVBCMb1vYv3z+st5BzCv1rzpkw6b9uJAomEL+dZy7fs08i+zOj5WMbUuw49ZlXT41r+
2YmEYiEbDxyhIOd/gRfxwvfKpl0ujjFni+kHxTWk2k4SoHepRVw0kV2htn13ZqxY4BxYzP3RykWt
VKMZ1kzAtaBJgoHFU5aVcA0u2ZcKnUiPJreHMu30cJ/gJm8IpNcoeHWAJym6QXMqLqJNkcBxm/u8
hkXFkhC80mJhZdpRCqaKXxM/P3LIDObQLQx/SEWVdeODT8y2CgsRY0KyBBApvATOeAlsatPeqZJj
26ow1ahJOvfdX84kVQogvr/+ipDzz7bIvdXbuh1L9Pp0YaPEkU5JTZTRQDPViU2oaivCHCm/rMoa
t9+eNRMEDSmoPjU10SRZS8e7svur4eUWkboRuAnKmRyZMxHy6LVz852N2dqf7WDvug5yJv0Hbn2y
ua+Cg9V4fwjv/XMfAXjbiiHwoC89/luesULkiix2yqhMyZvTUUsXOQ0DxbOKdDB3EcPpMnMyyZCm
8NDnsN2eCvk955ZNHvhNKFwoDMdH8iC/amSmbUuPPGXV5Pd4jJMZsfUQidO046+r6bDBuqih1mzD
E5uu/518TFTTarHLQkEJW/C0nFOuhFITt4uwC63M3/td2Drq1JjNV3oBkqxQMnHbz2XbqsUnshlM
pN15P0yLLhvs7a6XoZt22f5NTg+ldjmEfbEPS6v36HSMa9A6CDwWeVpvh7LwMU5oV5mySAqYvxdw
vZCHIpmbfCMclWP51mnvLCIrrbGFBXEnUFDYcnTOW2rDNpQaSxiIJFCWGS2KKpMffI5ukIIbz8Pk
VFLw/F+cgPpUh/lqo/OLF1gkUeGgeK/Sb2LBCrKFb49juqk004cO0Q5BG5rqmZeaazsUHStH6aj7
0qGsF8S2uj7AJrdvhjW+mrolAV2+GfufZs03/E0x3XrDG2L3O2lr4QjxIt/2l/pQtBqttrpICUDu
HXMHBsU3SQAiUEyf/q0TVhn+v/Dk0P5PqMxJe2DnSv3EtdqtdbENmFnfVD/d6IO7eS9sqwhzPR5/
pq5SPH+K4WyVFoR9NNsGwPGXbUvjV6+uUPZdcvQ/LIBW1ti9K2N5zD8yb2N/DX2K6rmLTUjit3y/
en5GbIwR4sDaIUaY2DvyiP+C4l2p+R88ntS9yneLINtq6Ej3489AsFU6dB/N2N17szpuo5r6nMXL
3mcRQH5b2JBnqqInefeWuRW6tRTOKjxEPgnRtGfsk5yXH+ShVkBjumg3GNqrgQuaOpHN3uDnxFao
eETugXgsKM4tXb4E2urEid09wOw9CXDqmR1A299W6fZ+ltBC/iAU/KC4ByFgrDbEU0RQWj1lTsrH
3u7dWa1FEjOKjmCujLDOpnrrES6iB1t9y9YPJf1FX+v2U0WxP3VWuuRZQA7bE9k/lOdlWzNdCCND
Ksm0HWgHLFo4m3lGUQyy4weJzWV9P8VJTJBRwoQJnsoqA3mFulDh/jMnHnZcLFfb1m6lJkOtLUEL
f4TCJXNHzqmO4h3UHVM+fd+FIuMjYb/Zq0x5f2ewZsiadBtmd1Bb/ywlhYtjFfz5htsilZ1U4W8t
os5KUhT1V/bJmXmEmgmoCpZKnDZca57P8kserrjaByDw+ZHwmvu7Yj8UjJfZsg4gTdYhX2ZFtsb1
38u0kuniGUNwVyT7AvHHVy7D5jBkM80hrb0A75HzSdyn0rA6axMn5IEI9gQzQNQ3LLWCICMKOnjP
goEPBt567BseILI+wk6bNgdJmJeRFp2ul/dbl2b/4P9giTSCuUZL1dmsFLVtlPhBIOdUNGJ5lyho
j4LLowQvrmP9gft4gr1OY173rn4V+prHTC445myJvmbds7urHprQOKTV6+g6nKiFPi+WRp80aTS8
P0kulJM3V1txE9I5tA2h8ss70MHkthyoVJ/Tkp4M3/l4mLbjzGWVz/bo5dlBQMPb3OPCCNegX9fh
SUu9PEL+9SakOle7hysMEfKAS0da32OKs5XGDZHGmCHofUru1UVT9rCgLpdyFNOuReRGE+p3NwCu
uaVdmLpYhhl7o7SNzjx9KJA+0fxcesVSxtPw+G6D0FjgwAVkvE0sjPgHnAdKxrkd6Ty2GU55+Cge
oNZb0boOsdBB6EZplLMTT1iBhref6WjTkms7ECDphnd9laaRACgjgQuV/f9fWeBl8YiE9JrUihnD
lY/18apfn+Qtp/8S+JzyO0l9NySCWIDGm9iIKqBkHR4KsDGwfIGvfbaKsX1jIvq06AbKHkwdfvaj
TkkZ0/S4NQrphcl7eoC81NiJSjhacqTER7UjyZaTIL58FNrYH/143poTxxwo7b3U0FqlCqc48m5M
HeHVOz34Ajpi648fzj+6bXMUWTFOgOqehMoogtVygHhC4hlajzxAyBW62QU1TxBVf1QJKtJDRWl/
qfTIzlXOiYGcl81GgqQTkoUrm3R+hJLe5y1anRSbS12zzHYxmoJzDG+26sNgmsjFspBfZ4PoHY/c
XQJKnKD2saipC/jMFRov3MIZzNGjrQjAjIFUs48eO0dgRXMygQFkEcDLDnxMFzq1iIhbP+X3ZAwl
9CeNxekdrm5+5qkhpna7sl1c4vbUWdMD+l+F+9IAbqe6A9aGqVuTVfarC4sgg9bIU1O0k1Q+nyz/
EP2YsfZkkYMshmT4GgK5WzlP5OHkGuniEJqlNnrS4+xmgP2NlBWvkkS2KYArgMWTkN5hevo05eaP
iutmsKEhe156WmoWRzdYxx9G6TSJawCI7ffKvusGh+e/+BESrJPjR1qu95f5BWA25vIYKZsdy9Wn
wpWpjAH6qtyltB8MarFaVd6sNxZk1UaLZLz1U0uTCdBJEcViFbUl6wg2ci6G+6fRLEKUPMX//YXf
+LXOYPujfJcyRpv3+a6/GAA0PyfUkMgnYfRGPl9aISBunVmElvzrC2MBQTqdgPwdPDra6D/eTQmy
EE6Vk/XxrqvB8Op6u+5maQnOhnRnFJof/1zLQJ1DadoeiZUHvp19np9FeBhfGCWxLpEVdWaX70gM
W12Z6st4EbV6EUwEAuqUsqbiAkiTwQ7iPkJaYaHm8CFINB/AWLxcEGMJINLT35ACeLk91/8t8U6z
GKFSC09+u0iTKSsdfAVmkRy4H+htF+SUjTilOMJw/Vj+BZkmNxdb4ZhgxD7/fG4bBkfMCWyJ26UL
k1z0D+260w32nvzhkLt/O+wu22304Q/8auOpWEuyB0Xr/lZAJxAjysHSUXBt8Q8JplsX5cl9lIJo
Z84RvMV/piN7IZLqtm7bpdaKq3xsVWZ+OxubWlbUcyZAxEaKOMXHByQYccDa64kIQ16EIEgkY1FC
KHHmn/gL+YzEScm/rcIhjc1UQh0/vmOQlsWbu3+vEqP7HgyjMSI5zuegB97x9dE1WoD9pA7V1F3a
fFAlTNiPVnRwkgakKABbmKJy9EvAbfmd9IvGLYk8fcOxZ1yz+4hO6fdWQ33ZsUlqhaNQuisROvw+
ynkbBzH1UqKvGDBNvemP6yfx2tXLQinmnZU0qF4Aq64lgAqaOkLmqD7PsYx2vSHQAXm9ZkaT4Kow
2WTqrcUlB/qc7Ev8ded0xu27dF6NBr/q0WsWR2/zGTtfzZsnG/hORn4aA5dfoPuAhRi06EGMMhIs
C0jNteq3WZOl/2WRiHxq0A7sAHYZUK9cHQhzP3G6AGv7IL8xjftFwq/5oH/Ca3K13DH/iHwuPkqS
Khwe1kE1pcf2gkuex47MzT4AanXrwsZsKoXEVh+c98s8Aq75xylsH89TrF01C42N7sGt2SdWXivB
w6ple0c4lwL7JIlXK8YrPtGVcco8h8rgUTb/HZt6nw2VDmWPbe65DjK07zjUQ4aOQ/rcmDORcXmg
1fLyObjzdbbnShUW/p0Xlzz4aRm5jzf+nN0lj6GWkQoLS6hcnfOx8utC8iFoerU2jLDZktfrkHB6
BSxifpKPnXcoE8R1VHFzA2AWDCehHSuGWPJALh8Irh4QXr67l0ZNkbF+qZGgkp4bGcpzKEXP+/3K
bx473r1L4w1eOFtiQGke6tamgEobc1b9+HxJmt7ZbLDVWn/7Kz7HrRrcXD/yybaaKmPK1XK7VKhr
2ssei0vFQKH5tdl2FBqG/qAjTxhQamv11sORCtwRh6Wdc4vtuU8WjGi0X7psX9sHpcH0/sK2XAn+
V2mJnk8newB/aS2qGszrt/6bXhugUjpcgLV9oFmDAl+LzqFmz9YYNsbwUbc6MORTMqC6n0o+eE4o
Rjqtoi0AcNsG5tZokpYdTkrqFR/3nQtb/DjRMz5SHkxneiFjCLNk/oqyVOkVXBePo1la5Go3byQf
Vqda++3tL+5bTWU2lUiU8/CrQlAIhlnZDxGgeyUrJ4UNu4WgTSdw5LOt7ABFXZWRMFuok2UrXjQJ
Mv9DBBr/G93PqDWg5M9pEtYjgNDbZJCSVZppzMuQ5j9nPmRnPGpBhgCEtrgjgJKHdJ87CfeooVEM
yUbpDm/5EkdQIO9gsjGXtj361lczSqCsT7VkwTOqFO9AWmfF0cqY8yUJhC8sBSYhl5My+9b8TAVl
PEOMRipWwO46YFfhIVqNYOdCIz2zmF9ZpejGRjNYRuHgc/T0CxhjhbglfQvmXvQxQiH4mUNnyddn
4bkoJivkdxGRyk9ag+oFWgToE9FjovjfIuVTWyYs9MUy93tYWFVwCwF6uvN9QUpGJ+89VjOQs/G8
7kxTqlS/R9kEPYlZPjzQi7CNQBnUEyi3kI+Hz93BItP0eZkU/xJ8xIV7+jxJ3ui+zysUBvgG2iFF
79Y+8IRxgUinsexwp69nUCEqQjmzDrmlcfgJ4VF2BfVbMmIkq7Y0HL+UicUh5jgOto/XUtv4nYTd
un7NW2fPLTT/pV/8jYBULd30o2N8i+T5gCrxnx9A9m5UB6LRqS79Yzh693JiYvoylTVBIVN/j2yH
/k/g0OGxZWbIgtNZK73+R9s/ua+naoLMnIsSL460Mim24vbXEILXq+Keqo96nfELXv1zckabT5ED
CquNkmTazfU4PIyJDeU3cKsUE+BwuL3++WPwvvV3LIXt9+jozTnJQRgL1fI89eyn6d1Uxf6yDoI5
FuQ8fJnaVVMQicxVYqaChiztHrW4E+NdozV5S7t1uO1y75UFzACplviTod0DAl6TXYToG8p5Kddh
UEWWYnbnV3mBI3b64tUHr1C3vm8HxK7bMG5EGxohkHeLfEE893n/rw0YPTAb0H+vigzuyAStubVp
u6E2vxSmhIeq2URhC45E3GYiadREuSKpG3H5S+f0icRVIDbXs0xu2sPkjylRof+YVilDjtUBs2c8
mluWk0IAw48tjNM0EpvSgGl7wNX1hkfoIMqBlGYtUbXB5S8ZF7/YdmKcQX53NRFVdnR/1JaSizGK
mnMZyCtQP0paxK7XHusGyp0yZYgYeC5VbBnjqDSLaJ0FztcDbSjGXho+Zka8CN/sjNVAVAjzT1bN
WvYQNZzITytAVMhvs3sA6HHLC+cWOmFUAI/nkVvzpEtGb16adkvtmnboj4VXioZ8344YVoUv7XTH
sdbKlfh6myJQn8mMtoU9MZ5xBy7TCHRDDgbmi1xFIqq4P+SaAL6sweDs4Kr80lrp8Ga8VK27A1/4
0FLg0gOd3rEkf3flwil0ClkT0Up0mAAHmXpd7xcLdJ3OwfBR1NFH5yhXdJodQolLdaDRslXMun6I
qBVN4Rn2IZe9y8n/g7MBXNzgKYeoiCTdxsfAkwbo6ucXIXZfr3G7YMrH3+R5RJ4MpcL2OEqJZhF1
VgoQFStkkdcLRwVt1tyYP9C8DuKS1F4ZMzg4UdKZQwTadr+McoVdGLgVIPomRYZ2u5GDuamLTAjo
amxWOUx16hgfjgdtlKVrdGRwP5im4HqUrQW6yH/uymUTO5kJHPSZRAU532KXXISUE0KEeBF+XcLt
yURMVl/Fn5tqfLre4kCrTmciNacbwYphTn6QhHQoiOjVelImohH7OXaVr5RU6XtiZ8yPH0hqU/wN
xGfsG0a98UuQpPQ1wJsT/4qAEEaxB8HmUzISTUBCe181XRDhA4lsIvLWbmtViTiKsobIEA9Byn6D
j7o9/9vCWID516ENzj6uBuXRgPYpnvkwwcMSds/M6Y0CZRgDghDx85TXWanqGMFYljpxFHKBuwA9
V+4oKel4iFk8/ooZI8g+5c9sV305LKr1E6LZ71o03f+MSCke1V1d2buuc2ziac9GNFJEKmTqJJw7
hIYMaUa1SyfHEAxMTxAyZscyuGAy4S36kaZqJLSQ2an9nUPY+vmGLbjmcBTHZxkeJzXPuMUU6C2F
IpiBDbz4nAXdlvPZLnkZ4o9445Y4g6fo2gftJfxjFItBm9Je6ZK7IT6BKoGDfZHFw4aUpplvDIjB
aM51vuug8OicrSxAdTMZ5mnE7lSvIqqW1L//quleEKvB7bZn00/9fQLfchFrJc4iij2aQHedDR/7
HC6A0/sYSSXN07rGgllHwfF9gDV/y/uVIjwAWDQA/KIanO0etJaEJ0S5dbyV+NAGamLCe+P3wX4k
+OYXOuKfQ7jKn0o1B50iykxU8rmNlXxnjlh/A94XoldyqftM8E6NxSKm95yUji7y0CrPudx5ei6r
UvtMLlPHArZFHO1S7ECseB3kx37udt0TBKkqmr22NDKXUz5gKkesQgW4eyOs91zz3i/FTrNA1OZ2
Ger1PhTPIpSI2KWkchclZ4DvR87rvTLA6I8GeUucT5IYukZ9p8eV0M6csQVj6jcLwY8QVklkOsUS
hbC5VJBbrXsr+w634wR0GNZ/9K4C8taSPRKrdKfEYo+4I7ikXc90zgqOeFWTpv1hKlpWtLLfnlPP
Cyj9xanNKGro1mLk7aE1UnhZLluvTzq8SgI4MYRAg+6dvO+9nW0t+/lwl3r11/7L3wz1cIUnROWP
DkQiN8/9dc7bGSFohGrLVdS5yaTAVkDJjPllk9gD+rwoKFqKyDqV2osgJHGciQTvDYTxBxYvnwcE
VMtI7EPxNrEIV+nRdjU3bQI0soZm8eKVOePdXahnEFQF2+p6mwJEs+TiVrEVCw6YrWuI4enBhxP1
qbNj1Spmvu12s+ruXmySniMcCxKM+An1cL5H+gZPM5yKHXDzWC4kyUWcQoC8aOJLrjhwk8orUWTO
vzUOCdqeS1JhDpcDIAevo2QCwn4XFL8r/6iiySw+1WafJaeLlB+ZNY3+ShDyMjLdXx32vcfjEgt7
Jl9AhnuahOLRd3bCXXB6Qpc42dSsFwGCYE9cI260K5M7rVTtB2fx3DhjhfJPV4mVbka7Kv0msJai
hgF21N/lDPwqcubHxwXd+/GFxb+YkuMeFB2TC0oIjc9bIHIOXRVTShe+IoZTJPIbgOXzvK7Z5rXj
GJxMVWnFCKqOsqneHbQjqhoBqL4nDQrN9avGcMAbrVz1iiYsBwZvVzbMPEcNNZI8O7D4XCJEz16K
zpDd6z8erUkofPZaxOIkGWsJ+2L3tNCJPzV2zBeHQ3qbQ+wdux9CHJBFZECiuiK0pIeAg7HLg4zo
eYjliGwBH2PWSX5agXwjbvBOgwhSQyKJwn3EHf6sDZ+RdlVIVopVntB21z9etLy1Gb/QiTVyPNKW
FYBR+Nb6hQ95U44gIYEeqIbw4R2HiyJtSdzOZZY75fVwzLwPeUVMgvHTOV64KKh2mD/FT9C7KKIg
+atkBjiziYuNwvSbumF+oCy49cNcU6mmg+L3+hevI1uatQF/a6UCvV+bP9Jr6vWiCuuknCPr8pqQ
YqQhzkD19pG8o0A1u8ztqt38ebXX6ZqnXqKEE/VIspRtNTI/3XwC+k3o1aDNK1mlXE7n27ghiqp7
wMTsyeBzX7CdUaeSLbr7CNplyGzCRWVEFVhuaUo+DE8bkt2dT7O81ihgzR1KOR/3yJuIequxkrWX
2PTH06ZGUrJV8tayGcAqu/ksfBGjJ/CCq7hDJBzpr/peg2WEM037K243N1nJbANBMDhwAiCdg+G3
srMvA0+7B7i1XAobOQ/33WjnWhI8wRzRE04WR1UNtzRSG3SusOBlsPsxMRLsb5fw9UNq7mw7A3R/
ZmP10R5JR8+AaDqZEx13+aELZvdZUjJqpFTuAC14FDNMGGsKH1Aj8jqZJPAgnvFHwXgXpbfKZHD2
LAGSHMyhi6jrQs1SmJ1p9zUjZMQfV4A3UZoN6QFRUPyx5zf80cVTF+jYqqOQGBGPRdUymn6upAW4
1UWUh9f3HsgZsJU/maUCqi2jGVbzHOMCwlE1WAL9Up/lnUBs6npLq8TLtDBmcwfyOmwsjS8dDdRJ
dy2uOI9yp4WzbhhdrREj5yGhizBOLJaHGLkntwFOvJTG1xU/c4e5OHeaf4qX5LTKyTR6QWE9TpJv
em54vfEwAfsBsPhWiFA+YAe5u0agOryguxOa+xGrYc1IYQ2RGnXue8q5r6UbPrnfmS/NTLyQUO2N
kB4Y11U0KOywQYe5hdkIO5kjwZwFx97pWiyUAmZEQjsIXts+igqzSHmnYCBl7Ynx56r6pScpr8+z
eQKl/x2EzQljaYvnpxOOYczpvzk2co3tU3Rudxkb2cl3xMUjAcl2oCSbrNH2AVhNix0cjiH6jbPi
1HtQYhGP5l/lmFzaOzXNrtbQfQN2wdBn4C+qhfk5oimvmT4hDq7vfYN3pGKID/Wa+QuWtbMkZvg3
dBNfaI9eXYSqiD1vmVxfbYdKR8lhhS/JEuOS4kSkINj/nBQwm58mEkYp6kKPqbxTltoc16DhVTfK
5180pB2L3srSF7geC95u74EUcR8Cf0o4mdRTBHPkaX+8aqjlC2y5H5T5/x0UD+TA6Y1R7m4MhZv5
nOvNzlZ5CtHsP4lvdTmQPm1N/+nUWY+V7zvRYX/C+HDTkJn34vGNymTI7IJEnynVvqAjcBkYHRNH
5tWXBTXxbBJP4KqowcVE0F4z9Zm70PMNiAd0u9sZWFwrq9Y1d90jpBnS0zj72SVLSQq8FAxZjuFT
GH0dQFxryTaWuAyFWn7tJQ6xtyUaYN1sr46HErVtRWOo6beJjt9NKV9lIq5j7rX/6ewxauozHes4
OPbJTxjAkXHp137ABHf7w60LnJKeDe2Iq0OZWymtPfjThclDnchrlbtj3VAZI30tMqfnmufh4rr/
04CyvwfiT0oZJROsKMC+mQWEBkOB7RvABuk3ycq9mXo4AuWui4yeUbkiD1YA5tlpg0SAtmF2mD9p
lgmreJBfdtYPb/Mg9Bt2d+aJcCi/25KE8uMdTGeEvQteLwY+9igl06DjALkvWG0TftB0LJ1ygNp+
ioOdbLeqSXOdSog9ySjbzZ941oPNfWDinxUHp8c/4aqxtZPAXObphwbgxywhBQKtn1x1DvDXUuGh
nfT/Le7J6mGnEv+kxwohGJfkWyrSZQQUVmA+K/wXM6UlZugQXy7yqtwx16oqVimqmYVUYTNSTO8o
3JvgTlz9jRrRtx8VGMEgsGBaD6ipXGY6eKYfiPkUWeJU8vDtYKq24W3/qqdhp9AsSWC6OfrTTAiu
XbYKLcvnZaRCKWKI6xEA01H3IerIZuVlSJmVdYKtTafPNvDSHIVwYSXAKuHyjvoi1lvpzbmhGeMM
i5Bld4GaJimv/w0v/7FYr9E6u/AZpOe4050w8fJew/rV/ylA+h0SFPrJCU52lKI5xj+JEfGQNBug
uAC1Ben9ow1yQkmyC9YbplM4m6DSk4p4rIuSTlJ3+B26B15Axoa5NOB89+edbyxlJE8Ljk0P7bGm
feJxRR3aIXQb6DwuZ7Hv72n0opLPxc/XdwSltcIRLPQtv4SvVQJkTCEY1uRaJbyhsShu9xaNMa54
j9RmLejfendBn9M8pSNHv+PMXMIejHcWNxVUuMfhLWKmA6veiK2mZu2flkovJJIy4JU7OQiooDAb
uq5k3U0W5J8/LB0j1yBPSaftXg8nx062T3++X0wpnzpr4m7ppd0RVbNopWE0lmlrGbXGCfWZoOXE
zkb5i6xZ/ThQTBO/flaVVTCsQtiIAbV3n8FOG5HBOmbrJpjXstqZu6mpzI/X6Z18WlbZkOGsADr6
7Cn+0Mla8lNeo9vdJ13FY6dNNYlNpmr5BZO2xCgGwg381nltGPVWMhTI6qs9GKr5W0TUckZwocUG
74HtU1mKGcIz5AQy4VBdikaRyrnoqprYhHHrixwTnx/LU43kKXt2L2gPB40ZTWIcVpO/3VzRHQSA
H0EtBv5pSzvbbrHrJZhKB4K5iFo1GIQvYruCAbJcwQDXAnObBmR+9OdZQuxMj2rZnzI1vkupwRyX
hAzF9nTQwJ1JKp4J1WtDs2V+Pr6HsDuW2TrpGDAvZjHwkYPLRWnWlH8SxLTiRqU4AQAaOb8UlB7i
C/Wsbcts8oNOFXyzkXkSmMuhY93jNurLVAVx9GyOw9Rf0roFUG6UIHi2RUy6aXTsT3OhzohriTuD
KcvvcKtTT6BZZK8KUODfGhJC6iN6neWmWb+to3FVOt41FvD7MMjDek1byDoHvp93pDoBZeTY3a2t
o/K9sgDKg7y9lfdLZ0IFcLnG81r1oUr3ne0+OZMs8yOwrgvzoP0JPd0Jy6qtv8/B+sh7xzI7lpcR
8jE4EwsIwI4IUuEOjt2ORjiXr8CA2cogD1iqrsFi32l4XG+KATFOqr9VoY3PMl6hCESPX8e8dPGF
uZyjXiWWBEE49SjCXtq/zFiiIqmSNCEBe+SoQ1UATzc1RpBjew2sdHNjmzzeZmd5hUE40eH3byac
5HYf7P9F9uA9nI+aSXf1UcLaAFYgZO4DRIRlaXOBI0z+UQzJXDQAHl7CWVJD5eXZVOvxYPPBDywg
7UXUDnRjp7oNwYIP7PaB0XN5WqNIwBVSa+VRupbixRT/d3plU9jRcc+BYcRwjLGu6V07RAmx2YbG
fRXJ2VESqUwz3pT3pmh6nCPZpy/LweiRSkXIBE+XOUGQbgRVtQiBJSOOFx2Aluhvd3238lON+3gc
sGwG92FPdBpmOI1I0pJNtgMnrz7RePD2Lav5N68XvCU7ivAy6j7lDLwyQ1ecAjawiYAkr+CyOEqA
w6TcA+0sMRYni7a8xkC1aY5ldztEbjK+8mX0G5LMbEgdq/dJJFfdZSNKoGFJfR2QwbjbKDSECwsE
S/KhNd2iLfqjoBpNQTzgaWVdPywcDrm+VUuXiLuIODyhpLvmE0UPaZPMhPmhIkWMBpcsZ9iXEH3w
Xkwh2UMwMocNgxZ7ZZ3oTC12ykjVZDUWZP+jofn4gzK051A4YY8VHb9EK3wqdfsnKUTvpexa1NCE
4P1XShi9rusM/R3Dyd3eoXzv2QLcgeLRrGpeqR2UAT/UCMXeOPOGmzII2akGN7RaKfqrHh9BUduh
r6+VGvb3ibPKpPvg7BjkLp5wBq7/ElW/3kFOXiIZuyd9IWluPsqKUme5jHz0BRpcQPXMLpnMgoe/
jf1y378rUJL6eeFLd4aTi1cxzEtTSIwJWkTHrzPQmavK9TE9/YM9rwMEJRdvBt3dfTXBfsLvUkFQ
94x48o30UzuN+sel3jflCnQER/c9+7Fp9ywlgEdLhibmNgW591k6S3lDZtN5eaH2kglbmRV+qDlb
NZ7ZAbRHgwd7YhpycUDEu4avKLq/axCvd0E0DRXW6GAUbj8GRu+4Jp0XV99fZr3z8PRhpL51WmVv
CY9yYlc5AlkJy1tkrBKz9jy/bchTmWv+stDoal+pdbwUrNb5NEmvPKoPclxk3MuIFrpD9zghuoTu
WzusrLWk5fo6lv9Ns1X54L3U9760AksQjusalmDphzQlDGbKHVBRS7sjqm0DFfhlpAW3/H9dJudS
+hR4ATugwohJWKZDtyi558hW4hzsIRksSMiM5x46wu1lUW5bvqmmUkml/jku2tRfsKH6iHwnTt8G
Wic3i2G+H3Qr5bjmNVAYPPr5mk1co4//p8WJidWPFbox0watq++SR6++uhR71p8NeR1RHP2j4ARs
BbUqbcRu01+Y3nX/8zu5zbtFX3aPMRkjiDtSNTUbI6UmVWG5np9hsxbDvNDFNxs0j0y9zvsvfgdq
VJYaTxLRFAVTM9idog6kc3PNmpQtzAd+c3wzPA4wPCqc89TMbbUZHSB4EgTPqmDwrZ77Fq6Q5Opb
OKsnSltyzJut+r/LQnwmd6QpKbXRwwteDV9UnXdyqRbF15M8w3SEX5zSzN7EgJsEbK9E9JUywjPm
i3gCb9xU4PhxU6gYBZjHWBgjNR3QAvJa4kpjtXnJN6HnevJsDX0Vk4LkzH2MbkhxCgFb4/iWx2fK
KK1S6bG1f/MpF5K/go5I17mpJAoJ5nGTXLXr0v6zfIggoWl2WsmyFRyNgcJxuZJYqoIY6nd8WUgS
tuALdN4KP1Dq8pLqaTtnmJSTMSiH3E4Rn5pxwcXdPqTz0pmW3EC5JF79Y/JO27FZfTqiW4r5bp+S
wMR/fFNaSVgGNg5Pj7fzgw8tqqwJEl336tckbxRn/JRp7ca2kUL9+I3XC5xSWS98bnx89sTxvrNg
NjLH3lZtGBjd+zE4ig0UHl4Zqw1HrDDw27WDm5ZaANu2JY9y15c9lqn8TPCpBD3W01bNvBE6eVu0
bCdJJAdPBh6r6ILhQxIrdT6RFJC/4vGrslAMaix00LsMYnaijISUhcWSV1CMHsjrvBNVw43Alwsa
imyu7Ncw05KAYq4CX1u4ZR88d48vpYM63YGTeYDKtlc0G1fPbYNuuqF1P3RiMFXtytgyBBXZVK4Y
jSiifBW8atLLmaOsAHgWZ2kqxoCMWUBbJy5ZCa3b4pVJlGWlJ4hZ2hSmiOXMI1HhlgKkleSSqjsn
EZOweJ7ENvSf23UOx3URneVyRBUPlC66Of6rdRRYPVQYe389oH3Uwx1akvtZQFFGh2VAbSe3PIUI
SNxKJ57pLtVfKMxK48LPWT0N232zXCJhnI40PL2x7jCG1+3T3GGQCcCqohCDR61YGqPCjzJ3DPOI
C36wsspO5AJrIbKq4yAz0OrQAYQH/zqux2u+PdSF5rRe7GvXYStkpw84dOvSNRXuzndjHK7QMP61
8/dMDTKR+PKcVMwgL0UXWge4H2H34ve93dNqabp12r7SQUn2BLPpChpDsmh0Hj80NRb3vM8D8GzO
tG9EuZv5lhrW+7C7bRG/1bu3BPDhk2H8IcSnuRJtxh3H2w9b9zDsYVjBQgaXlcr26MnztBuIQAGS
H/LAB6La1Nset5wGwVL/FlbeFlfUvwpWT9dBqqZ97xx9INav+wEAPEp6l+5NWxcUmFQ8La3ahb3u
vj/ZoRPhGRXK6lg8G1qF/DLUjcF4/NgpP1YtOlpAPiz9id10HmynuYVuZYVwp7LmP2PsPok0RJeP
MfHUfnGdb64+hfwNIzWe1Wneyw+V5DqX+204q4GAD9t3XJQo3OGyi5RoOoJWztdJwlwVF7obGnkt
y0ziSbe96BmCZ5cDBfe9p1Px36McP54As63jUI9S8FWYJRkgESrg8BCPL6xGdabDCY2URMfWXoxu
S/407K64XTb/JZ8pdXxF9eWrrefz/k6H/rptemG2FuwC23njqZ4mDIdMVHRuB/6ZwRc9y2O3XIpJ
RRe/j6zw95puq/bViRRRTsfxf7C09tN+c1dk7/+xHmyfmhhPpC/GegVBqWQBKspFOJ/xh0Ei9TkC
yuePVQzAxk+TMzCdDsXpCYxX2cRhlBcBdiEeI2LQddmNT1N0vCnaTxjz8uxr6ql1ecWpSBv8e7FH
1WMcntNyX1vr7x5sgLao0BUcDfn5DqEEaU5U+aV2BYLqyEFGSkRsDwn7KZiS5AUaYjN0E7I91roB
HJ1hT1EEpB4s6pdyglKkP4vK83ED6dKlR7mVLvQY9nQK8Qw2XufeRapWQ77ZUE7PFDhTHwdYr8dD
a2jQNhNDieMiPawTDH53zeBYjvaBdbU0CBuXzWFzh1pNuDlgTy9fZs1tkiVZiAKcVii5yTILO8YG
fECh9+IBLqwqXR2mWbfmWDlOAzF6UzhDHrfFGL+lZx+CNQGd8LLlfjlv85MNpZL7/D075Btj0nM+
veMpmXJBtd0tdHOqO4rILWbnADC66R4xJqhLthzC5zI4YFGnJdEUm/Z0mN9jeXzgvnwpw+N0Yqhg
NdPOlWBcnckzIGxXNKy72bgBnIBf9qvlgUhytjEBdzcZSrtb0EU0h68mu/PGrAZOEcGU4Mtt4xYu
1uF26vzhWKKQ1ktT9S760+fD734Ys7M0ZMN2TDmrbZYgIGelrg27wFluO2QjxiMlAzVDwL293U3I
AYJQs7nxEHplycpEZ8+nu8d4Zl737O/DS///UA/wlB4ifbAgRO7ibUArxv5HnT0Qc/vVe2vU7Nq+
ZY2XumghAQz7ZkOKrVALJuQ5isGk3SZvvGl9xZBicIhLyCcajoUwAmAFE1zGsunUXXtm9p1iFdJZ
m62fzQw9PnBIR0ybsBxjtee69NYQ+swGWGhAcanWM9uOe4VqYhLyjgUcUyaHhK5UNQJKnjks1+Ba
I5IrjJjQNeMra1Fkd2nlmXP8GOQ5t0V4oshRrDFIaN4y1Z9Ark4eatgheVykEEVDgLuUPQNaAQM3
ZaN4bjkAxnsk7OzmR2OeAgWknir3NGSfctmXttRQG4+Pn0oxCkM6xvGXA8oEqxbMjkN2KCVxgltu
KAN0wrPtRlXHbJUJbHu63p0bR9zv4tOaxJ/JU715p6OJ/qx1ugC5bK1rUgNF1M+cKai6MeuO7NfX
uJ4GSDzVg85SJNSAQQXvTmt9lRyo6BgRR08Ws4bA03IOSYCdOdkweg4jwewRcJcWW8sY+lgDgRzE
4qyLqVovg2py/F7lZgODvZy0X9zcQ8c1jejdATMY27/B9xsaj+TzuBawGkl9aarZv7RksfaGZDO+
yst4v/U47kpzXYe+fxjlgf8ZDXaCWvoRGVXa+WdOE+DmmiKBehIqFd9dMDeiKxkQdxqDbw8XsbJ9
nJlPr6mcixt3y11qAURuErsLgJ3Uru91SeHd2h65jjJ1TJjY8ZXqti3CLHkrH4qQiw3Lcqld1DD8
knlGbBxEaeSCkcUVX7ilEbhr5N+pPZrESBurE6EgflvkNdoxDIBXI1JjpVOoiTi+/lmvGNJvd0KL
UG+hOuRGgTi0S7FNpGtV+6N6gJ1AFhkcgkhdwnueftzjDET/lsXyY8pJcASnsd8L6VhXbCxv1z/4
Xm35zt5acg90kSbh/UEzh1ilVewwXDNKryTX44m2xhkwQ09896LaW4IUHh0OqWy2d+dxnBXEdWJe
LXFDbj0On3p05jS8pfJ+d/LGiJ3t8I49NxI+hLXx+7hJ15XWvG8GuSGQnITa0eCoyklW1w3UiwE8
ZufKvF8jHdg/ANsk8AfKzClBWSbAAidMWDCkfZP0iIn6NiDLB7vfwwNqzT7CiDwU9PEo78Aj33rm
NiJwIKrZGFS97SZ74H4N0+NZUmByLDku7RBYVJvhp5z3jf+aeAHC3IpzGu4pqlcAot19DexeDw0c
HrqgG5FzLJ//5uMffhNyBnbVZHChwXR85qMs7FGh83oK0Z8nQpLZLkyQPWi/wTRxLliyMfklC3GB
giZL8hD+IyexI0CLImNxDlya0xqPhL4EL5tUg+gP4BXstsw4tkuU+GpBnm+QUI2x5aWxHKYOk6qP
TK6mH4D01GaCYP1W6iQmAlVxE180u5TnPXFydYSzyq1lIq/kRxXOoq3dULqiSRkMXNinY5HMHGaw
DgpqgcPnDOh3PdhmBmkNQuLKt4wVu5xn4tZHBJS6QAYmDeY281wIqMYRp2UAuNBCg7iZfgbkqitX
NHW8ep2EfZWKCFZ1b1451iXxEEgQ5A3Io9AOHgx63+WfPpXF3eBLc5eGWNSqgghPkGTkBCzYHVYi
ukxi9nwrhRvUCiaF10EC0Z3AeZEtBZQ2ZH1N2EiD9LAAc5QAycKPRgJFnyAYmWak00t4syYc1kou
Aiwk4wVWUCKdeQVfIoF8Q+GwrkFa9afPGq+vuQNZ8I4tNuKGhb0qYM3FkPvPPxxNpJQ06j+QesnW
Jg4x+KeNCmBDBsyflrVeJHhCu0utX2DGx4k7YwE0h23JLgNB+Ct7n7maXGV/W3tfVoDuxQGSaJwz
RZeLAML1wbLy5ahU59zIa4feIHIYxFfY6N8WpL4nUlvc6SIHTMmhR0QuyjTJ+rVd2Ojjv5M4XXpE
qnkYxJMlvl/LbntOpaSQ7x2F3exSRM0M1gVoGUtj3EllUXRc0tLh+qp12t4VvlGVxNvzcQRHgZLn
Lcr5HnTykjKwo+/MDzrNRzz9oIqbr954FsNt4SXGfBS/59mFA3KFUTtNpDta9UdDrJydnR/ILVcO
ppOoj6jzgsMnlbps0rxLUSeKhNdTGWcr8igHBRWdHqNxGf9o2L2Nr72bujBfmi96h2oFic3gXGX8
Goc+LzfT3TF30wqMgtKcGvsIMXL/Vweavzngk99JSLU2rPalbqbDhFCTyKt0rRixh6xuBGY+4nXl
57Wd8Tx8gsj70jsm1v3nNh/8pviV2t/ByxvMyz/JTJOYE3r/BGv8V6pXUpBQoXEJddDXIrhByaM8
UmFxZ+jGb12tI5DvxfDw2dPq04sXDS4QaOMPmOy7aukCC705E7UVVD2r5ixQKQzlM74e2GbitWhY
Y0YtHFMcox8Eo8FlB6WqQRJgZkt6tmOGXEQqDxA87v8Bqs0cG/Ri7WIMEzwcq16SfyDHu1FJ2uWl
tUynYul1qZvSO82WnWjhkacPcgY8w/EykYrLXHXNNhu/6t8PwcV7625E3KN4NH8M3xFCHWUhNDPa
1+e69QzooaVgWeWyVHTfEgxovE90Bo1W8pQm6Jcw9SXlQCHDhNYGgQHhRH6dg752CSrxFUYg12f6
+NS+R2BCf6StoSNSZl5rBxVUIZIq/wm059U6LvgXqFmdkSNzieFdTjMLMsrsmJHTtAPelFzw0X+o
Jmqf7ZvjZWOiH3sJBpVhOXUX0rOYmpG4JiGSsqevxhlBuJlln4gmYdyxu8h8e9pWBBMY7CL2vJmK
0kudlYCzhHiU3DIuHEtRgGj17EdWiFjva4ahn6qMgrkq8FAUJXCHpWDQ26XG/6fdzg8epCAxJthY
Dd+8rmNREYnRzpfPc/5U8N+4y+1kr7mmNM9jXio+DAE2Qo3x1TPNuZB4Z3MW5HecJ+27fu9uCzDp
RvALjIIuXG8F03l57qWgqqL2FbEFE7WHDq4qgYryN8t4K4NQ2quq0neuSJP+XYv0gn3ASPfxMfT5
VNYnnVolEk0c651Dh7003Wr1SiGiFU+lBE0nGvQRYmKojllfg9qKIGwrNC0XHS0USk4hGSt2s16l
p6yAVkd5Qp4LQiKZFOG+JajV4nlKzX5BBeRQkn3qn0EMU5SS2ToTPZbuOmmixOP01kaATvsMckQo
fYOuHsl5e14Uqcd2jqE21JeDccZCKCfg2bC7YQpoLEjn0twMhIiEOcbsrUxzJlZlmTQEtM6sDazb
LbUVZ59wNvMvmTCgtAETfRIkf/gpJeLLFAnuG31Aaz6/4q1UAENSBZwQEazWuMBJ5SnTUqMEqgzq
prdfDQnFNIyeSWVTe3BQ0kLKGUJv/EsgX0ydDDpAvyn4uC+qYATPVFrMMi6cD22F95vrgm6/kKrs
HBtynHyZHnVBzNofPRht+rVg3VHHu/CvmaL2330/Gc3qH58lWpK1fYJz07AU/Vpyr+yf4PwVrTvl
9T61HScH7nefoa9oRrK0Ki+kcHZwDszYT8LhBx1bWocdKuz+HMd3rtWZsKyHVJCeQ+XCRKrbVzA4
bHvgE1wHmBzo8NEHHCa6mYMRO2om9kWjJPvgrHk9PxHDYNQaPU0CAtcUsYw4/vvyBiG0VQ12aWTm
fCmf8zxnKy9bBwEcv4JZc6PgGPomtwIjNtJtBbYbWHtuyiJD9XBI19rB1tn4NctxjyYbxQYUXb/B
Dq0xvvsr2uX7eZEIP0drKBHpgBuULOWaZ39pX/oTkr3cqmjJ6c7F5xHU1ts07+uveVvm8DzaKMBT
iTOamaDCAnSAoB40GgBkRpdk3AsUrzsRyPTIirUJijeOL26NIx28rWA248io9d42chZeLTkc/AFQ
ewuiCn5YXtBsNc9OkGm6vsJCh2iDNfm5AaN7PcyCktZRpAsv7v5L9aIHr6jHkXvMCnCYRz+1NSDM
AmHKJBAjDhJOesPLoH3Wv/6c765J7GqSvi1StAI3mi/b4GVv9FHlQsDGhzEhcQJTjH+/gR5N/J1B
x58YkFFgqjHKZkQrjqbmYGs7GFufhqBZiSkodYgbqOmbuBFNxU28gQNInROes4CRnS/HzVc7J6df
RV/vLBG9tfQYJoqtL0PfyaxIxyhh2WXzHDpkd42JxRrxSbP9g51ADYgEbXT/FHfaS3yYjrRgqWY3
veylipUTxO9fln+F9GhW+KWSafAPiRHjMgk4aWOl+kvmNV99Cfq8WN/Nv/KfnkpZZ594LmC2ZUK9
gwfWDrLMDcHJXN2YBy+2oNZMEJdXwEQovZEVmFJJTs/1YrR6bH4hrJPNBbbNukJz/D1jh8WkKCEL
HoidYrV8vgk0pEjKNmhMvVK7E2RwgfqOnLK4yrdKWIYpmTVQu1cd0QgzOAqJBfCk/T0OHqptLm4u
KxAjn82N1QnvIwfymXiour9KPgXUyVFb33GZxc2M6B12P3zAqmo6dQzzWZKLVKCBf0lYQHX//7nH
zDHNOe/xtqMgBV0fSIGT2fNRIO8mR62F1If0j2Yfn+S3pUXxNoqKatOKRRco+7/C3lVXoiKZXJJT
vtWIMlGJPOeKl/TX3MONNpqtz8C7f7B7r1KMQIV2MWvR6hw0GzC1hyRxUop7bXyixgkH9mwbg9to
1xB+yZELXebuP6L75SHzOdxsiFCpIRoVIdlw0hvyWzwCHuWEGz6uWm4bRsaG7dlvdFVhsqo6Agft
nLMdjvJ2uZ20rA8E7/pOiq2eHpuEvKJoqP3wmioXyT7bhYDJlyoFzXvg20FAimZnqgbxwXiLTRUV
pBDgGmxobPeG0KracYyyMPqnE76MsQBH4diYp1G5WdU+XGhj/WmlUFR7N+7ox2FoDBItyHphu8Jf
L/QazFCM9JiU8i4Afu2T+2VRBM1XamVXJapu8DDBANJrm4F/NttYGh5YJmHaGNeD/GZVWIKxEBlz
Dn2AwByiXMPqCXji0xR0WjeDKjlBLM7/Dt9zwjpzwDPf7BJF9a2flGIH1U3Zcf7cLnw59/qriZUU
10OTQ16kSMIkUYcIQ+dgH1QWLlRGAotTSaGehtrogKKHEXGNFF0n5vJB6xsO7Bf7hVKKOB3i0oW7
hcJqLL2ijg7X97L4x6hc9G3UWHnyep9XWb+0vg6UItkySxnuOBWu1ID1ydkAggjcmUW/IclUV6Lq
WTkvyQb7Ejgt/3QOTlKSZzLVNG4PBOOMtvBy1j4MBDuvEfoDO/grLg+9tmrkNyQG+VPQx8tvzXxi
MPwkOpU1hG4cjGxNoEgV4l8yEwVr9W9+EfMLYVrsJkG6cofb9wyB6jsYR8k6GOHo+BevyNZV5pld
DQsTE6vI3bnuDv564fxyomWCVO+ZJDSHus/PWXHx6pfarXxo7QaNo7fQVPacBCA0ThvmeloqEnqX
acRIhyFy2AilXHZ2HsifWimyqbDB9cPypVIVbBeIrbparPiKz1nh8jgF14MCf6VgC9E7h9yOgjyc
BFBQ1Q6J2AFF1yjBR5yxkWKAeDRskBJzK/trZLyaarRUBUaYP59NcZDxWbCQENUfZMdD+s+yYvd7
ZgJvCI0/mdCwfzbwcfO7Sgokd9+n8ZcI9EwJZt045gihAeNy5f3BPbx8UESKTI0zB5FT+tHK5l5F
mFrjyIj9LX5lcUXAtPP7kkTIwmcELolXoi8oNCj9594cLPP04vgzSlktAKL7YChQz+67EJIb065+
jFQxF/W4DlwZrIIzqjIw8IRRyx1WPOxkRD2WMm5TkUTBNviopdAjtT5XGHcPkIvsBqp47LiQIyLk
4iYcsO+h/3MeZhgiNkpim8N7tzSad2/UEL0X9fbT/mmpENeQXhgm77Qyn5Fnh3/N0rSqVvs6m9g5
bvGu8dJouMg6IMQtKie7o933jT4tc1DkDq6Bhq59mN2VfZ5FqgHXqFmzsN2ZJWeGZPr7C0ZgUIs2
sc35lsNKtYXKmVkwkg9L3kiD0MHiQfM3kOnJPSerb/81AkE0qYrnviJgejLmUX7SApiW8RquIrrI
+cFPbIOxH+ZLqtPQfi+0TRM8PzrzfW390lNgZojJCsBNe+BTh7ZQZrcWtgjjb0iJce5K2mjHwXhm
Yl+qAoBTjYY4lhepPbJHVSBiK/cr6bPLjiy9pIMQGhAqKDFVNsg4NPRUXnYOSB2rqIQguWB7ASSh
mbyoQqGDxa2L+xgR/KSw0bUelJdwtqTJC58MxKgQAPvM21Cjjz/hPEvfhu0YEBrkE9vCcmKuU9IC
wDfjCb5kJEJ5yaorm57oZrMWDF+IJKhmqDc0PGSdXA+CSLUyno3Zb/QJMYlobTe+0ZR1Dp3Q7fBZ
P+dD6Yck63OD4S/bQsJeN06klj+n80zMfdsf2e4pAyVkNnHyQZZue9ma3eAiLCko5745Iw4HwaCh
Gvlskp+WWFya+gso2FnmKY+Ke8lrBtIienucK3PU77uqILCM98daU3B2yYSBysS2tZsBxnc/AeRX
FmFyV6ejCn/TaVAIBeCeNq2BlcgTfyY6fgiJNntLhWTZxhvrqHwF8nTCDCuwb+IgAW+W8nntc/M7
ct0zCriy5W7UX7fnJc7bu9NPU6C5+H1MWP9IlHGtIsiLB8LJ7L0My/a12BsCWa1uY6unuAWCvG3c
PngoZiIl6re19Bu7AuTC9XIGED3Nt2E/9TDbAdAZzD+JZm1hI+cfAipCw1kaqs4BCCPQ6+L0uJN3
6aVdSoEoputMfGApW7cJqjGRioVu9kT/QIvA4v6gq8LYLEgoKrZhc5OSjwyaA6rAOOYjpQVjtCRW
WqyEFyiFe3c7LO+pT8fnQoeSewFeB7fesp8Y4UkIkdITa445KpSdnyMakPFuNeNOrpCvAJBOHBA8
sCXL57GgMHTWIvV1CaOptUORR9Z1fusUxuzQcjbpRvn2k8eMELj2xxf3+FOqZzmmX1rikbORLv2N
0LW/X+njUPTxxxABg8AMWyDhN2f2NiSVMElupPtFgE0CGdBufTiW37DLZVynBI8qqle0w33895xd
GSPAfbTbObVLh7dtNrjXK2CgpLBa0s2v+eGMurq59USwcKaWPnboawf2hfaTRBmP+OiqY2eLx3Lw
Z5Jq2irujGb6LytxTWlAtIp/acZGEbDPEyH/3qez0P7FIWy5scQMmiQAv70NhNr2xRqqmFwbCUEz
VdMrHwfxFBgJrHzUam9bWLAu0mRAOqIB7pS/yaowbm+o7lX8IpVxGUmsY1U824A35FO3G3FhTsuz
AJgSSXhpdiFKISyAhgxNcSbDb7puV1aOXwHWZ96KF+BT2qiG+gVZz6OlB7B40ZuZv65lZaHlYbyf
ZsIW0yEUjvh4AgYdySwgUZvDt85TKC5BGPnjmELZSzAnBEywwRnlflaOXKOpK5GqGhh8iXv4gW3s
mkQfrmvYuqnMxSg3z6CDz+QCu+P6i0Gu6eLCjPlndwt6w6PYLfvV+WgbGwSH/Pl2lKnnX0SOA+hu
QE6t5B7weTjqJ1Flu2+9q3pl6v53NT0nKzPZ/emegC19ND+h9ciTL0Kdu1eyhowyhFRyQsDwcCzg
zPhOUK/AvsyjWuV8doQlfl6/WV9GQ3p9C77S6NPfOaRaan84LpZfX1/VpV56k4TPkTUfMtyp34w3
AfkXlqH9VF51HdDVGE9Smj9s18SCjadqo15LyLUiPbdfyutjkvGSdCGCrihFFQCSr4SlchMD67mG
nIT1VLEOEvibowC/89yvv/+b7BdRcC2+txuA5nq/MXvUiR4l/KxZ1lfYkIUkScS5k42SgePfwa/N
3I/UONLuVB0xE+ve4/I8plrcA14J+GDFbBOjZ/U2fm65yQPbPHYuhWE5bMvf9b9E05Q3GES16cTf
SicEfPZLQUYwKnX8Xx7jJLpuMBrx6oxuXs9TtZirhfkmscJdhvbFOq5Xy7ixcHk1+RZpE5vL6DiR
NoDcmAL43Kmzm2AkA/VzIsTCheYDciIf5oUs4HGVFzB0pmr5fRJK10dd2huxHT+EMZQZbdbHs4Gw
7QctbRBr4cthPc54eUfxN6HpEuA5LPmyLFoIoyR2dRCcUQGelymtsZy3yZzqbi4Sl2LTtwtPO++y
KjhE46A1yFPRzyt62zRauUyasNSGJkwclLbns9lJTsxWs0i2rZ+gXljVCv7+hGzxixb9AY5DUhDT
iTsa9TF8y6OFw/RNCitRobUrMlbonaXuQ5UEEIryeCZPE7wE0P0vLLc/K9svhqB6XCFUDD0Ojx14
AxKb6NXBeK+USZQoRybrnuynlKOrppgZ5wGDiAhjGQGWcDFhfNu2qQkqE7slltuC7tACZZEZvr0b
mwCPWt7s4fgHa/2HtEak30WX+VcOHTTSQBpAW7SFsQXuZszW3UASIbZ53VAEv7H+9rt8SzDHchS6
39GKS5KmBPKZMZqFP8Yw5e0Tbqe40YTMp2mCiyHniR2d569IPN/SOV1Ldn65+zZf8kYhx12NTInz
pWRYC/6YWgvbYkSXm9lR3TY80UwlS8NgLmhBgYFxb+7IvK72gBfHMGwVAF2J8hqTBLY84EDIKqT5
bMHqyO7nixgnSXK2up+6X48idON8E3cXxmeQpoXM9ardB3CalLqRwXlOELhV63R2Aa81e+5JkVgP
vyfy+QK+2xTR7LhnmffM9UPTILhm/pEzrROxUvZLYHfljsxANqfjlbPPs4XAAYMUK+JLGZ8QM59B
DSZZ6YPLD8NTzTcgZtOjSxpFiVxxFLEd0qi5hTVJwIhYIH41ACGdUiz0IExDKn1BI6EiuyAPa0o3
mu0+CZXz+wINlnSSz3XSEID9ZgXLHHbS9lF1wRxuPSYy4WEz6muiAHusbccsCUmv/BbUkYX3ZQsP
mZwI7xUvYit8cEO4gCCvk2gp05y0yZX6J3H7ZsqyXcBnP6YejYwIfehtJtYbkg+11lagjhx5BkWd
n74zxeCnjxGsOrUf5FGh+XYpysALnOHnqKdL0G9Z7z3WHT1O2jSpZsX4WV8/tlOTQucUDiPFafNK
Uc72cJPISZAyALZze4LDNUvTnnTuj9dYvdbeWRNEANURsTW1JEkF6m04PaHXyFdWhnLvLgo+4Y+u
8iJOyt8S811lr7IRHJdezGeAzEk38PpOlFMmmOqa1egh+DZM55n6mDYqcB5uC9fWl2URFbPRAbgL
yJkhORAIrCWaErp2qDahvq56NPMmn7aHajqHSoZ+trQJCXYP9WsjOUVkMC0ttbc9A6pqo9VD2UWd
J4joKjH1br9k1CxIhVhZVAw+jXAbNFMBeJiyWV9SsryWIAyOuRTGbFnxJ/yJWbf27fRkPgUWbYnY
/cv8KIT06zWqmrbNruB0RwNGUat0iHqTmAFkVRua0iEKSvjvUSkea/C4wv7f3SphZnR+p7kGvT9O
LsVFefjGyIsTn+CGwaUVfNW5xRCwvvvziDy9xJzpnIVsVPT4WcTLWDeKLnXoXo+JrHKXwKfK2L49
8TljdqAjfofEmKXFGUh+S4+WtNgjGc/gK/BxKKiWPXgqnZTVe4+un8bnCDesd9FbMSLeMmuzekvF
dhkKXMhDhjzeXmzjFT/akkFVgmohjwdJ8KQRtgxiaiDDITH+dNODwPqhp+alhk+X2y0DTUr4au9w
llRsFfDUX7J2V8PMofIw65sP0PQ7qhQdJkT9ylwFYgOX40WV+J+u/CgVxA7ru5231Wn3VSl3OeXq
20lKdcdR2XhsvhBsuIy1s1F26+v0rlBvdhlls0vZ9xME2ptfxFDlIpqUXK5sJzYIFMgX789juDSt
Zwmubdukszl0Rk0zTxuNjo3NNrVbHwaRIaU4nI+L3rTdUEEewKZ2EijKFOB6JIGAszFthCCLc12g
xVNE4SJMlCPSYKpOFaw3N33fZtSNIJOV39A+VRuWR88V30/A1sURH44jFA9sMvWhzmp526BOLMl0
iYOXZa5Xt5zSI76hrUDxLgY4jiYKFNwgAGQuUbDlGSAMrP6J+iH9bw4ZDYhnXl0ZdW8Peory4PcV
tnVgaYKd2jC9xxz3tPplyRAtDVgeFLS1WubjOefg3yBIajAQFbZ13yIoXUv8XMkLo+fyi+9In/E+
5viHRyjdOWYbtHdzdA2IKcdwatMR0mTjypgLw8M4yMDJ6KssJrN21Hr7l/arburCbx9fSkg4Vqlz
y6t65nAD1gIIqf+wH5wZY62nTm10DHrmdx0t55gP6b8g+FQWyAe8r9gfwBj88OZMv1HkT9OOX8um
BDUJC1FabkhTZbNL4BWLWhaxk9QUsiohwlfuFIm07UyihnVAd32p6TWWkDYxPypV4awPznKuyIpi
0O8kb5HB3fjtSHt4n9hxqGQMHpzBy8KwUS6tLWCXC7rmLY5mfruHlPcSmd/kGM1x9UPSgBdTLhne
Z7H+xbzxC/V1eXUdpnuvHLArHQ7GzxnZmJt7acm+UGVeXvTSDA8+jo4+jKQ33FLH5lkA+0s27mc9
DnOqrnuegKb4uBVxcmAvEEb7IUKKHUhmdxbAwRHZKBee5r21ZPpif/3YLz5Ngsj3+0ZVBQmV33MM
klw5OoGrc9ha0Uz59twxad6VoHTbDRKepmgtQER4RGy7LFRDcBhaBe5paaeRlbs+Tvzfd99W/4I4
M0ckadX04G0KQA6kcTNk50a30YKObCR5ywq6vqVRNNXS8/jT2TbkTU93tc6tDMRumMR8En9qHfeu
TxgZNhB0YwyhGwIl08p1lpEO0Z8WidnKzK+fAkzqShnJ73MhsjAPmsQ5/m1idlkhx1s/TmKoLSzz
K4+D7YljYiU8JbOFRtOkcIlSNioqYLN5fR98v7jlhY96lZsbFmdPuVAcwOGyIVEqq7R6m1VibGYc
lNbPYum9C7laqZ5URVfKySf/+a+sCXo3u0pSTsSo09ZG2CvjHsjVl5UDvIWNsH6iphrCZ8swx0R2
NLf4/iWYQ31dWphCWzIlj07E5cN0wMD5Vaz+5X0xHpTedb8WpNmYR4aigTnk180cBlDlVdRIE00l
nIN0mtR26Z0f9yIaRCNeGKZJvioMOkc1myGeyrOgbWsa68AUUsep54Xvex96o7mp2VgiXJ8GFuQO
hp41zb/lHls4mNYKmCbYTP48X6Euh0KrgLDXTm1cGBKnVLFtEGA0Bsi49/G+YtUXNW1ueidwobWe
b+qSBsNbwEvcvy7qVqtE7ZYC1vAk2enb8A6m2gwnSPphTx5dY7Ovynym2CHuvcZ+p/1QQmvnKuVU
0L6vgeBAOIbztCEp6+kAx5pxbCcMz5g0U9GjQWSbaB7ycmCX4NfWnu6wEMOFak9kf71pGio3h2Uv
jtKlUSfSZT74NuO4tzgxOs+I0E6GDv18rPtPY3V8Xb4B7gRzw1TUpqy07lbGoYy+M9MIFnxxRrSj
02IK+Sj9KUz9upIL13s+4U6cjFYQei1Jx/akPrxXhUgvY8TGxnhNe5QvN9x0ERrrCrKDGERcBgWX
pMrV3hrsYdhwtjkNxZT+I/eyROjNqgAAOHnJ8wo/YOYP/kKGrJI/WIdXgBwcUdnq2UfvfO22qK26
sdzuTkHLThRh/2joymVOpBGP2gYwP2FygPXs/f+XOykYex1EvPfIwvJq+T7bxdF9ZLdjzjAC820O
ThkbZfx9DRLFB8ySQfTLQWmmmi9upz+TG/HAleRmreNWpxTBT8fIcPqn6RwYAx5AfIqOPr74pFw4
AIxBppiVBXCwkzS9N8hTN09SOX0IGDK+ijm4K2PUP+CZwHkSfwF7rlby66vjLbuOjxyGxDBLKW4+
BIhaYxmheSjHmpvjO1NkOnudVxc+2QRMkd6JUq6cNMSbnIn90N+04iLo9VRe6axSirZeZoQk+sfc
SXQYBqat5wsoyCva6ZRjGHI46Sg15mL13/10WEHsBvXkJzOwLz/dRf+eCHx/BjIO6eikJJeoOMkX
DVhJD199sU6lVMVUJcdMA3Rpgq1jH5+8UvyAddjXEPEcb/p7FqPYY7S+iiHEA74zLoU5Xm0vStXm
1ZbpE1c/Nis2mRZK5RStbDxWT34G6S5zRgecIAXWpq6dyhKyIcva/kRTGnXnZIb1puTqA8cVaBJ7
CxChzAct02GmyeUE2QEwcnXUa2kyOMpRNSoD3o8Du9rrwFq33I2hhDKqSrGNJCtPTfNWctGqzluB
yE2R3RS/3uV4NNNHKE4faZLpO+m3sGhvWWFKVwQqPxFNhehi/fJRDYOJJBDxJhbgKLbbQOaNCaRg
K8yzYF0hveYnslKgTzifTrj+qtB5dGYSy7h5t2qnqAhkE1V9aqcidIQx1aTvLbiJ4c+1DxejPkUV
pGt1a711V9fvJSWM562tqTzni6lkEX8Q4+beDaneyGcKtJDEUP1+A7xVe0BC0yKv0mmt8z9xBXwQ
nxUEKVfzmpGZtx2MC1iT+0I5QWWVTLOg7X5SFl/rulsaOqhRze8OmlRATsOJ8OdMOfoIgDxW2fGP
KvINoLoz23+tUJlLeAP4+QFFeMlMoJoSRLzcsfTr56oFHKRAfg0Br/XTMUSFqvGXtfwZ9PMiSbzN
PUcXhUohXnRAqPx+Ttnl4ZHkKnV2nf2r81QGEPPWrDZUYnHWPi/LfXSeoP0M0Bj8xyzQYlEPV9cz
1hEXNhopWHuWFqPGYOxiTu1vUV3m+pviNxDIUeTBAPyzvDBlBMbUz2HrdpfLosO2LA8euDyD6WIN
tQU8UzwmDUFaNbxcs1Eip+rxi2oTE6jkFaBNjDdn666V8SAA1bRmp0Fq5uJWSaQdh7Zo0f0B+4J6
e1S7aFc5xJBogMYfUYjlX9fz4NKn3d35Apl01N8H/Xm+BN3vlFHByEBXhQH00JIwOtXCR/e1/R7f
CwvIekwdNjeUnSSjGhNHZizMoYZhouwpl/hzQSDvgiHhPvCVV+ZArjcN0LX6MassCaXBXwW6eKmQ
SuWcHNvtXjLVIIatYm1KUKToNYzzqow5AvxFBPSLuXRfRkBHVtCL7lVroQ/EnSNmS55M2R6QxpfV
AI1FRIcyvL4Br01QcKN7dHEYq2JFn+azg65E/Urq63i9Xyvlwa2/pBDMbBCTysQyHmTV8LE8dK91
dYf2WomIiQOUI4vdZ/bf1LvfDqP8VwuBVEPeb3cjqwMz8pCZihSeqQa/oXAAYjWrpxSKipDj41SB
dFdlLZCukWd4tqFWugY7tDn1iTGaplNvm6GBVdf4cmaMz7YvMmpDyERXEe9zR0L3Vd5KhWXyaVUG
Vu8Bd8eaaiWooVyDTH6lmNqvzYdMnSE3N8kp5w6RHXwqeGaiBCwBZghRlxp0hLVCBrtrK426hvMK
3iR1+UR8GkU0z36OF2X5Oa+ovTzQ/i/rszrwn/u1XdBAXL+5TR8RxH6a9+TX6yE5GDFBgFExrhos
I0A1avgcY+jl4UqbQwOgqS6YRqk+68K+E9dd52ArS4QWH2hj705VWGv+MDZHpNgJX5+ynjwi/roH
C1I24jThTUkDOtGnslLkD+R8in5W3nigbE9k85A+Jqz78/DDl9AzzeLXXuxapKNVRHZYvX6Q0otz
jXbd3yv2sSxxMUiACVOSUA2i+/vZKsIZmmYFwc5S1jFYDaNqbt3jcUBdBq13FlNLrPj/nL6veVdF
qq+ob7brEia0zafRi8Tboe36hiWDyTsXRZSZ/pzCWyCOxoeqCURwEJWBLc7EjtVohTG60qtyMq+9
2PadRzRsmOHbnT8d/uGesw9V4E1M7V6alR0pcclgN58A7s8juIqf/TOreDxwUs6fXvq2N8q7yvz7
q+NseGU8JP219Y9+XO4MOkGjhPcgVnLdwG6hHnjHLgEncckPLO7MdFY78X2BjF9A9kpS87qjwK2u
kkmsEIo90azh1YOHO+yUuAGKWNOuX9gFctJj1t9962W9KaaQT1+NcLMb/8kKPpit5nJ+Hj+Dpk9Z
5668RkIlHvxFXYyIU7IM/MlBlYySMbDwoR15vcvqHOxVtsh91PG5O6F8108VQI4ezg5ciXPTe6/s
J4O14T7k4rr2i6NzPltim5/OYuILxwXpDb2CSw5xVUfMejhLyS1DV50blDUg/zy64bXQzkCGxY7J
C80Z8NbqtqvO94dWSm9y24BSDHuHs0QgoH4qZqydbamHayNckY+hW+AU8SQm6AnF53w/qMLX+QRp
MVX9u6/sR1nM6JICu8sYO5vvwa4G51BbpJerL6AGy9Me0SjEsllWZH9m9c9E2JfqjCYV03SrPCfb
J3n+mwRSP8FX53FFVWhOqqwyBCzhXEQaJz7CSRjDT9q2Y4Wf1pTc7/AfcIiLylW2zwCrY8O3QeNn
UK4UtZhjtCcIH4W1h3IQYF9uOAPelj1QWZOyDInkOq16QlF/UteBbW9dcLvtLO5/pl9lAG8XNCE1
C5qkCzZpu6fxjVBZO9kK5tY7EICFZWLQ2PF/Qf09xG71mRgJX1yPcNgk78hOc7R/WwDLQxpVeExy
tS7wz5VtdBLecj2ss6DHba7XLXNgNAY2PekP7W7E0Xxezd5faEnAVSbT6xGwW82+ocLLIzvBZZek
Z/nqTcmCMDkn1xYYuHO/UF9Q/UJnAX/I5g6yeaOFUUizLpTRyDBazrL7kxEic5vQlWh3L3H+uhYY
OMKOZe3GH+/j/527UNAUwYRVtzXPYl2TDoeaytIvdmT7VklReUhkUg5MwixJJ4K+b0Mm6b3EFK2a
WZhlXgtXHpC+P+DITeuT8OZ8aEPeb/qoxluYvt7itB67RMV63yiMp8qX1fRu6WKBfyIOXV5CWBVe
EXRkd0rsImxZXMzT8bN2BNltBw4Tniv5K2iHWwUhvLeDxEVb0rm+5fmCt/BsklY344Dprc036W0O
6M45/UE3F0iEa+HEIGZWKuKycHPabxZrMxz7gCB1YvNtfawDsMyTOk2UlZGNyR4B8ERbbrbqIvr6
8GsWXazuoaDOmVryP6/2E4Yr8I2LXpf3n0mvLDi8um0OqrvYWpiRQgoWfdwNoJh+xiKBinQf6/zz
qKqx8iHR/wG3qqot0FCD3HOBg4totq1RQopFMi7P1IjwkiGATGmDj8wPIru+csUdTNQpyD5OIyKW
AXmp6OJC7MbVTgpxykq/XHnQdO8RStDnHeszgPuYj1ldAZbrXHoBnuGEKgFJb4OI7tv93kddN2KZ
d4sr9vZYeDIUFs4WvD2pl6fgjvwCaRsTcsVsmSMuGYFt4lCaX+QfSr/JySQDZbS2Ceh5o2nRiRmU
IrZdiBDnQZGmas+/aFOknrN9WtKua1FDYPZGmKg4qKTphqVsP8s576vo6txoaotDLcL2EpuJb7WO
qipf5aVmaDB+Qea+PwzEqnxN3r9rDqvfox4I7X7J7cPRCxKptN5driKtClkMIZvMy6gnPqD0v1/a
9511I8deYizCaAJk5zWT+5jIMOfEUb124LwNHUV7Be7glsImGxJ75h/qFhm/nl47VKBBArkdCiZa
WLhffgu/Pa9DNbnNauTN/Xb0f4mLqVdt4mmrGWzZHokjjBCzlrXMOex4MqL9jYebA1NbswnJPs10
xehDv2kk4zr8Auqp3DDBlUCAx+3Pji+icZcRMVBj+uYLgFr3dGl49/T2wt2kqlszjtJ5BDB8cJlD
j+1dVzlk0X+bVPucLmS5XcC0/Vf6DkKTbmRUv3VKwKa52t4O4K461wznpf3j4etDnms9grtUvQdj
5TPern8DHQ4z8vOO0NC/mwaIHjIe/UIi6Rpj+WRje/UK4QUtCwHCUwGCiC4hhNLvBXql39l8ghHr
sq1sFdNrK8ZaOXrmUJOjU6F61m25njjnV1WsgsYpWVTdOw9ognBCNOp45Wtc6AddPZKsnzQwAYii
zZlk5dOaSk7p37Sa9mb9E2fXn4ZOvnpltobMWWHhRsGQ8IE46LWP7+gEqQQBTZIs49FZeaGCyLue
Q4c+UMceds8mHtJHCbqQYFPBOKxZMBBV3tDHe2bGcH72C9VkrxP4789GnlgJ77bB4jV/guSaL+JB
DIHT/TYQIaEpQFXIajRY59/MCkwZi9nxzga0ay7resylZ4yguXtk5U/wRoezC2K04l+rO4n62ieg
1chGH1F5ORkQSONZZJfP2esnd+GgNMUI7MC2kJM3aboWqYH5u6tmpMIqKgqVfAm7NveigGsflsgX
1MEx1d2c0DaYVglGikbZR/w6NmX17UxrrWGQ5d4I1UflSrzOLSivGnWOZP62zWYkd1Av5+GlF5V6
bm9TdbYHzgy0CPcqfLdwOQVo93KxyRMTlO7qnqbcCqvlnNqf5OX/BbJOxhX9vxMGDnfFAybdD0Zp
5rNsp2sX3WJZJocUccvVrfBUJch5cIV27pdk+NPcSoVkqsS32C58nWLTHSBSN/8QJHku3F3VMBDp
gjIucwfca/DQdrTDwYI8PpTlbvB1Aitrors6oNjCs/HWzzZrlk7P3GvOdrH0o7obZRcywRyGb3Av
PEOhYODsssdfXTKa3BUulJ4Ux0pILXEdXtMS8jHhMgGKO2kwadVMjYx8MtQKPj7lDsUVi8mJMhV8
EcdN9qRUz5WHkjx3tCT7TS9eGpu+WCcP83Jja8JLa3GySCJjzZ2jN8f5eSSi824R6jcEJzNVCRfN
FWgNbuo3Poe5YI17LxKXeYSdWFiTH4VHNit/Ar7Yo//eN8PE3i5phaK9uDeK7GhUeMcTm6Gvvx72
2EleE6l2epSazCbS/seZtr4kn3kCT9ZepgP7xTvX5Opv9IQZNMxCu6fklgQOI/YpuoWtnsGJ7tfs
Gmbqhgto6d6O59yARE0WHMw3rRJO8kHj2HNz3x09ofP8zejTvtyae6RyjOmCNqTejVSyFhpfRgio
lKuvamOIEsvRrQA5+7kO2zKB1PgpcYBJZk1ikZ0j5SeLzK20IybFxBCDfCu1BEg8deBBeKbwLuRO
wpG5ZWHHLT3Po0BRGdohnUlJICrkf8r2rHxOmtayFqWRIxBLmGA6zosKpkHsXcYdbhz+xXnTbCD7
XWX1xAHJ1amu2rMyAKdCYeGPn+We74zBO6U25NwWA1mGFriKZMvqvLO1dFV9HV+dPqwG6LpcypQD
nzHnq6NxMTwmYES6pwcA79UgWTuc8WeMCMkFB6oeFhyX7fgM2s/FxOclNFeZGzFayeGlFLWjZfRO
k044FurF+kctsXBvA35kgVqdQxEYgSVPX1B0J+NGBZmUlgNynmOmHeOLyZwK64Q0W+09LWmtx/sV
OJJWVvW9fT3glZrQv33D93QM36FwZV+q5cydCzi7gvUU48J8kLRZ3rPHHkAXhYOsLDJSd+UgKJWA
vuuGd8SMPIfmIE+WitIg3Y2nKtYg44ahIe9hhupga3d3CYVEzWvnrLzXECGOCnp+x/FwkI9MRyOR
Ii7Me5hYaSubIKVt8gEK8y3lDS5u5U/3xB2G5tgZMh7TtrnLpm/tZU/c2Kh7JwHQYJd5KNquSAMJ
tIONvTsPs/fpb3lyNHVDN5F/zW1nVQheNzn/emr82gZaEySfKYjf4l3gWTU9/O0bePhg2vK6uDJr
zQu4VhwL5Xh8O9Hr0hgUw6jjpO/8Tg75AOkY4mXc0V8+5uWXKrq/zH0SdoX4mxGCENpRC17gCsNP
KdKAk12Ou0rPlBU0r/NKV/NOOTZjw2qqhBl8ZjIYeToEoDcJ3Pc7eUMihNanTu55atssWNgOoej3
CTFqsL085WGQGbC6MC83hOAyHYeKLlt3kS9QDe+M7aDR47KXyYD4ECzJhy342nXGGgp+nGy/EBw4
SfOdysDxofvbKnelxmRKqCdngA7V73InGTWBNmWGJNPzBbGcN0yP1lwdl4J5Xml2H8UYdRP8jo5W
jgQFEwANfsreQ4DNzfowr3yuUz680tzOF2nGm1XAN+NEpXV9YRWnjCqVBTy1KH/3hI4z//dzqGDQ
MX+MurE2YQQ/XAJVTRAu1ruD97LV5ru7ig20ZxEV73+7XdgYA7X5qba4f5Cs4t9zn4OVrxOo0AIl
TUUMTdo9oJNbwbXK4ZK1g6+FiMBsSVpsmIdJ2zJTcQf+LhrVdXa67JNEMeWRFtF7eq/7JPx6qowN
O3xwpoJXiP+DsdvNAYKt3GaFLwutx3o5QHC3SPoORLDLHoKZWDOF/6YEwLv7pvI5gMfPi/MXBmSQ
ogzj9iYLTpzIJUfdiU6UZ8I9ku/QgCllbRNR4FB9Su6n7SfblJylxzpfxhFNdXy7QSv3bOvx+4Js
cNTvQ9v/6N0YwGGoXoOEV7DF5H2qIybQpGoVxsBabtoSyyk00NO5dorrfj/ih3TPDBu1dJV61qoE
uLdJVUHEf8yXuwBCVsJWq50xOjPJC8XgQpb0CKSkpbAEVFLq10q7dnSwqeF5B+yzSgQI5f5vzxF3
FUAEJHe0uLaiSXxuTpT1hN0j5w7ooq1TBKwP7puzJlhBv6/U5Xfr7/faAQCe1FqMg180FEiiTBeu
XBsRsKAclSCkXRQoL4MSwxuoxpPr9KjXszVHIYGu9/IFqlzXnarIMQx4UPZ3mlgavh38PaOf+fxW
KB2SxNwlOuqazfn1W0qI7Z6KKCTbMIHFhdS1vOHRfZG+WWnsiCzv+Pj67Rgof7bn2souu4LR4H/9
8IFYglTn1a82mG7IOs+y55aUtAWFFa0SoNOl7BxLqdZsw1yFh8apqRAHaeuSarpIKbI457RBY2j0
/+yT/94JoJqkGS6YtwNwYXCi4VxNyQc74ZyJecZEr7VywxiJJuM7xltWNb6yEvbM/BVCmYdqICC5
qyt+lvJMXUuV1kPtsEgAf+Ill2EDVqwO5g3Y3Cb/XzT8bdEseOvwOzURLk/anAqMSu9MYAWgchCB
70SDaio289n7n4X86mvLBFlujne46yVx9HTDzNtFV7VCGH+GIMzJmOcnLmgL1t8nvg6HO2VCoIbv
TeMHtsLlR+aCA+SPoplPoWe5Kn+MQVtbO55bKKx8tX6QfnyaaVeP6hmJjIbyOE6vv7doKzZXwqkx
fIYvfHUGYwXpeUERx/3SR0k0+RMeWQsf9UE8Xsyhf8fxpAdU071LnoJbiai1TEPQuonqepikMd7D
u3CeZd0aYK1tIa2Up5lUITNdYh5xI/k/FYDI9VHRilkP+O1g6GOgwnkSxLh190tgmlTodmr/nfKv
37776D/R7U9lxZBeBz//UaEhRktdrEaGdedQM5YqF4Ott2selAgffmTDxEua6xX1KPXUpiqWalo8
EBdGO/Tv8EvLCLxh5ecvEQHvbeuzxMah50ZU9SEQ43ZBRPpX8ujYfUJ2DcklGeN+4sEMkoOf++/9
tU8es/lxYwRP4xatn/qy62NuUqkd7rEvo9HW0UA8Miq4zEm2HtCbm7rcCb/nYZ5HgzogZ8ZZcVwA
pj49J8MVRvUiKOYCncYek5zNll3KM8wddAK/AQrk1z06hmW5cleHM/QEZJYnHh/mRldBtxUnMHPy
wxuTw9D/9lX2QEd+oq+Y8R65lle6ZE4gFGUNkp1DQX8Nri6O0BMq9DkjOFRrSzdQr8J1Tp+xbXP9
SA/xO6i6lbHyCfXUpaWBI/pfZh8INbhrOit4WDSFCqnebuZltJsYhMHyYukKnujVBLntbDN1GDpJ
Iv3lNkyxeQ9neyJOFj51yNpjYp/ef+S9q7LjW42D0zB3PR7Xp5dx3Svtldoa1DNkq1ghkMvbj0Ja
zfsxSAGi5Eyb4QbSDX+xvnAZgcncIp8ME/G8WQEAzS57wf8deg4a2ON6J9NBZY6ju7Xjw5EnruJ4
2auWM7/daMgkz0Nx0x11gpJCiGYozL01o6wTbXMMI5tn3NyeNehKuh5hqXOUphKEWUIBQR0e29J+
Zx44NSCmIlizrQCl/mgs7Ei4O3gE9hHYEPETSIJbm8qCvO+3u4L0UFLlDWs6zWgRrQ3VTEZsG9oB
w4afJ0oGfzeZw/6Ur8/ZQ/F9SZcpT/zxGoZ2b7mwNkorXOzM8B3Yyf2itUNJMi69pi7xbnFTkwkW
Q/fGrIQwLx/Jk1YpWP3C/3GKtXisgAhB3JHOUGv3uwcc9xo786IXdWaP8xzesf++7DH1RHS6idIE
O3XBLhsn6UQXg/yPXh/pUyI/sPO/ZRpBz80myqxTMgmO8EOWpftKd5ZlGhrzWXBZKtNRdkPGYkl6
Cotlv+b1AUkdSYlCzhLJ3jk8S/5bVLWcXKjx7ozOxtxWKe0Iwv4xdnE1wctQ/+Kx4k9F/GaWGFU0
AmzSMlBhpktC5Ee67ttNameDt1NM2891oaCQIJrsO70AE0OosMo+darpNvGIY7HitBMqor8lSZK4
MmhwtlsApjz0Y1F9lHPv/tmfk9w3Mlk235eE5CGP+1n/Btn4XcOdlFUV6RKsNdzVUU61luUGidMO
xfsGdDt2CCkcn9YmOjXJ2KwkgKDZrJId5WrxPXZXVafg1QtpWWqeYHDiZfJmcuUU6R0s2/j8MhCr
BHswcEoLo/k+uMzv/VkL0Dc18pt9TSdaFW3zainK6puJRULnQEsNy4A1Y9CcWPEp8l5KKBgCNCKy
ebWKbc3q7X2oMT6Qf1iUwL/k7NfSvLIWCvdP8Uk4CfSBUVFfcePk502cVmRrowYs13Abb7kC60Td
iO7b5f8HD6FfWaA+A6uglH76Trdhenm9LskBe4FLFMlYWhRedLscisecFm2PTcRqqA//y52iIkr/
6m0SsyKy/YD7ZD3mEYCryJtt8J9CPGmFafv6eddN9R00bBGnj7u1a+6sz6eGemLSwyZU1U+ul3Ve
sB8mX9QrZNx3UVTe/opAZ+PdevP6JoMKf3TdmwY/mtQYpObb+J7r/90P9TRQUMhWNdivuxJ08g9d
egiU3yMbofr8Xc8iIaIiLgNFfRGFK6Nl2F5rVqTGywpd/nE0KkZfshM7N5xohLZ40wPSy+Kp6Ti1
ecPJG30u5y9ECt/Q8EnB6dhzkOP4gAFHWoUNPwghmfCCGQaQJcnFIUNmn9kYwxzSYbW4SvfmLAlQ
uLyxY+92zxCJLJG22QvCwA5RnyNCfB60rhEHkRvsxT2wJgHVSXkN57FpaWz7AFDhtCcWfC2SbDgL
mQZUpJNrBHmJvGdTYOs0gHOd5PwiH2dKBEr7Sj0R+a77XFrP6G0ChI4eRckPgdzGolwJpurVY/08
RwfUf4M9L/me5MQzjlmeHDIMInTX9UaB/sRrgSK2IyxB+5l+7QNnW6NFTshYKkOzuSRu29P1vOxv
9bxzVTmBD8H0jRJK2t1QTQ84z7hMcHw6y9L5PT1bqUNDIn61yLsnXdrv+/sjApdP1Z2Qq3BlqC9o
oMNWAulJt4AxnPqbyfJE2jnF+pEQeovTr1g7XGUuziohXPd9P+d86GHI9iO85i4YJsrAUzrI6Lae
aXAhIQ2lkbj2qUp9rVPfQdzIwUMiBm6h0lQs29//BZURrqC5EYtsPEO7ztrZLBM0gb4Xr5GKKwZA
386d9hJnIxjZpS4S1HVnUU8fdgNhqmyfhIpyrzbfWybp8Vhkzf3GXCox+oqjEudZ6H9k7Cq301g5
shClEVqDlu60WSMChLqt4lwZsYlDEH/Q+Ib88QkllG1ZkTGPc8bz44mTvbWk2l0c0K5NlM9Y7Zpc
faJwurpCYTtEGHu05+05KZLRdEiRWGauxu6jT6jVnUNLyLU+szg2u3N/PEgCLfZdYpxC8txeqyjr
MD5xku3hZVaCWl+2vUyy21DzzTgaMyqRViZi9uSfWFKErgCdYuIGdwVATxBITXJRdOyWiUrtBKUp
KTMlBHF/BmMCUf94Ivhi9lveO9kRdIKAeLxrvUh4oZWeDzBQdYK6hBvxs7K7EDku/CVFgSwBHupD
3shiXRMU43Ez+/a9v1SbmDihpRqX20fGP8rV49bpkwRWfGuICH69OCghPPBu7kMjJE4Q2dP7incq
+Vbqv0YrSm+VHKmQfhd5q6UpOH8a8gXqoECJUq76JFbRWPn1DVLxDiQM1wFJ88TwGNAf91vn/k3I
TTtVwVmwDHJvJQwbGUNMbqUgPmwqsIuMUfitZdIrDU7eWVj4tqlxJiP0trl925xK3BLmFTiFqsFs
PLj+deULKobJMZ5Y1TdyWSx+/ZjYOgpXuCVXrAVnXNuJWqHmnIpSulneDO4gc+aUAn4xQw4W/pfX
yqOMLuCn9QGp0NKEZo6sOqHeLYKrSPMa54eNHNViLZJVBjhlW/0LYyacO1uAZvIR3UgRUmsUxA3e
tVRx1a2Zsrda31AQXZmx24BUaftJEbyFbuUgBfLjKhIb+cLhgCx86IXnGdq7kq/RMCtUhdsPmhKz
2t1cb2ma8bS1FK6EBLDSbXfcNZYAKqRunegHc8xfi3G8uJdCeMhbNNnOwCDxY7gQIJQgzeeZQ1nv
nNGUjduTX+dc41FyHq2e3DV5UACthQyh0/KEbGAVvH3UYsGtmhWo4QRMvJdqIjLO15H6wWV6+3uw
J6dd7dsv0OXNQDwWKYFCulyz7vOCYL3jFsumrv7D1b6MEoWC2vA5twE7xrgQiTYsyY9cFvsS/CsL
wlUwq++FylOXgThGJvOWrdbfGrXnwpZuEv+Qzehw0N1oa+qUftJ4syCZ21H6IgUJJqOMcg8VjJ3p
YGa+h+MLUtzYHTl493O1FgLgkjUQw28txWudEK3RYcrupOLgaNCTaDsoLl86FrG0MfJ7lImrxRZm
lSr0RiML+gnD027mILuCP/0UuDmTjgQkby7RLvyXbxseM+gqk5qAG+XzQCc4pnJPFUWCnSuU+VAK
sDIzBfeoNpA+z5dFKm6qd2c7GzZ1nbl0BSMe8AqjXOeH+peixW56Ca+ZK5eX2kl37JwVL2cwguzc
xDALFRqW0ztvu/QhKJpv3wJICAKeL+cZDaItasiq8dGVRagxz1AGYV3ekHo+GTB9bkqwC/dtTkGK
zb6cXaZF4e6ZEGbVuzfSTtD7NeSbLbuA/zQtE3mm3ABFL+VyLmhiD0guKQQ2yYQKDzgZJxde7NgG
wdIJvLzc4NedODZdTx4eKItxsE88WNyPv6Nx7LHDZ6+1tSHxO5csJP/Dht62/kyfsjsmlm3xgCRW
JrBmF9DOkI0LSq73LNKMMHyV1sENW012psOUwM4aNzQ59ByMMNcV/KgZuKXo0EMSga/aTB7svMMa
52RYQL+uJ9DVMvr0jLnceD/zRDJxmqOwcVogp89af2kSb3jZzlhsV7MVId5R7tRUoMcYPK6txm1I
iS++YL1NNHm5oLkoSbHi/p3LSEgBPqztE7Hdt8prYyJKdb/d+skHRWbUQRo6u81V04mSHUYq3J2B
H3xauGYhf9kW5VqefYyP3noVRcAOWYMKno43TDV7SxD/fMtIDMhi7/islvKS4NuzFOx+q/MlBLve
98r4HnQdHUwQCiNym9gEEa4VMPtV7l7EviF5uBrK2sZgv1Dz/o3ahJjYHXtQ5L05CsnsFUNUaxhr
Wdp1n5NKBPzycLdPfkJh/tfRV72WQEzSheRsqTPGgT1AfakwhDboUqmFDYymc2xUcIwo2eo5ghbA
9N0PAQGfjmnHQ4FNfV05bG/voQUUe1GOj4ACJCajngrt50B5kz5L4UIqfkx2DSC23ua+uvgBwNqq
06nnD64rDJ/yT6sDb/9RSrVVo20TF7i9zkNaplOWRvoN5amwaaBFNkHestlYN1s7nKLNclfMPFEl
E3cqJSw3+4wpRPck1BpOhpr7pMXpcPsC4YJdB0ssJOTmZcbwwT2tVjlQDP2dw9oTlsNYsNBUVFae
qiCk+7hrogvNPJc+TZS9npVXKj2kHTMgFwUi0smR7d3RJeEwS1gBsUvPbQh1io17u5U5LKnwUr35
QmKYVJqqVaH95jkbIKMN0dBOGtrRSdZW2bXI1cZ31EaxuSsUhr0evtRR6tu8JtfWiLxaDWBlKgO6
LwO6VKUjlU3FS7q0398+ZV4wqHRBYAZjOT6EBcwifZRIbSdYDinbIKh+7NKwssizPL31EgVn0Tkx
Rvz6bGzYvQPL5WhQsCYP+ROHLOy5xuv13ILMCWV3j2WfMQN3ISCl15i1ZWEjcuvQjBkllzl6YS5H
8plYTOqwLclc0TFgrxEjM2W66+Tdja0kENX50KhnrhaOBgU7OlYdNSb/t1IsN7LM7P+LqzQqpvr6
RIL4f+Fu898CWeaW71fvzIGHChics2xpZkkQ/y1qUZutnCbpg1CrEuVpb2Gcex+Al0XOAnOWe0jI
todX6+L/rx4ZH9SACiMvXC6H8MRxqaoxE5eoMNrCwirhhTpz/ZNAA3KDFxoP9OV0/xxgZ2rkY6BP
/xBsju6o2lFzQ7urJ7LaVyE8bsMjwk4Hhl21AyJ7MaORn1W7oOrgrzzMnZqcLPTlw5EdOiHWDosV
kK2Itjo+sLOf6E4UYkevZ5p92BODljZ3+HTDn3lc2vmYYF0cCmkcSEV994Pz034UkVS+H/z/yePc
37mMz1yyUauV7EO+RorMBUCD2Z4QdKZ00F6NYvBuZbvGVMp7yFRHKMOaHyrfKBwC04Te7xLyx/ck
Dtvwsp+ug076Txp+Reu7bE7Izb1h+ui7C4DglaoL4ozU5I9XyvGO+ixGDFfwcpUlg1nGdWlDRe/5
6BxaY3L58gFOJpB1fKvE3auYfwpRzZcAvCB5zlZhpGBmY+o2aOjmwYBTI/rTzL0/DNC2a9xpNrRW
V8LAbH91EwINk9VY7TBQMdjqGtgzj6q7Q2qYe2fRgUnQxMmWjot4gVgDtoI8BdKWzUOYGTAjyr/D
aaUx90vdfsWL82rzMGkjAiQQD6NTh5s0hgUfIiGTPHC/fy6kcZCXCNCIB/3rSDjZiQSQl5bIbW4/
qABYlpLiMm5GZmLgbNWcTyWmcd6553sG1ZHZOqG8Ay+3+dtgUfFAQ5CTz8/XTS2oRHb6QxY2LeFr
M48eZwJTJkNLrbWRkxhAaXQBCfhtMah7AaVCySS1429Oe4Da5CwnZIwxWdItowgxKVTh9et18B9v
9v5Q+pShTmdMsk/wjl5EHUAtrdt8BvCIBD6YZOvGjjYTJjutnLYYF4QGiNV/0VSPNEHRwGYEGrsl
hX4d+kKZGEDVK+S4jyMkn56DDuKaYHSl3l9JUWmP8Bb2SU7onb2Yxi/WtDYmMLabFeWcHYkUrUbZ
/Mj+RzyAWaOwHYOBpJlAKurjD1lno3azJwE3Ym2mrPi/+B4XbGc6KuhosB+OPOlJstmny6fK8W1z
YYhj8b+tmg+by6MrxT8nzFhXDY1oCs2RKhLFzCUE99ARzzEBLcdLVocFX7T34FApTI/G1jAzjAjb
eC76ajJG8mvKHg7nz4aXelgDb9NdeT2NFK2GNaukCkBzKDactWEWNYDdmg+TrUb7XcVtz+K+IRzI
PWJRxiqrBZ5Sx/9CK1Tbb+rrJ/B09fkHaNceZIkJukvCZoy1gF90+uWGk5SrqX5EGW5X8JkRCx/5
3Y7+qQ+2UGufKpGgZiI9QRfEeKvogBorPhfInp++xrXIYvqH+gzOvySqp+H0JXQ9LCevart0yhKO
3ogcHCO3nAysMDLO7fZl3qt90p19UH6mszarNKFPoWjmV1zoePtrcvLECvxRxhqGlKv4xXyZrFmh
zod3q5fuofZzPHaI9Q7YLAG+S3GX6eocoytTy4yT8KXIvUh/elVYCQm6v64nAqNM5q7SEA0eZQHg
Fk1G1wcN4/y7WNH9M4VdUT8W7jZkkqbKuBoaDBKXc8BsUbxT/Nt2lBKHYA5HNtP9ffafvLbwdn8g
BEGQiz6jj3lQWRBoZQh4e6rogs0d0z9N93OVihbHgggikN3qVKS44h4FWiCmyRDyv/JUVhIJVsx3
LsacjthUGh+3IOXJirSk9OsCXYyr2kKQ5SBPPt0DLuE/tdGHQUVBlvYg748K07pb2qxDmpzkON94
qIeMsKkWOPoI5zaB0yr/KobBIcLxRJNy5cHru4u4RZLLwDyTMHRcsxjm5D4cMCNfeG9od2SVJKrT
iUyakO9lqLhY6cD0NOgnRonTB6m5euNBq2o77DTt/dELNkSLBeMjLpZEZcsKZZe+gCU8ZM9agOeS
1BpRVwUKhLOwdm9/EZJ6Vu/sSdEcvrSggo/kNHhKI0Cnfl5UFyCORwxfUa2ZqgcX/s6YDPhxn7O+
db1IPWxEpZyAFJ8zbZOCDTYCdNZg/QmJ8rDS9zvhsmxHY4+FFGG67cF+jLwWQZX3lX4XHi7d9vdq
562eGY3Yey8QSGpnmGyie+Eb6iza8oaiHG+BL/onk4jOw+Z51eir2iqC1My/xgOkAs7aIkFAJ989
jvSavoW5pQLXHyUp1qSJgXRqAuXSiXEDnRO27mY9ranzYsPEkFtQffmDqHt6XvqDHF6ju926fCvj
hnzQ66Ttm8Yb/OGFVgX1QmBYAK7DYMpejqDRusRbuIFwEG5g/DQiCD7B8HkX19aJTDI9UERlXyv3
3VUalwPUWlyqMKuC+T1UL/mGu7nS/Qy4tTTMuFVFrAh4BOTv3MBiT1qCnE7D8yayXLMwKiLuDrJd
cyB2bTwE9YiAP8Gp4ShVjPLUsOtPwfFcVG9AMpBcokP67670t+cWS1F/uC1UKQdtq6tuWgCthAoX
/31yrvHIDRMiwDg4AFLWg78yehrfNL5h7+obY+OrZCwopkjaHia4rNQJfEV2CjdnRLz/TE4X4U40
AU+f18eZiOddnv2jVJpUgmHdxm/lcaGIswLmLhwD2gA7bKUbdEcr1JXXRQN6lnlhOwsIyjvIw/U4
ZuG5Ei8K9XeF7ahh6w8QjU48RjJxSwr9I++48CbQUbCnpSpAklNurptGY9srYt9ygRYbQdixP6hO
x9Rccl46Khr+uRAeaigrTjElBPemXq6pT8tqUtT7K13/PiHPY1709CHWjyrVBbpuWYxI1tVAPtuE
UA1d65GM3UBTKtdjwur3anZtJ7RkK9zsz3k+anhlwGWp91J5RGSYGPmFi/Pscnu2vzOO5vWcepWo
plgulbsM9u2VvosN4auqHH4E+NoTnB26d8l+cKLzA7t78yc3jTcvtzXnsjF4SDwD7kspVu7z6Fls
iRG9ZZ7LuSaoMAsJvsIGGJnSXWWhaFLcyzyN9hc52A2+f5Z7yJBpfMfCswhbye5ujghLKSGwlTeG
aG4H1KhkqBwAaYnXP1nyQt5Y74FkdfNTgJ60Lk+YjcXiUd0lLACuQcsRw7zqehWsQYlbeAm/n2Hq
eqvppQaz56j+YsUMNsKb5S951OPBgUyvXcDh0Goyu4Ar70jPOjy/8Ozk1GgYNBC5rhJe9nRBgxwq
vVHCfUlKaHteYDtNaxbVHWGJ5/IIUKmwFljrsFK1g6ytpaxai1JhHjufin5zQmHHHQFluQALdsCB
wHdW+yk4FOtHitFAeil8YelkUfrcMpcwC7R2iGdDW9sejt5JSVq3eu+l9rivEDzFEUeffRDB74Yc
kuirgWTMx0QY9ObNi3tSjI4FR7QSmIWeaQnIQ9Zf/w2GgZ845trnjS5LjOUxk3b6TY75u4a81TlY
9B90ZPdpRQHKgbvitEjEYQchiPrjrd4fNP6UGXVRvnpXGPHC7Isbo6oZPTofOWHkC5cu0IlOnT5A
L8SPnKTAibhCLZQsPNCqv7igsLfuznWAt0ttBd8KIBq48hdJwm7VFVbZrnJ3kBY3GmtO2i/pK7WA
ogKSHyfk3cUpwMkyDl2Z6sqo3zFt4N4WiCesgEVqz1g2G+3YdI5GRmaavXVgg19TykKfS1gWFeQq
GHKuIZEI6/oGbt+HQmMeJzjLsthJq0vgbe3pbhRm+REX2L5vmI8vxEqbjnJ5fHK3qexBxRJeUtQZ
Gv8wDuxLMnY2NB8NkyDy/YpO0oxrCakmQ/jZCru4cthpI2EJQlxUJGEGWH4WCWCwBgWvvBCqJiTu
1p+IUMD0fcBbfG79/LeulO9csp0/z0jFyoaVWaz1PlP/afVAQKQKfG/85mEFQPBc4ck3IZ3ni8m5
3FW1t2NSK0AR6HA3q44BoL3mYZUxE3M1CpZj8FaA0XCLTiZp4nE/Gvy9HLr3Po1YFCLRwa+gjztP
t9mwkOLKUmMmBnzG6kYazSz9Ev3m4uKK8UJLSiOsVkvMkcceH7mqfYhTrrWUhs9JlytrVYY65f1G
1HbZSJKjbHm8wSylW7Eu8UEqY1YEjdU5L6oA1ki+3R+UAjWNlqj7KGsY0jZwwh6b9eqvkBJnYG++
IAL1Wh7q2aG8Namybd1fd0nTDSWj1npWCOTvGTJoU/Z1MtdLKPpSlJklPBFiebfRcJ8M005wx16U
uuaR7iUJTqVu8rh8Y+n/faAa1A1upR6geU3L+2/cb715q+oyM7lNdXxPBCBLvxh3b8rgtWS+tHNq
wtBvJAjB4GDz49X6dIPUx0opwkBokzSnOrmxVuwhA1ADb5lmhgrq1kbybYNJDFqdd/XJPzMIHjGt
N5ix0gzZaYqASrQWJe5rg86uRoc6iWoKXTh6oJ8vKFcqdGwaMySoRXJHbx87Z6913KvJh9Zd5X1H
pfh7JTgQ5bkyxkdCptslrIDmpbi+qjxE5Qdgdlymh+shT7w45CuTLtIGIokr1+eA51uhucH7+wuu
hR9nULzpB0Y/OrtEdEp8k4o9XTenr6Gjrf4dEr2fFcaSG3KU91m2Rcbl0OTfgTbgNgnBeObiCg15
KPvTDcV1Gx/U1vRLBcNXUd92kXw6JP9VIehOd72FlNCu+EOuyjxqPIXhPnc+QxmzoPdAyLaEZIuB
NdDbdAKYSPzRGJLyWN6ujZaA+f2LMSXM7ufbQM7E2JOZZU5gFW+x0LGecVFNFvr1CYmvshS+cRr/
hJE+SJ4MloGxrwvfhMPW8Zc1Mi2PR7sGINYHP3Tt7YQCkrMwcte+vAjpjjE0cNPcWinRhv6wnaxO
wsN5FL0Zlpv9hUYpQ1JIliO5mFLZz+pPYhmzjT2ZU5jViswSqXj/OQXX6Zs7wa7ksiSqXm8hhIqp
qIwsSUtQAu9PlnK8Il8Gbe+fQjtt33pxR8AELze8iVvhQz6C8o2kEXuPU9Ww3bIm2qz8vFnriR+A
8JcwYWjHCY/Tbxij72axY+l2iZoAOhbcHAletlGWgBF6rBY8+NIhqRL86ZnGpWaqOvmty40KwyoZ
pBa7yAvM3cmFXaIUyfyAyaZ20HVguzwbnkamEKL/gnXTtmzvTOKdEEWI6lQ9yryZ3wnF9mCSUB7X
FBH5clBhF3Eko/Ot9xwawHB0Wq9yXdjZfERXHNEJjo7dAzppcGEprIDOJNH+7oL255VVJWHbRqbp
CrZzGxprj8+kZpixJGfn9ahQRRaoJaN5Un37qx2cOT2iJLduu0R1xnakxV64hjq9QcwT6ViYKbQ+
kJhfrrgpqfcwj6wxT3RSXY/rYMNhCAGJb+BxLG0XlnLi9OjngBd7x6FR5tTrVy5k6K6AzkqSqscl
K67hcLhOV50Z2PbigNRDPDetqpwFC22/gj7rfzkJHhQ8r8bNPR9sYe7ThKo1mTI7GG4tCjHYGQ/N
TiejnPBYGRu/UlnIIpiDuQ5KgIzRbLQbtG7m13/2NCoCczLqhuu7JLwCjNo6DkWMIW5IubXUvPHG
obCWu1zgeTgQLG88yA7aV7rbkmIEyPhbNZvYFaeXhPLOpSGvFsnBN2xV2psO30CecM06VE1GKi0U
/LK8LdGiOE1LcREWlT2oHG330rzBT7RG0lVjqmBbnTssGMpnvHzUSoFYUABPfhtxQjaYuffMu+r5
0GAudXFP8u5RTLB2dEBIgAhVIqWTxUNzQQSnSe8T4uu8MQV3g0j6h9hva2WOkSsKywf2nGM1GeW6
DHAq5GoyNnilDDkgImcbKF3+lP5B+ICozrLnrbTn7i/vDVGnikM85nB0EmUuXEiYa9syr4VQ9mQ4
Tiu075QmLqI5l3XdE024aOxNN1P7Sz43P/h9Yjuld4Kwi3/U/FaWQRd62ZAAhnxWe+153jIVW8du
y6oI2gsxZ144ny6BMMyPwwhLiLQsi4a8D6BtH0cYdYxkNigVJA54GZ7JIyEzoCAdII+LXm46nTvy
qF42G5zaXU8QB1lRJOt7QRRcNiDJFNqSX/BS/NYp1K+UQAVZdPjB7tkV3LuPbtotWakJEtb5njXh
8Yup6PQkiGqn8rOj774VYKQNHtfKGuMv54cWuBghEpoUyKzNA7cxGQVGzcp2TMUy0k8FMzGtiqdf
6S1S6oTJEpyurCKUQ0obG8yfR0oYTkG9LCdvoyOUAVgq+0Kzx/O6YVk9+uM3B0JWmPXevyHlo9l2
qTGT9Ql1SC+Xy8QShb4IbWdaa2OAxpiW8gfuE6NPA2D8noY85q/q11BhOFO0B+Ni39XQaa7xozBt
ugYTI9gDrZ6zbo2zVlsFusHfD6LGGN3r5SUYae7YEIHDT9IghZ8oFE/ruA7aKfaLheWuFxHD+voU
4cTgQSM13UPwfTYpKKIutvs17v5bAayXbNZQZOc2D2Q9iRik24EgVnBBNXEI5JyecNeJcz2xOr7R
7RTgjYp/Cq/PC2FqU5Ipg01P+GamO6o3gC88LJLVvq+KibC5O9ZjPmeW0mvMwLtPWa1vqMgPa92U
Nom3EvrOf8COsVVKd3a7JsKdXeRryeaeK3cju0vYuaAsVkGDRKAoH3dy9G29UHpWAO3OBC17hGpw
plAX9uXqUQzCr0muvPktmX56TSSgsQ6Tie2rB95LTxbfq+8aEoJPHH3Wi27E1pM7WXSoyuD+kq7l
ZMB91+b9LwyXBv6v9lG/vEVYeg5D/e9QFxewBJ4MhbxDPGB7AmiShsF8ga7Hc9tSmlaI59z42QHt
jWzHLLICAnShKYYq3gviv3X6Y4DOiy7cSqj/CenKcGqOxJe/4ituSmq57CdHkatlryb/t07aYEyq
Xn3ROSasTucehg/SGqCnDU5COuyc7st1D6wSsiP2eW3JvJssJArq31sXRaWv0SodTLjBC/pnl4Ao
o6TW3OKlwjRNVFDaB4deOGhEEVyidUcP7XA6xleXHp87wxX2voBikXE6rF5iZ2Z2K4IJhFnTvHvS
/mXo8mFzryUS6hnkP8dwepPxtl7Yw05l7LqXflcTnJaJ8J0u3Dm18U3RUFGs4IwBSYNrpQZRFSnv
cnrqgmGVqdxaDUSGH83ulwNex26d9ZvbrHDBiq9eFBrWSeRzVF48CquKrKkgxrkYerwvJV/pYRpH
CNMMpW1ssvwq+5DoIUVeTEPh+WgnTalKhP5S8B3mwKUGjV31oVVO9GTOVmiZ86sd+ufvVyaNbeq3
ONKv3GKwV6u5RABsX50BUBtikblrXaeu0fBuoaBIAWpIXwhezVG107Wdrzc/+RubnppiPVW4V1EG
S/0a4Yv+K1YCEyb1gQdTkNycXBdOptjzh6+G9iaXlcn0Wnc9bedtGlGtJGu+wJGuDx2a2mRKFMrn
OWRdQ2L7JeiEciYasOGn23vFGYHkkL/+Qr5srwN8br0wTNu2zh6dOD1MSv2gPUc206asOKw/b0d7
L/za4spax4gJSINMe4PpkWzV+IrDTc7GG/M5TcG6Puq5F9zYfePWvOmJpKfyz12irhLtsfXWFKU0
TE4b8YjI5kwx2qHrqfyOtglu0YkHPlSdVDQo0JOZZnz99d0yxfIvbSIYhAOYy1JpDLJhg10crpL+
dCEmzSlXvcxyKlfYolZIbL6xRZ5PBHrGPXxMzzhrh+7DHGMtxs+Bx3K+SMUbG7KnraQHFflrAWer
dLnzD39crwqBriiUBMM8RlpyFtCfvjlpBFnM4nPwEq5dk8CZPknCF32Rk45tuAcO+pEh7jB7EhaR
/hWFw2fd9fvORBOEAV3U/cvxZGgWTen2J2gWrk4Pm2JPWlQk+Zxk1h2o4VfZuPI+ft+Vh5xkXE7h
w5JvN9eF5w6SWfxVNzvx5qjthOLm2PlbnyGjxoFM5en0oS9WUKIfBSY0tp/qbXTMDmMKDA3UyEcf
mIJ07BaV/CBjFh6u8e6HEjs8xL3mtCrGvuZ/N55A4rDxsZXfCDJFeGiaKr88oadFbmsRrRgGWIxc
/vkpsOOLA+TqiJnzRmyTqf0vtC64EHb2cxvxeKKdU4cdt7zyMhUEvJTlhzLX13TEcw1VLrWj736Y
8zl5oggx/KA5C0LUPrkpkywIT2i1AXxD17JNepabVoWXCLbEJxFjDoJq0dWCFtdTedApfmlkvqRD
fkJwZXa/2y0QeNBHSgMVESX5Hq1kJ1j1PiCB6siYB3TrZT2lmQmkx/y0QZHlLuUtPVtzB0KPy3Lu
LuCEDankdquYL9pl28J5M/DmgaXZWcIJYul6eJH657xlA0zEzxKy+P4H2jvKao4NyS20tQbzUFgc
AUyUp8SHggS8gQmVkW3e7yURvtFFn2Pns9MdW14LqTjpAdTAp9kd7y+tvawxMJktiZdnX5q64mbW
V5WkkT3XRSwx1sCvtMRiRqBVw5lsxGT4cta63mIL7aJu9oG07VQK2CeZR26nrhWl/W1jn3OlI+yM
IGSrmHswbLW86zD1rmC9/cnqULg9o1Pfz0I4SrYg4IECYut95QDQdZYZbuz8ugBJwjEVchHh8cvb
xt2yDpx3HcKVv9BfDUGTItFydYHxodcimfxaqgx4peDwbOP8dvtcPpSYPfEHNxHGwRAfHRE7JGV7
SL/WEAcIMA3xu5LRgz7UDT2dB4e0/tD+aZ2LBG0alSGDImBHxr+/ZjGv1zADSm+AL+E8/3kF01Zc
nIzQHJWKgU3BRKsyOxSjKI/rbDnYLCXUCG9tKrwgfrAgvUuW8mdo+Ey1/jjzGfD2PhzuBd78W84C
Hh6EPU9lTBNDqPDWo0V8FqnaXXDBUfyWDtKIJWwTnzWgJOFuo0PUBlyu8c4X+ta/yMfuzWAvCMX2
zp2EaP9jYKBzuEVg7bH+voAFdJT/6BB973jnPaNDJUza8rcbgFMeKKbw/H+knx/9Jn1J3QavcuVf
AUZha0Z63IP0InVJTwcaiSWhJ6Y4fkJcvtBbsg+tMtxRW+q6GSA/+I0Ev62PGKWu4VDqf2OxHGJE
u4E6slSg4NpFOakPDxuT//3WEB+usfYr9wcCHN7m7i2bM9I2SzjyKIkSp5Swrnfse5EmqY7DQuA9
v5XY2IQq4OJ11ML+41J8oDwXjs+mv2rU71250qMzPETW/xP+dZPkecnq7Bo1qr7H9gmngyddBGmZ
C//s1xXDP7w3Fui7I6tWFqQl87CRE8KAgTHuzLP0RnecvZqI5qkWl8X9qavR+yPN7hQjy6/RZVyx
IxYmKvojPqp/7VMMT7IuZKkUKCto/bGVjmnz1NS1qjWHqpBcg7lR1nHu6YP3HIkCAXtSrFM73PpI
gKfwp2J+6CXymS2x2tQs6c7RFovvn93LmyJojEhkWLqDBOJgN841kFN+/rKbTCtwkSfs2ZxBiaDt
KBKm4Y8+Vt3Lj05c2Hcvouzl7DVY1sNaUuHPhLSq/ZHBaccMeMquf4AvFenHcpi2d88PaZJ6VWcY
yLX9aMHqmpvJ2BSW/XobtovIa+ylNCdYnSR9y7W97UU/zZz0c2BKRFc/pshnPj1hIBz8nN/5+7V6
7Tx6K6ZfOwmarMRpLp9pdi3qf82dCvFGsrqNlS0qiili7fWnhaRCCwl8iLwPGsC7F7ooFLASStLw
k69aVyFDyR7KVLze3EyvUDgxMQeOzUP2Kghb8Ltlfmz1lREmR1/cXm7sw4DOrTTLgHBdKRbACkFy
6iuspYM31+M2odgVbSizq4mH8GYkG+GsffSRxGuvX0ptXNllT3y6b8S55QDLAHP2sKJl3BSqhksk
FS9s6HZUBBjnVcLASXYmNLYzB5Vzxkgjo/MfFmIuVZukBFwExv2ckaeRBHbKnrVZV/2t3A75vMcO
6Ptzf4tWVK4dCytpJqf/ATPNoK6pOPvzBtDKrvu54lQqIfM3jDjnWP92XIUeAsKs/OL6rXmC7ES5
bUrQ5fgpr4yV862p+Y3hp9sFrLwUDzADghc64xYlP8NsYbvN8WkcJTKSwoub4fmRHjr0NSM7B2iS
45BtfC9hNNoxZOcC4XWy7WXUhruqMmUv52mJ8L1HyFfygHnJFAIzJD95Rn/dlyU2KsOElooGsVSG
noBwAtnB4F1GMiRRBpIBoiRJILTCbxT10e5YNpfME9FQaPsGUoBygKZeCs5ktoZxbbQl4taz+Z3u
q3o6eMRMbyVJZDlSXhvJ8QJV3xIDmbVMKE4EA4b2F7oc3EzDVUTFDXUeeFUC9bhyg5Gif1bUDLFD
8wQk4mbi4gl2DBYWcQFZ57nve95PB4ycRO5XDDn34AHrexO/mGhDzfscz9Z8Z/c4573sQ8ueX561
19oOAC46MBPGl2UDMKiRosJI+9ZqHTy3wj6jg19LlAoQRQcU25MF8tzfxPLPOabhFwh4QLdq5wQc
3gdvG+0wcTGlgVZa9Z05Dk+rSD1ZAHHWSLFQyMxggraNgyNsq6fg1ZnkFbyXGCZA7Vh6crG3iA2f
+gdc7Ut0spXIOVeEyN1HMYZb8sbzuNToSLvVz2w/tKsollR0f4vHDqNUdnmt1UDAxrL2N3lgHD5g
AyRVHe3XRRfLiNdVgjr4LGQNvaZb6v0a519XcqRqKMDKF1sfom6uMPZsg0SDoRP/kQKm5dC+Y/vA
ix10InvVTOMCsG7F2Xt3bxBO2FzIqO3VQ2hXJHFjJ9cueyUvFlazOjoPSWT9OBrE/iGqBECt44Hq
JM70fSoJFKLbs2/5bDsQK4+4EOss5Ad3Y9+p4NiJGdY+/lIhucYeQIjoNW+ZtFDx/y2ImvEBg9AU
e/Ma525dzhfIMmq610qpTAVCnQcG0vsuiQKZDtCDWPJv7XU6FiDs293LiKjDb9Yz3BRtFiTvrVf7
gN7DDqB41JCXAvJ59TsgYxyFKd4GrtC1RZ/OP3aSQsciv4GxgaKz0MKCMTzz9WjCKn1rEQWFQWNc
FeCz+SDaVT6SoLWuyz0knTHBfe8yaCNYBoDhjsBv0tjRGL5uc1cvdNSlTAztMsZIq6XcmL97/Qog
Yk7bBS9eUqyTvKnnT0oucztBILFNEPvBGrn07mNhzQct/myfNDbb8Wu5qyTYllz9tQhlNkOBE4D+
G7BY+0zCaNO/luioe+276gwsdffT0g3Y3ZCTEGzli6ObN56fKBvb+qpuJQUrJWaGVVdPT3d0iyFU
fKV3JzcWY/Kevf5XT3SExht0X9cuzf4yEW134+NuRtfa0pJ6SMP1+wq41R+FBnja9tqvR94ofy2q
idfc6lXvDXYUOKQtMq2EZsopsKlJS0yfE9eQzC+cT/tskV6YnG0t7SY5cK907idjRFUSpVsLJeOF
2+p6YSK34sHZz+8LaJI+FpH6U5vHXOpcFUiohzox7/zdi5r1MtbdW3DPc83nj8mwWDK9Ok/Lgru9
7wD9vQwOPNVosJ6nekLn5G9oy27n7/2NLQzf8KYOJGRYSSJuH43TjK81uraB8XhJq010xas0O1OQ
r0a0o6Zpb2bpCWFt3pzkJXh4brxsY3Urt6lkE3hhnYRGS2JRpXV3LcEAJQqSHs1xwJYDAJwIlpu9
8X8aaahEylKc+ic6zvLvK2l4XeyD5hJZGVXtf8TOKQYKaZ1l69Ppd1hI5iswOJaGlNjzQYJykwxd
CBsvonsGG+X6FVDkL+SLCxP8PF+VmcgVwJFzG+PfiUKU6BlMkNss3CPjleBdZ80MWTtOYQ0fm0ho
uN7JWWBxYDrokc6YSnHQ6GEjp+V9w8fuybiGj0LtZYVE04ZDb9fmH6M8VU092yQXyiv7wRGiGZdi
pd6F+Cf8xD3frmqsK92HcUGhG3zeJVGaXG6T2usOUkSxq5LeQWAUK5UTsvKEB9DhmmKeM1rdwjzy
BWPLqnj8PxU0KP9AL9LtzLh8KwCJ1NQZrKXjpfU6W6xBR9MXAr4dTAbegRs2lDud9qYwojT92akt
rh7uY0u8eZ97zgm5ZwbHxV3PGmodt7bmSvO39BdD51QIj0FejeQrJWMAAxVBRHr0Ma5lAU4praQT
pKkZaW0K3jYYpDpxePA0kMe2Y7yrhFX8vMOiUL16iSo99j5yiA0ESTAKv0jRxsEE4dH9CQpANoS2
UqohtO69uwFpiBvjdpu8n39A/R5V4uC+Juz3D/qYGxTy24maeWr+br8mVtABPY/trgUeVwc0JNPd
k208KxCnlnNjGQIFSoU/beFNvJb1dzKZ4s962/yIlnJ1b1GNCAB06Tvrr2ALnahuk+lisb1DO1bR
VaQDTfq5xBBknmBqqm1pNSA6vKyjeyAVjW55l3uwR43t9nq3M11+raZLUfE0VOrfXKHvV+PSga8j
jrdvTgf7J71gpqeoTf6BwzEoW2lBRG5BSZSiJsqZN0D/oGCVL7UODfEAF67irhW7nM5QQr2UcLxn
l5uc6wLPqRX5Ey2AcClthpQaIKLDhlYyj1L9qrEv36y6ITHepLplzYEDXP9qftpdN+jS2p+kVNjp
Ks7GQA1cR59PsJrZlbgi9aXSOvCh7hE1Tc8lfqVcYr6IyK+fOkfJOHICHDYhI/YgnGaSl3dt3KbP
Vznj5kMkcDRUVWCdyJgzWTDLT0pTNYIM1Dl2naTrV4t0v65JnKFWxzJhNRozdhsT0KAAJoCjgpUT
w6oJ3tBVohtHDs7gCQdMgNUbQ4K+B2Rd95FTXlgNxAWqaLgzuz7txg1o5ZeEPsjpa31rC3SYmP1l
YN0atLY/tw8bOWDtKFKlqXRRCmTZzvoNUc7MamR95/jDt3ELHL+zy99MSnOr4at7Igy4Q5ePg++R
MSYf50bfE+ayDLMyMycAJVlqD8cnou6VdpvyFdKKLlFP9v3frZNFexKH341iH1ItfxUxvIFaIp9q
yyTUlOPkLIWL+x8zx4A5QE8BLBcPWGpbBi66u6RVbVEGe0tp8jyqUTNgxpjSZnZXiAaOfc/IOmGg
fSfidFyzochkIkuYjUUJQ6SpQ0BPv/NAJgmk79kvki+AAhi/PfxbL8fe1IvvuRyHfjo+k1U4bSxm
9Zw3BKFAEplJDlmLB8yDsIhk29UA7PXTQ7evzc0MwM9zVAKk24n9VoLRHOUdQPq2y/eLxP2McdBd
82GOFJV27yiHDv5cJuMUHQlB02J1cr+e6rSuxVU+if71rKXGfcViMZQzShzw/iprUS1V5V1Uf/mZ
kTyBCwlk9+TvCX7XdCGnSj6HrnZncU++DYLWxDUKxiS8FEpUcDRNwQ90IiEb8tvpgnNuDXXzehjd
xUCRoGJEV6ipY5e/jihlRSf3lNgWQa4isFiHEYvqBWPH+DJmbsUXXNuNOz8SqtDM9Vjb9gO4B9Z3
nz1CBxhpZTUxQfETVT6IIoDluAeXoljElvxBKRicNsHBwrkrmEbvMaSGB8ONRMGRSxBu++R4PTY2
H+z6kboWp8RZPLedCTC0qlT7kCApBLyp5xOJAGbwA1+AJEeyEnRsCjDJJz1f2LfOf81r3DQ8ahiD
3vATqebRyFhXZGUDNk16KRx+MSlbrsT7LrxQ/x8MoKVJ+aNLtV24W6l/TCd0Za9vVzAmSkiUklY5
KvQWdOqRtyq+FkjsIhAFKxrb+PgWFUbL0yUK/w0js3po2ZW4VQL4rssEyubaFAoAhS+hokU3S0j1
QmKb7Xh1hieKfIMVFb1ojlTVmBKKXk0Lkcr/8hdbSHhMd/GIGILOhQg8OQ0CRPxt34cyNuptF3Ni
EMNSD5Rj9AnG7Wu9b8VbKCHNrOKtNPBTEx2piTyeTFVORgRXb/kzaXb0fD1qdVWJAxDtbt0Dcvhg
KHXzS9GhUsv17S345OUioVO/0oeFzMRIzk1gbXtbqt43KrGjFAqBvH0z6JbEtLPMyfxkBNDTHfCN
IVOFxxyKClIuKSKYViwLulkPq+MdG/mrdwBWDxmGorvhd7L6mepmYzVhHudEqP7TtAJnfWHIJsD5
+iZWmFtFSV8Ot2u6PZHam8WvLHo2/PBLrOyJZpS+jJBkzcArZz1tKiCrAxRdE2bK1+QHhaC0bTmP
qEWqzWuje6F4VLsZdr0EqN6+mw/TIxNLAVepBkarWq1kAj6sv9dHsebtvZBms5N4yFiqTJMrJm7i
yBNp+Kk3//ZwnY9opIcVPNY59SbQ4reurK8DJHseKlOZBQFrjVEg+esMMf2TGSVX0+aKdoyOyEeM
tmAy87y1wBkslmgUkIXOsOyUVJNROoWmO7PaKIju7TpausuKlLiMiEq0JHJJL/IvhL2KiMzXZSgk
Ug2PTCUA+qqUHXpU78AiMyEaRRAsJRj0a1IsbzAQC0EQBRRXOAuPy084IwqVYF39XkcdbMETURBC
Y2X6Kb0L89pMUaufUFPfFru8Dh+6FisoqIEGH1pBQnQmI5+OnfC+ob80lhl9xI1Nx3df1+wYDSCx
lrQj6oYMuXfRicw15UgJhM4qxU0M71R6vsgejydcxlbQn73kYYQuGutfuGKDeAxlwLDEj6obx0z5
LHRppjPfmovCZi+C+LBwUYZsL5maYj8PnEdP9i6S+TpA0GawLxlVETwPWP6QlUrOP9PBXGjiQT6S
ERTxusdvi6VkIXyov46MqD5Y5yfCu+qcKo63JCk5hXkkpTZkdtDEeLA8pLtug3MTA0dEpRMWyxvA
Wg7OFYviyX1qozc97BoAui5iHrP0To/cjDA/pOLBDc3z79AgPtSRaxAHhJlXqKepvj1jov3cvS+i
b5sO+Wk6FR6vw2xH5Rhc+fxAtqnySA7LOk6ZdkIMxm7zL9dCbmWi64i5O1hMhXt3BP+PYcoPK1qH
S5xi6Bmvghrozb7b4OJr4REiO+D8F2fOROgMdkiJCMp6lT8Nl2+deRh8qR0qCc546ynEh0jg0+oN
+uOXI0+v7SL+6Wp64irJa8Kss2XEk7YXZDIOn2KaiC81IatqdTNXFIs38LzI2zOBCaGdXVqcJurz
8fT04fNUwaUO5Vm1XFbOGM0xiDGMpehCpPHpBps+w4Ccmlcn1ubxGroFqSz/rYIoY5YfaNzc7x4U
+wDDUwQauc97aLwoIhS7lKHUQQu36hKl/3IESwNE9QX3c8dddd+0fSnRCrTy5YGrPxYDMGvKl5j5
qcU/qOGlrnvC/mOHlaKUCDsHGudu6ObrgN8Fn9uBVzGZKQ2WVZtGWt9u0vkKLIS+soDVvo19ObxA
ajuHAUhxkbHG8bmUqnboU5xku+AMvikfiVzzjvduDD5NJnNh5BgKkmEaD71mQBg42o/9Vmc7WSKn
HN4mf3hEZ91+M6U+tqz6mBP8odRXVnzph5M4k6L8tImvQNBYFnHyIf+4x5uU4Ox+3cMP3vA3YLYh
UaZwgyz5OhntAC+HLC1tbjp5Gd+Eivkn9dhLi/c1ug4TJN3eftvhz2htvrPsxJd6Nu0/WBYG7fKH
6cv2P+YHGDAicMX9CWtNhPebpnBkeLYhwr4dyzrnWDB0ZueYgW3FzFsKWU6Euls4XvnJZOEsnzT5
a+KSDZHnZOw5P1BToFMOSM1FCxe3qL/G9TpPwAKiEm9qnsVhxYJvDcMZnVTIpM2obBbNB8CJNj79
xI1o+xWFrIzLYVDDc+DmjDpVpBJzV7QM+YnUiptIYWiw2wGMyFVl1XxyA4GYCqXrl3yor5R+5tpJ
oI8YBU0rwgUa86MHgUKekXZI8oWmVLZjIyXHLfYuT2pBmLndtI+7/MgDN5HwMZgQznVfZHhauazT
ffFP/gdAjcyrPN165fqQaSt7P9V/evf9eD7Tpnw2Ndc9qkdSJKIQNjHb4PdFHhcsmcEG36BIP1oF
Dq37tVJUyXbL1KC8ENC7O5tyANPEtbIXGrlZcpvH8BeQYODU2LQOcqug/VW60SsAo0XA0nNxXQuI
36T78WWS2Xo/EgD98Jk/qi+IYh6eVVgbcMKJpELCeJ+YyCtqosDcP77a6lRx8T3cGUpUB2Sk+32B
vg4ZvuxtOjjMBk0zBNtQFXEkXoS6AuAmDj+LgMDQPH/9rHQ66lG9DzZYUg6tVA80xK0FQKLIh9mI
atNbFy9/UxE0y56oZA5Ky9KsRJjHfbZ5AwXR4Y2WLSPgZTUc803JAO+UZztm8EJmrW3SSxli+FXZ
w1CEqoUX4nx08Osq9CXJZSIGZeOe58qj38E52dNiHEEcXCUlZIsPyUpL4RhuxoPYf+Dw7+ApnOZV
iK40EPQqbdB7VvNmerLxIOMUt/Od6X9gll9xv9ZhciYtFnFSpXJz8wfPGcM/Nn5E8dYuEDbGNgS+
5Pui/xCVM7oP1RWeQxGOhSFJjmfQCkDRLQFUTyo0mXanLU/nVt1MWYoDdu6eB3TpVORgIy7+2PWr
mAQLH55/T7W87h4175M07IDeY1E5eMJHb6/cPwNs1tFHVA34EjYckKzR5RLHydOuFS8weO9GJBwZ
L8OOdvjofuQb+5Qk6wrsHVdjtU8WERwSwGdMSEojaAaaS6DDK2HtOcPMYYtEYKmCV5yoVg0j9dkV
6NA16quY9MkYKWwv8E9Y0+iU+Ck2BYxHdkzgSF4JajsC0AuoyseN0EDFRNuIErLd8P5p1scB4dYN
8jy56rYe3PgyauVkwzRAAeU8aPYMFqe9Ccr0wsP4GCTLhquUlnx22T88b7xVu24Aq4Re/o2Hyaqm
aylMJj6AgFXa/L2Y5a6SOw4nIH8a3Fu4xCHxTWZRnR3XYhz6eLObGyzPouTcXZBasFdQpGWQSa5e
Ghdk7o/lYhkpVQ3OfAdBIlUwIzJ6dj453OBDOqoUb0tU04n6/T2PDV25ofFBDuC6ucXoY101WnUK
u1VYnBhOcdPtuFLoJ6p7lR7xm9pMROKwlP8b9EtECsHGZRKy3J0JlX15tOsD8ZvMy7ap+lLFn22T
0CmX7tq/d7kYHtDXXsDsNgvpJ9k//z4vOq0nO1CTnLWqqD622hlz5EfZg5ccfeckA70FZcPMC40X
9KMtspJQfxjyVWO0iATu79F4LKNI4otl9bZwkySLXIMLfYaClVbGTyLt+cLLnfiDv9cfHnHdnFXj
LO2Reilinc4qVKIVzmAjzuq//Eb+HaQCwa8GaX0CnIUrcOK7oUznkqIa9OVm0A6oMbWSPh5FuTnd
hPX/pUAzVKNVK8QJYSPY/KetYb9qdkIEL6RzkxPNUwjhmqTaceMsz2U3vhmsDn4D2e9jd75493rd
LOUahU3+9NDS0FJpk9Al/aalCfTaCRpcFmVLbt2bel3XHrEwEzu4xHro8OY7glc87S2tD8sePtGo
rJ0PAz6EYQC8VPWFURCiwRv9gsQ57YwRrP7+JMkqPa8bGYrPfxKKdNMl0Pz2/xg059HJprsjte/r
I4zMpwldD1eAwInb86PXZBuKCzY3BCpXAKAj3CsTYgPwd1R1PtXy3T2NatcDEUi3dppgEdOKjOFz
qfCvSj1rjmuCwGH1YEXavnXan8/vKXR98rA2fgtzeBaiFwb3s0qU2KKE3uRNWVdt5ASecQDPWxq0
uSlKO0Pmt9xs0eZxDt4piK7DG5PoDdT2tiWaHlqL5RckcTmqUwU2pZpR7wdMqvGry3dGl8ygXfU2
N3ch4j4PF3nus3Se3JG94ZsgvJaoA2XHjTRM9ax3OMCYmUnrxZjDCpUmRRXf4qODAb3yqmh7C+Su
reNT7qNRV5IzR3hqgyU3jeCDAwOuyPcsUEIj10YaITgU2jNwGDDkqw9GehJXN5Poewtky0MiPhdA
zvsmHrfpcDGhyMovxX3b4BP1c4fl/yMd3pCiKmN/QMYPxrB7Uq1NZwmucmaqq4A5NpDBmLT26Zm9
5O8WSdIKIleMEFJf0SveEiz7/N4l0Yk3SNd+7CbkwtK9lrlRPnaaqKtJoBXgokDSVeYnRSdA+7Hg
/URQGKF4oxJZw8oOMupi9nlPtZ3bCmpYmtgHtCJ/wDdLATvI0Z9Sfs1s0Ihj50heNhDOD68J+SkK
rAkHL2PC90XZWgaJISuyHCKH9SuoxeIzdjsFQHBH7O+Qs1Be7EZQS1neMhZzT1dvZT7FR67x2aS4
+d0VWsDPtnIiwb/ztnR1mPYZ0HOg9jZUEDEHUkRvn/UFamnqrxO4TUxBxIJcEijBuqPqkLkdPF9t
YCI6aV2+L5dmGmBeeX70Qm4wVDwq6b+EIHJcdgJbK50qUOPQcLF53j+yv6wxKGY5XKNtUTgJcGMW
ZastZodpMtSdCdvWTdoO3zl09NaR/t/B0MVm1JWJSxYT4A1lML3TAYSjJB01hyxxfDrdeURT/bBY
vpIeRTCyxPqDffStAKCp9skfshT/l90JZuh4+ke3lfJNgVmc8Qn7LoliNu+zgb520oWj9CvNkGnA
iAPsCayOBJpB9IL16cVPMxXpjCtC7Q1Sn3FujUamzxwKH4aQ9waU0N1YiyoFMBSvG+0jb3yxFCSh
feTCE3tpI8ngnnx5zyNZmxp+kcg8uR/m2DDwiKWwhY7gAreFl7j+p9hjTGT2J9siE+ypcxn7+u6D
mBaeNomrdFVV2FUsP35tMLJZq07ZHYm8THzkpd9vFEb5RDOVkUTtT0YMS5XV7wp1LuFNjgT8MufQ
a2oQr9pMPNyqp3wL9PrTVaPZHM3BmFPw/S6272MvOp8dEAr9iZs7CXrY7KrlChftLR+g+AwC/uU+
3g0GGDZKNGL8eBnTbGp7Lqr/P6hKRJttIRKNseZMqxc/nJ+LaPCDSBhVYPeQ96WZEclbyKMktXjh
ka6WAgXv3cA7wcHd5b5lTNC22lqlBzTWWrO3DOLG20pxFSoRMJTO5fCauDU01TgAvuW9UnMdc1bu
MgDNO056CZ8fhVZBpwd0UaijX+oWKqEX7k/6JLouuXWK4rXj2KY1lXzpYDuHDyQhT9a+6uWJxw5z
Uu2ndlUR5B9Zvsbspx3mrxrMcQmvdpaLa4O4oSh1RS4WaBZwjkj8gNXvBHITvH9RypGs6xd2nE43
HQ9TkyjxdmEoaoBordKxKadZuA2WlK16AhWuo2v7O7CDFKeFuGhiKeG+gCw32dClNGJ2f7Rjv634
H8S/Huge0mNWpMGSkKHHyGnS4vt72xAc2c5RU9a66azBRaKj34QcPNbiflbsYsjY1tyn5UjbyGxt
ap7RaZEqafZzqcQtWndEBSnmzKzgA8/8V3AGw7PXOCuX7ZHzhsAIeRcn9vThdPPk4xoM/sNGvwO8
Cgq3iubP3GmQSofyYqIK/jcmkoNrnHiV9RrupO/4jzGr8EbSF1cNDTpjIRMhO1QkzbQRREPERiED
vZxADB6dKFO8Db4IpisMaAqc/XjxjogVoREjIHWhGqcBDHUsb5gnIcLLI9G5UEaU1SsDb9h1ZFuO
qoVLXeq7S6HyubpIxs5KOaVspzgUc6MyY7Sn8WMx/8zgm1D76DLQVJjlwzudlop9K1FpgwC6OMOM
a7aIfMATGCENsmNbWRas1kmbduGSKaI8N+KPaYn0KrEMIu31M1EpS3YjuQoAn1ARdRZbyAXVhv5h
/i7meDcIQ3zDt6UyBVUfoCgFMKcsahaDCy7lDBOqHCmC+ihQh5EXaSfQvtloxYF8fPYBD1FG5qBD
BcKxZrtNzmvmiWIPU8rkKFoPL/1RP87WLkD/Ls4ifBBFrqYDg9Y9lTRhgjGsUMVKgdTrkCoPgmee
9DRfNeLDjgwFwfT7KGbMGbf+cjtVSp31taHU3eWYKmaPN95K3G11PFb0KUm8RLaFRUz0qD8Tjdjn
Ilm30xPL/d9/A8xMqdvwTXTFdqolkK2Gx7H6j3ZXHvPqUxpgeqbsApz+SIa/8MS0QX+lB7vMdQhG
Bylq8aF220Zaxee/rJ+uo1T7IRQ23cbjBt+fypQD+jAAynTgxMwvLPo/vQ1FBvGgPsJx35lkSBa2
L10VW1J1O62e+TqUQVgyPE/Nto6yUSKlg353QudHsP++nJvM82Pf5lg3dcjhzlOphXigvzJkUWEQ
KJxzKKrFeyZHZaGG694U06pKhf0f54HSmyd1gfxpnpUQdPYys9IxHG/lNS/QQcSEQ/B5XUAaHHuz
TKJu4Fjw/iCU2BaGL3Uga0lY4jJB/dKP2IyExskajkBqC3WypU3ixsrOpiz5b8ekVRDyQ90elB1/
Cu0BoCeyQMCLwYIbTjLiOhHXT1T/XIgvF1zKsuQLjTK/Z1mlY1GmMvdyVdnEgAWW38XbztQPLDTT
zbjw+NR/pDTmrEHv6Xh/BDjpo0vz2snTf5kZbZyQY9pCnbmFvD3AM7fom2t4dG4kA+gGd9rrnSmP
vUcwE+xvqbK7fYaV1VwqDCb5b74VmmAKUlB3bTnxZoo8NRJQYBIHmD/7jIPMu5iD//0hsvDVBZBe
OHb9aFP4AOij6rdUJYmAzoO0rzi/Qa0ZGhuvcVkDmk27gn/R7KQaRoZ8uIzu9ne5QPj80zLne83p
1YE3y0OcatXwwvD3zJwEfSqMg1y0luqcY/kVOrLHPyaYcv72cN4/8nLwsr97IiP2vPgHBdzmWzeE
tsjpcQnELa5Nse42KRotpqUPFEs3w1IXN3dZUEaddYYndXFXOYm0DL+CimYYB1KF4816lrPmUfmK
GlUMBmxE55Nsk86AEHpMY9GPBsYz5JJpaVNlggYWQ20y1XYDZtJy7mr2PCVZcy5WyCEXnUFGmkOl
8y/g8+WMy1+leryWBeUw41Et47CJwHd4DAHqdiMoZl7nQ6MbtFkd8eu5FRPvExk48RQH7iLixVta
klQclrO9xeQqDvQTv13QTNRp7wAo0ayQ7z/EV1mrN9P5gBkzB/74v2ZaWdMdb00T3X/V8a/jGBGB
NPbQW6Z4QxzvUgpBGvpzXIXkV4mOC0JOX1bO4FWhP8EXgxxDBGQecNNSoYr3aE7uwkWfHZ5QML+X
VOOP5iEon6kV6le/6CMe5aLtEb0p4PGNNFG5j4roX8EAzBsSS5qOica9+QcDMU8Lonn9XakVpA/x
z3GxrEhufDrZ5FP5M/5Mx40rmRQ7XlzkYPHcdnfWbFqY2+Es87bBkhtspnl4pc8rYMhfYVtGK/Fq
z54ZeWvHhN3J0LhaMrEjJG4AdCA0Kc75/0wCC1cdxMe4FbJaci0R1JGciiCk9bZCeRRMqYoMFNGT
TiGEkCd9dgTsQlSXHVS/RU+D0wKiZEo7A49S9QrY4SlRc2A3fM/gwV7nxKPlxgYizwSibBoWdhVE
VDBgJML+LIlkjvS0OxvgyYmiMZFguRyxBo2IPAafalwx8QoRxifbj+VumqCITurZP6SkHGCUt6M9
kkhBCZMAGLAH3vkjVxuuJxr0hKrpdhJlnOOPVYSwacIdKviYki8ncOCpae64aLrynRIOdqe+NFaA
5VKcZy8ADpUn0uuMEoMi5tWu27ejJmp1al2MvcchvHdcZoq6kKV4Uauu8WXcKVEGyO/nMyMTx8bh
LWVUPVPMausn12l+W9LFkxxXZJPVdkdSF5Eqi3Kj6v4JInkrBMDuuioUGRNGIshI+//AoxcQdc4T
9dzsOmHeXxiRTtYtwXSYe4CyP4kMXM+WyqXm3aplk84ts3wHV5PvYJgX7ci3qQdv83aG0Wgk9Aqx
b9sdHp2NngVzzlus6iMldkI3k6Garj3Zn5HtjkBGK79qXJz4Y0NTDp99TRdHCwkfm9o4Lup56g7t
ov++fC6lweGwkcHknJb4pQlbpMyzCNEnZPXnpkqJMWEsUG21WpOox9bT4nJ8biXBy3O/GVf6j0of
ZarXkZlm+7qdQ1OgfrdaN2Juh8XolnMLgcXXEm0fg+eyDWd+hWni4/v1NE6ZzQXv3G30qIKDIIGd
OXejGfKBF85zyrKQtO9zq6DzZzU8EVYjCvPQdXgtRKYa5OBOR4wQOdTZy12lCTvU6LmGIWn0f9BB
v88cV128pBCMAxPh89eK4k/JCIp7L5FJ0NAfAZ2zg1ZgRx80PouzVlOKBtRuxYwJmPQFZ+jC7GPX
pGEX3QIx4EZSWmLZZ1MIMZFdNNE9NHZ2vncxyCHES6y5cG+Fmov2eGi1npm1X3ttU35tbdnjLaqV
vFDz0wX4MqVZZ2kNLY98bVKfespqkKbBGOeszIOpeSVC8SdsZsvHrtzvS1FMBtun1tmnP8Ow9xKi
bxHW9SYteWNJErrSdDe+EInfawJT21/Wu341SBqBil/2exvlbGjJTr1rdgJA1jrGYk6FG27GghYj
dQ5bb7K2XT+TjK9tnWv9EQgn2PSKpU5m6vhjTphPhoeu1owoyyrLcQpBKKeD574WbIcKHxLjcIoh
dHjvaoErgRHs8jXKf+0Q6J+DWny/J1pmohj3RhqG/aXBuO3S0AWBVfZdSxkC9YJYq7eel5lQsj3e
Bfq0tfLHk1LRdmhLiqKJeBrfqHngWM6aYnm6NesdC4O5cdyE/YKNUh3jwYFQOBvhA4Tlp/H6BXqr
0U795ZkvlnDsbtHzH/RbqnkF3S6JVhjM1E8eiEvINWdsYapPWlFrrHmFrWFEj710I2mm0O26On10
QRPiq3A0B8aGm1FhyGz5RLoGHASmz9IPTOMOLcnV+oM6L5nGESs0MVMbtWU/znSxH/wKpiWC5F+X
Zw4lmTaYEqSvUPG4dEeLD8exV43kVqkKhEFF4u8Y+zyoinlyVkFFN6sv0Kdztz+TvyMzQSM0Wu+x
/6f/eCEQvcccaChfu503vOF9nQ4KB0AaTAyupEo5zlgRM2HVX23GuhLx0+9hnpWKrQEvNeSLQWCW
WkO+KQWaRpv4jUwthwfrq1s8ttdItGv+kaHC7pBONLVFqogIuKMrVd5qMLa1F3fJWB/DoEihmFlm
nF+fbHhBedCdZnTRkd5gYuOWINU8oCBYY21hDma/rRj+EwLlcic8kEq09r2cC1mWMzTLtMnwB02f
HsR8Z/G8uo+d/jvsftkOAcKquzo1lYPBQgaP9tT9lQsCxZ59YYWqA03FM3eLyD3rnaRnjmxsD3jC
wJTTOh+H3llGisp22P00iV0H+eStuQLEPN+HZB2A/poP13bTijqrgL1gtq+eEMgGVPWbU/AFo6Be
CVAExLX6tGCcJGW2IqIHk3R1HxDkmg50i3CzpsUldQ/WayV7hLwTP6CdrBPS68abKrIA2Pi6ETui
ZpEaHvONr1nRuszUNNyZAJp94CSPU1oqVjHfbPZuAajrC3H25Q7cTMLCQzdyrbIy7vQB/ABDf6t9
H6YiXqAQWfjkqszgrxZxwW+XrQab+wF5Erj145ve6kq7Owt9i5m/q3Kvwtx+tozCgEzHvpiYft2k
gpIAMWZTbCq8Z1x0iY9tzu34F3fcf+pNfwNRPv2oBHPdbrfwv4LBVb7Qw2SdKJCo5bfH/pnJqF67
XplIh03vsen1xml+A/y99BC6v/gC9sHuWC0M2Y7xxOhoQDAwXbwbzJHHBJ1ysvlEPfHnaWbDLlCf
5uPzIpdfUPSHM1S8GYIuDcLnGWivY0m9swVnaAWl2eJUd3mQ7/VLSA+k64SM8Yon9qekPSLc/dxT
5ITAS7fFrddqVuXh0vl8vqGBM2QyMIyc8THjI0Dk80FgNqbbqxESM6iWjVHwbYu1p242HQtSEl9r
Jlid7NEoxaeBVbaU5uHrMKRaxwOXRPtsDcMTxOSXes62KrCG4ho3NDKZSBKjVjDZiUlQWvLhq6aa
RJBB1n1lvoxJj02pD+c3C1mwXh1b3TPZD+iEpMl65nQZxzpWUbLuPa1QdvUC9ar7Lh/OCYqe2AxM
wM6Fi3vxUVVT1keY3kyrT8t5UDtf/M0YgLp+jexIVctU/AWx3Ci+hgS5dvXv1S3JzK+9LJtlet1M
ZQ/4clut96KUxV/VkJyPC01g/kK2x/CpdjTHisWkUw/wewfIx83ux1J6gEhUTTpcHccxrmLRe4C3
YNlv2sGYjs6EjS9FiJK2MEEZqVjVBTcsB4BqKrYgiUoq8WwPqVSU7Ep3mVpmEX+c0X/cuGcTcAAg
4pKrGj8UrWwnoZuTi7536UDFe4az8Uz2uM5gwPeg8bqGjzpIV0twdzlGUisViYczgXMAJR2ddWYu
oJANBhpOW4FrGSRmsRFVFWpAnPvsraOJNWtqrF8mhS7x+iUEGtIBCvHRACokScnxSpZXub95jSQL
b1eOUevh1MTkd3sc5y6flHWd6pA9Ljy227dU/FrPMfymQo2sVYO4gE4PCzNzuWEBmkXL+JykLiGz
EGUrea1qCY85rNJjK+p/41W4tbQkexcqmzOwj4+hKtDyb/+PxjGc+Ahjihas9ts/OTtCXcf/uLfj
DLUqZlyDkzavAQdgRQ+lQz2DMO5HxWjeLtTvKrRSsWYfH6RedzhhU1fbs5TV6q42fzLS1B8oUbwy
fR+u9PqPJjlpqdSg4SFandJb5SgLozSGfHA0E+QCk6wMgA1SmwpJgokUbd1cyqj/QmBcSuXRW1hK
jkW1z8YSbOR7DNdlkHoeXthLDooyfzDNqRiiQvIYqMhNiUpydfIgeVl07DTHwgRR6ERbg6Hr+JUR
Zq1Xh4hpWnI/fMcGVtxourvnh9RPb/NUWaIfPESa0bjDHSzZdr+op8hst84kPfe2k5XJEMB7zwwK
nPxjRIyrPdkoaN/8GFNqeg5hCnFzChKKBTFI1FWKBkLKy+5RVAO+rh4WjPRQAcs7W70kMN6a9Wxv
T/tTVal5/9H6uQQUtzAwl6gc2/3TkeafumcI9gSuHJNpCwCPxCw+K8SY1Upt+0jU+qEl/GhgOWyJ
njJ64mU1rxTnTtI91U96osk/5DTYoQvJX8uURpWqqyXu2qkEf0c1LYbP+LuqXzf0GidqImmvyIDp
uPQU2ZpAkiVUvZanzIO+ZtHr2fu7/+0Kbhq1gZ7OX67Ryjm0yRHZ7voSINGPXvE0Pm5tTIY0k00/
t8Grw2QLi45+4d4LbEgMxoYIcFTJdC59A6Sd1S55Vi16kqIngjiwJUkgrBk650sSTmEOAszCTDZW
rJSA3DaFKzfEEnwCozIV07tDBvtPY8etuBhvHWKLQrf0Gv5HDzMiO0vC/yrquX8lgUz9ntq9YOs6
wC0XR/Y5YIaMFZY0KQ3MCXQnWDm/GKk8R1o8/yisVFcNYnADmQCcEFZ+DsO1KJXADE9ljeOV1YYI
90SYMkXfXaPe//JsaGMxuZczeGpUu2XOz1YlLJQp4UKPV8a9xe6HEa81YJ6rx3se+wLhN4VmgUfY
ipupDZIkzAmAm6Q6OCA4Pl0hDRwJBtgukwKLONrZiEL9uhMwMv36seaHJ6TYnV/HgF3Bllce+Fto
u8l7b4VMY9iv113mQQc6gEST+wFVWd4BFSSRONRIjtrH7Y8m6t3t+4VSFWh+RVPjIcAkjmAF+7PN
HwPtuAofzX05jQVr1jL6PGblIplzfNvXOeWHIdBzZRpVuM6pkbqnDRsQ09UKWSImH7tR4TbqesEg
93IQDsi8HtXv3X/wfzeBMk9x6W4WY1Tk07y/goUovgGXEjGqeb06eP/NtBg3/2TsEwjKhwumJRSB
a39PeOARezT5eBcpo3xcqCV88WTr7d4SB0WUaLdqu5m6giBLSAAbrLiHE8BNhJJjwwByJMf767ru
yGexbdwP4C5O/G3q7+WMI6G74OGceyGuFm1ZsHgqkMp8T81pxi/ylKo+1iDKkFx0vqjkkZzxMMdT
kQ2D/4ZauUqPMNPguQTjK1Jh9BmrYd3lTZB2mH3icsIi9FvGCbUQvI4RcRNNJTbGOxfIDdJwYKOE
nDFp8BqPvx9iE+WfvTsqKzlbFIiikTcwytvrtKbaTHeDKwv1E6mZp+hpKJEZwVniVYcx3kcUtHJN
7OsjudGtd+kkLUvOpFToeJrc94WCNg/k+y+4qmwMBPYjwCNah5KgYWGCctrAxm6cxuTDGSVbyDZ1
iM48SBHRRecWfQkZzwGYGi0GdyjkKdq6bc8BOMxG4Hu7rA/SDUxoZQX4h4WHwW7kH1BhC959Rq6r
KkxsAVZ3yhrg9a7JI2RWlJXlSsHv53d3wf6vUlIpk4ChTFn9pSp52vYwoUOzxH1DvUnThms2wPDY
05h0oEzFBOMUQQzqks6/jcM4TcitJsoAJgPJdF2GwLvc+qY3fu1wuxbZTTACoOytB5nExDS6xCBl
AH60rJd0xZOcm/vIeBzOah0GIFde437SSjSw1L5vTw59qxRGsJwLZsmdQhC+Tw27IMvag++MwBzN
3PJKqtC1WMjsXB8NZ1/O3ODPrJ3/mKNNyJXWWmmAO3fS4sg5rqOFKlEU1zGE675ZQkRF3aXwyKII
hJ9re9DdIrXQ1YVyGwLmtveSReG6MvzVIfahYVQuRcylmFWxky6yzQUcXi7qZ0vpPQGjkkfVY8bw
m3o3BbK5lwI+GXg4vxYEd1C7qGn/ubRfaqIbI+Lr9KdYo3BroJmnEleasDq3wcdRUJjXXBnj/Tr2
YnbB4Fi/DoBNzB8qVtbhCSSXBLd4D4YoENfqjU2Q1VuEgf6gxNbSnEwFErTAuLL+JO82BnxwOheh
3pOrANmIYvrgSqctaWMIBSOhVuaCPmYAGX/XlHmCAXgxyKI6JT949+rMe3NYdgMDG28IKNf8NvgM
gfauNzI02lQO8y5HshGvEpCDIll9jkNopCBY26H5Cvz5S+tuyK8rR+ZfuFBMmgshMclG6nALWoku
YtTfCsSvYJ7J//RQY9sz8elxzj5OuKZ3q6BbGOPb8fBu+JwBzNH/bhA2zw/1dvuzONG/VhfiqQva
Kh0njVDpOnZbQ+KrE8XqesbWSfYZW38LakT4R4bCO1awcfg2e/cDC0teVvgODSO89dPAC6MwnnEd
4nlXsv4ZIgeEVBp/5za5ATL3KWyjfPU3M7HiqNJPO05Phg+8Ymwy3bCuSUFy1n/Na8+9g7JCF9Ji
74DI2BCrr3ryYF8jMvW7iY5/4yR/hAI1JAWEDKIWCwcw8HdoXoqvdm9oArCCQWBYTBpfiBg23Q2Y
0sKV4Wm1TE4y/AHibIn1fxDStcLNG0UXulRAVnCp4scPgA/LFf7smd4vwXq0bG+miKC20evBnv76
O39FsqlvYj7SVIvq/oe/f+1q5Nl9Z5Ecjou13eMJHHA0O3rb+Ye123zkVJtozQvsUabR0QvyOtd3
juiUI5rma1wHxF++rX9M3FWq7BiKG3TebHle1vgnDy5baxSuuy5tjrcUdHBSNLEYk94/M5/rzGRY
bKGJN8oAxgQJEtTlk6613/xTFWjF7OpKTt7oeow+ZSMv52veB1G7Inh4VtFvyq0DT8sg9j0OwNbv
G7pKPgZf7Bp8u3S5drnlHcpG7zuCj4FQ/J1CmYsdD9GL9tBHw4+s46TdF534+YjJnOJcQNSE5TwH
89tQrjAIHnK/pJx78bXyp20QCuDMMsgZSD/IdTkAq2qNvJDIL1cIwnrRFHJgYaghjymlSL9Llqgo
tKt5k1B7LXCNjFABFgjNDgs5/P8YcCh96Ykc4R/IMn1ePR+rZM2vhHD31+bddAJCrlBzqVzc0P4A
L/16My595V0TCsshSvOxQDtvuW0Jr4xmNYEeXC/FIi7IGoO+GmKnJdiRem2vmClRhInYULdrHPrp
vs0rC1AbHEo1YLd8LU6AgKQLyrcKUln/ZodXXPz+Y1IP0oDYwPmmguIXmpRM8K5sxxRoyzSwvjtc
rX654trrE7KZU/j6lGIBPFCLF5LiVbJ4szN8q0r0S5cYKcTfBbvHEtAvhmc42pPyvDF+7ZanjFPi
tAjOqP6zLyyzpqijIkod4iz3f34v7vMS19a78SdyJk6hwr/7Q4jkJk3K6yUXx6B464yMxmUWie78
OYEA9+KWg26Qr9P/VSsPHLG4TahE7Al4zcYyX5Z43v6YvYuhZ7zQrDHjmtiYLqxVEM+ZmKQYINz9
XwqB8CHTxmKknXZyuAf+IGPKQDT0hazQOXcJLnc9a6MW5sLjVJWKMtJbONikacUhMpqyfbCniyFv
EIXUan6BCZ085f2xz7fOtRfKKdI4v/D7aH6kmWx4VbmopO9cyj4Xn4IZZo7H3dwjHuIOIXcFIMYb
ZvHkfJerkg8gsmn7rbWU2303ZkZQJwL91McQF09uTae4neDpjCe2rP/77OHzzeLEBRJTf5bNj3pa
EYvdd+UCn7rwEGjTmiZtbFpaH5ed8ILCqW24qA0tXLi2PWcuTsXVGyiWhImZ0SszePHcbr6AVRP0
JX5BAqMBKbUTx4sxk8PHPa/BMI45iZA/7Hhyf6ZjkxjWmoNqeaisz9OqL/olcvCJ8PmaeEaadrdG
8LBTAg2zI+ZIEIrPvOHNZX2LSQD10/J9REOaqiq0M7w0IgrJaCwCYrZLumswcssqMcekCw6+Duxs
efOPJqGAyxUdB+YgSK72l03aRVsqN+Pkh2cse/0CBaEuoZkeqaNLPwD7Q38KGwq41rfLE8i+zP6o
mCWxNRdsnEZPy0ZHrZ4SZk0wDSnxf8vup0uyUSQqoe+MNr0SBoQXDhGQItpNQd4w5Vkov+N9ihMt
Eje95mkKhcwBA3/OCgd3aZ/Pts6JKfFZP4r75QKef4q5ylhebEU1DP5dg5c+J3XGo9BqympW3dOb
xLujeBE6xXLwFAT0fChoLRSNjcLzddSxpkThYENTAUPau8ASDKYIsNQbSTmWfhCz2drXd233lsN3
FYunbS10FstaF3kCk/FV7UTPF/tVafn9AumgYxhej0VG8tydUkerr3tOMNj9xJN885b5tfAke4I6
+Da4UbZvfj6X/wI/mRv5kdTjHXVN5gLd9ezwx/QTx24rJvjao+zNI9ZHq3A+qkyKtN7DLd/ivD/c
lCaZ+GShBmDQwPJGiaFQnE+PJfR1wClHhtfzOwBsLb/0EIUlDbQ+MoM8O69vEWr20HZS3EPdK+wt
HoMpKRDFaQQV6SjGwvXj/r0M4jp+FbK4hNWVr1sexQUQ8/6HMOZsrpmTzHlQvBzIP4ZBPcGTiYIV
syFAHKWHfNbJCXj3XhF3bEDHX5GEA9JUlLCb3lNoj6Torl1JhOVj/+eVNT3toSD75qIsH5tGkBJH
K/7+AG1BZRKn2/Sg8Tz8U/4pkBR6aSZN8X3phvIo7odoR8MQ+n09Vl9ARywdujh6ZEw691zKFoqH
grWPVzkKf/a/oUV7THwzZDZ+jbaR1lYfE/PiWXzfmy7mKSe/V/IuF7S5D8WcqMzjxQSA55d4d+Ry
85PLHGWonKIO31NcEi2oWGtVWunixmKkUJn6eqH8Q3scYLdJ4YwC84Kh2Teepx8jKs5D4KPAH7qv
j3hirn78tdb7aGdsai8bDOVyrZCqxmtZim/u9vLPdW+cSySpXg3SoKMCHLliH0CySVPBzqkSTkOk
/oeDOwFof51TPYpTEE0+q4E+aYeVGU5CdbxV+AO57vqpcxsU/pF2SxAJKuEeCbaWX56DZ9K9l0rW
3xMHSoGtjkSf8gd/KdM0iDojQ+EQpj5DYBVM4xS62pV+4NltZAA8FaKCMo1WYbA96WrZxFoZiOgc
1f2UwU/3sXPn4Oo7D2JmRC4RWPPm5U1SgF5AgjY2be5fQ8czSVYfThEzw6v/Mq0m5e8TFsEWpJL7
Xoeeo4PwV1y4Sd6GfXa/LK1j9TC11SSxli+I0yg2cLpoTpBYNBOaKA2WhjJAoyAknmHCWpvaQT0L
oUzNOuKKM3wYWTlIQGV3nkDliHFMNZ5aPhO2SJhNu2Fko3gn6ju+Hsk+Hxhp6qOlUFagNtRM53XW
Mtmzn6U8yFSpZQIzJeAc9xYjWiM+HIpFqrD+c8MVR3fgqpvRJxDEyouAR56F4xr081S9LdH+lYdJ
CxsEaP/gUPXU6ZnSDL1/RXFX+LthN8OYYKChvbRenfTHhIWyqT4qC3PISjCKi85LBp5IUptDF7Ow
Q0zE6t80Y2YqUp4i1qSwStNu36YRsZeHBkG+XBq/bqjBHtYpkrezNHIg4kqD37FwU6ruiW3x67aS
vG9xu7NxrFEkDhpUEcfL/gRNBmuALULL/DtHKoO4cjMYPU2DffcxOOjuAgeCgPh/FIrMgUhxbm4q
j1s/fVE9TsbYKc2JaQn0lQ+jYTPeJSvcswhc7FLkR5uBGZ59c2rK6tKJPVWgw4uEF8m7FZeMm/2M
iBP/QLiMezhSUw8HiueTmCvLHMhLuxF9dMUAmkXvQSFwrx0JxOugSaa4R6EhfMDAJQHgL+o+bfQQ
zKY0xSZ+Ebq4nE4HolKtFAeDUn2etEQz3p+PW9Hxx/Du25gtxjssdEfrNckeor1DGym0Xe3EotET
g/xqVO65h3jBz+JEq66SehYgsMJEqqhp1ax2UMpWhS96ceb1k1VDYzFaMUK/PKNq4nJzMEbtSQH3
6C7a1Ji1AY6Zxj5ocO34chj9wS1kwfyqn5+genBVCWWrGWes4aDlkDKvKWVnbRH2v8wfKHvrYkUD
gv6gNInRS/6UHsBpTnMmyRLSNuruIvjEAX2uSeE3EoPYohVL+FEVEUVIzH4a3jTDwXVLstkExYvI
h69qKMcVvZcBy8p3b5SLUsX+oGOBh8DsfrDXhJBPlpJMXknZD1YFoahnd6VspV+EBCtoy/rxesAZ
/jX5ta0puBll3OVY4Q+yeO93xAQcsW1/3FY1XAaVKuPLS/2jkUcgko46uN6vIiiUI0VtTrVgdkia
V42NyQ2C5zvD/6DHJ4fSkutiMsxorb5MJUE9JJcyJpfYL3GGlhd7bZwRL7XMMJn88ISuKjf548PD
xVJKy7hgV7fX0sZdU3R7J1ESd92+QZc0t9HNRXdi7gVXhAyLgs4AD6T9NqdCezpx70CDesdwtzvB
VdN9avJDlmmVPxpt17LOvHe7BzYf96TeXzTDW9li7kSp2hQcZ5UyN5G3PnB/v2C2E2kZnUZofTVp
oHKibWDJOimcziTinqOPkcH3ZymBsxfCHaOsJBB9WW1zyx9odflDYEKsggXknDwsEyOD+nUR31Av
1RzF5N7TdkqbnIWO5FVXN+QXO/Bi8J5lduuTNM7AYE1Fh+X4CFRmmrnI2PCAMcZt2IFoM9jhw9Jz
5xrHijJ8ROsSoVATDuyaQy4jk+RXXgLZ42KX0QRRXcHj7PMTPYUT9wLpvavU0HaRQn5/wQf5aapR
eEVSqBFZK9WrZYqpJdeN91h2tejiDTVaXkw08GA258B0AqXsNisyicDy9UKxKQx2QnWGdlJdXgl+
MB1gjpoPAkVEiSCLPMqP/B2uemEk5oE9sqXWa5heoVsGcWThaASK9TPoo1Ul/bHH/fChwQ7j7A/2
xczP8Nx8LbWm76dtnEIU3Tcj2bhZSrHxNs4RDagV81F9tHUb6kZtafU+OlnI8B44yQVEA9yFBzKh
37X9EStZDqtGOjAtO04Ecihm/K2gwuN6UAJAlEy8rTF5ZiZRmox1XCvaarmQU49pdrwMoYK4YQCm
Kr+x+KYzvrZr4yeCYLvJh8cur7TOd1b89XR5oYSFb3iziGfXxO4HvjhSzOxpD8n4i8/c9VsWmbZr
52uWwM37HeMkMJ+fw7kNUBPvyeo3HHpZl3HBlz+HcHPYbTVEBsh68/qqYisqSlojDnYGpaBRiw+a
3dnim1bSvLZsOWG+lCXjwOEqC78mvo7Px+VEZwaAYd3mxaSHZtHcCHmd4WWZNuwBUkK78MYhBBw3
PI2SC3GbH8i7G5OYUXMkyrDCxcesGF4VS7wVff9nihAb3wMou+fnmNRpO4QpuRj/l54F5X3DJ5R3
7ZpMAVkiLlZkRpz73aD/p2A75ePrOqRi/meOQOXeV0LpUrBmtO6yILcSEausbd4xxxaHQSgvgFD2
TLXXjKUYezs3s1+Pc0l9LV4esdMY0T4PNGy+U9SisdjAVWBqK4eyscMImMy20KTbSXRBTgg/trf2
dpGSn6YTDWYmIbI3kKSjxMa94MkoGqFEyruIsUZ2g13hAEdKjp+vnkby+/m4VdMCROzVgJwXmSjW
HaZBcjqQb4e5SiqTlMsqf86SLj6zB1sa8ZGB0UiLKepBS+mAUpdWv2iwNADNyI3rxqKk4PuOxc4D
cmMRnrtvUy7MQ8/Zf1UHxLy3Q/ydGFyJd4ithKlYS1h3yBbeaWhqleESAGotpVxmw0C2aBxN1XR7
RfY5t795EtxIlQNNX9XnXT3tPF6X/Fs70GMjPrLFAFAG06Ld/YmPllEGbIE2erV4bUv2dS6I1DKs
DfCHMnD6d3Ws760Xb1neoQDrN9soVk+dcGYp959dx1nDqfQcTaRxlsqwnNxlxoaQREjuY1AlGZtw
s5PcoHwA45I+cQWXqv633v1rJwytC+mckOw20lZBhzg5qApZUV9LqvLbXWbpph4o5SXi48l6YAO/
QvoBarYaUOwNwAwIXg1D5TIGOzbQuWNzYmdy6iQcVOmWwWS/k9eTNYUVa2s3baM5rZmimGPzuCRB
+9AAyuNzEWNbqsIelw2jamps/ZJ0p4lGkn4S2p3dAP/rA9+1BIykHRPAYBRWZinvkt8Ec9/C0UVZ
sipeAq72Ai00FKO7JKIeLpyNnrZRK9L/IG9NaLJvl7VLJE+ZKC3u2aP4U4CxX4o1kMjbE7l9g/hm
+8c5T+7hVcriIFP7CNG8hXe0ur3x/Wrwd0pNFFnJlmcwb+FWrwWpwQZa2IhuvuWOBI+AdoHdcmM8
Sb8z+NHN4rUaz7kDYDDk3yGR/k4kI3Z/FzXoH9FoUlquRtWv/gg5OF2e5I97t94X7ixbbZ4B6eJC
uMOQXhvI5C622g+Usb93z3/7c36kMRIt55Mwt228gMixEfkoBtpubu02sCckmAZgdI2pvGoTCZYn
h/jYogYTaf79TPT0Bt9QMWL3hKxpbvxA15jbEZ5BB7qxhjQlzerKBMuoYMLZP1pnghDPxTWqc1ar
6pWtxC69icA+NrGAb/uQgscwKu5E0YwdL88cG+lzJYGAlcV6cBmm+qa1Ka+FnjsZT5Ql3uDNAh3P
8vMlR14it02OHY/++LccIX2HP6TjaHTrB9eiPNgSCbJtaD9qNMDCSHqpdW/Brk3Pvr9aFnw1Zubt
YmV9I2mFhZqbBWoWGhPyzSP0V9us7bD1Z6BCEdmoEu7poU3kw9FSwB2SVTqpJvFWzzTjMyobtWnP
0KH3Qfqv1K1Q5RFj082GUlFsGamJN2uU1f39G9ndtekoeTtRh5t2ZBUpcn0bec8OZg1Y0sUSgTHu
3/envwURK3g/nFV8hLLiHF10vlqBe9Q7DJZErz0qQhJqYQNMLHUXpdL+wiooKhSIPCA61qyqMhQr
8shJMvJtqddmefLjZNg++LsBhH2EvyBpVz4Auo8KxNg3lonEbtAv3l+AvtTY7LVPXyKwlHSbyk0B
vH7zA+dvp25zEpXxiVaUfx4SgpMahaXlKfP9N49zxloOeAwl7HWN1jzmKlt5b3ljzSDs446x8rBk
rYjG+mIcwH7thyPE9cuTqmVu5DDf0g6bCBaz4v5mEWA0MUFBvF+XNtz2N2gxm2vH0+ikseogqv5A
9XxPNslLkIVfAvkvN3GLWBt18BrFq7L4CSsHBtzPTCLB8Rn4lnKPd9Guv6S0e1i3zwvhLlF0xRcr
VTPQ1nk/uPL09mR540G/hNlne6zuD1wFwWINsaTn33k5pMGCwPa/BUx+3+p2KGe74bKuSGjwxXzl
HQtSF/ljcz0aIuhdIOcxl0l10G931FlQBjF3Ib/KvlwvbLzUwpEklgdSeg/w32p9Am5k6v5avo+u
mdUYgSwZPMhggsXKg+uC2h4z1F3aqG9Ns75D2PNYDe1ZJBvSwqt0G+jncQ4gPK1aTpEB69vCAl0N
Zomz1npruZdSUK33+2DDhE3/Lm18SkzyfwHBkv2OWPAPD1pa2rOXOvYNj0fQan/u356JO/rs7ptW
Ds6+DT3S9CdGhOaqXN3mURk8EjK7M4l/uYzoAUCbzAubzxKGUsIz94ti2wMBzWP1UwEfk46FJC7b
l6taDwEj77hQqP12K0pGU8TE8j/AMPvOM5hX9mAXrNsksYSNV+9viajjd6Buq79s/4eIw7QpGl/z
g+M7wIJMfVUEfjLXYlXMaCnDJ9T11vx2jDZ/dx3vYLEXICJwuIhz2WpHFuG3oHtH5VhDELwAdnAn
0bGARM3y1d9XjAinaFeIsTsFAnDTZAayISTemd5KGbci1rkTZmJIV3mlrs2qFbdaSfqxIzUtWmro
mMioXK2CZWMIU0mr2RQSY9j+7FXKta7a1HqGeRjzF8I/hVZoxuGkrKoHwB8Q7pOGXxxshjM1IQiu
VLtoSiXCIcGGMYBziaV2UA9lOJpwQCTPJaAkhZOUugDahbuQIg1SUSEl2WGX/vI3/4NaJlxkuJlR
tW3B3Bq06v3j8KIyATRacCxe4M4jdgOYtn+aM5OcsYaGv21DT7hWLfPaXzOYY6ohlb9lQmCcIX/h
d+ff/HTdCKWakHyGCQkYu4IZBn+BG8nxzeZfgZIvWhoN3UfWv96m3cQZP7MWkQTxDZy8IjEA9L/W
yu0+QNzj1CgQrPUfpG7u9bpIeXUNeey8nP2jrG1IGn3U/l7FPBF3aeOURxEZWWjDXOr629l3Crfc
LPukjltzM+pXz0Bnl0iRjS9izIOF8DzQnjLBzB9BLd1Q5oewQRbwpJ5ot6acXjYKq2b7zmFCNEua
iaL5C55QMyTRgT90s0smuj4BzjXxay3hzdL4RibfivdevDHQZA1vZTytefCpLru2sLZqt7iDt5eC
fF8mKKedWAvGpIzySO0osYrB5xmlL7zc66jLfOCDz26z81IzLH5OdY/VZsMrlDfegmlpxL1HddRW
RSkTfE6aet5aB53UBGTvbaXaEj3VJYIkDOmcTbWh4Y27lsvv2B/OqEgvmhvOaLxvILaPVMlZxIB2
qfoMTn64kIGgFHdWyilbAwru1Yp9lxXakpSRz4HcCd5UzQsnOun49+/rTZ55HDvCKgJqbtb1d87c
FJkiXISc+gGpgY5mBuSq/xuU4EUdwIXIWgu4qZAB48ELfKFaSfU+HfsPT0wPuSXrhIgXQmfKG+bO
D3CJEfl76sRAEinz6iwiV+0u7k0TvB1LNGJidU4V4vF1ooRvb6wyGsU759sUbyDEWH2p+RnuSK/c
baRlarE4WtUbsgp90V6YB5RBBq7e46NJFyeX6Lsdp8eDH9naonGKAMER/NKxuxGSOOxLTYPh/1Hw
hxQZh2YnAW7tkegM3+Vg37Nx/M+JeXowIKQs/OyuL54kNeeB+12pPnjds6J+T+a2Zrebu9WElNpz
LVBESsU2ENRiMwE+z1MJCqAWV9xAFZmUJ7KFfffVW/Cmf/rGZ6XdUFXsv+vAOj9TK2qF2BxzJQ4g
cb2xnLrL9qp0GPdsCh6fzbUp6xoLctrv7DNYzJd2UMS+ciOsJXvledn1dTxjkyuQzJUlyRoxPgAa
lpIquuUbwtBD/OI81MoEMa11MiiXGltCqjfUm2Ok/d4bl04x/5cUhCQoMn8ny+TPNCOntZ9IIc/g
j9/dC9FDzEIP5J/Fs5gv9yM0oVRaT1hvEIMwbj4u6+8FkAeVNA+Ys+ocGvEw5JN0Dqcsd/Ca+uhe
cKhbUe+Ox14F9tHx6N0SeDFgNQQ2wK6bGwubEoFHN0fl+47NWXW0T7ag5Jkh1yC/aw8A+rk85nre
nQuBHTrsaGo/EKoDTKMMzcn+6tRt4UHjcZn0dstnGAwnkjYuGzg4udSQUjdc53ZMLR+tz+14R9vc
gUyx5d+h0fo/HEWTXopPBEZd9Xw17dkOFOkOy5NBn+ulDLepbRffa7Ft/6+eGB9OmNLwCCnNU9R2
F+wU94TYBLL/AU9SR1Ome7N0JA2xlpj4gg6xJHEvRSSgmn2w0aaaU+vY7anbb6xiT+rSoICCUEpW
HOB0vJciQMMeTSsb/cGRdpnVyByeIUEdcMo4mmzZTUXdG2hA55RsZulHUTGKrqJzx21sSQ5BR1t1
7dIQX+xUWLI99xfb6jJM1rdYCoDf3E1KWQHUQMoXt6dzHLAhOypa84tjy2QVnNuGV21EsHooKp8Z
3qkBkbLIYt3tNN6DOQOdMnHFAUKMn3rDzl/SeS1AXj7M+OA4FWBUIIb+i6rQxQjIXGPguhq3m3UF
kJheJVB1FfnU38myn/I1kCTD817DWQeklhDAlgMdmgtEult0D3/Pmv8hmVQUC9SpzCORErXsmOz9
5+NqLYLpwS9Pl5UfTSFtz6a7uXhgMkb/Jr+FufsBgnh9uDuRiLOY0I2aVZq8YCZvdSF9H5XEVAGS
lm8dQuXDpIKfCJIb3bWhi8ElOtoS8sxt90sT8BmcKxETyCeWVcY/cb03kE9QoTDHb1ECcPeeT7At
HUaw0SQ4irohdjH9iIMDGSnCcZstmFtoOi90dB4IOGUwUmnjoXvLfmisGQUS6xoMZCbGSFqFZ6DD
uXrroeuCKqVRKv5SbkGt1RvLBafTS9gpIGethJoA7FTTmDl80CaK9+MbEZjnV+9Nc8h02Nigqd43
bbscQM1r8oPsSbyrVjAShzClnosa68mAKZa0q0so/wIVBc9dwfoVK5iOlqROmzESoHea8IzIhMlX
8H3m6u0GyEU3ZSj1eC+4ifUzHcnxZmHITZYj73yV+zprOoJK54H7O61f+5aojGqJGuSR9yX+MFzy
jHxDrvPhBKuQBXal1cP4cuxqizVOBipyOEGEJE1moq6dZJrGN7U/hLoJW+K2aECWAAf6sGS60qVj
UYXtrEzOyHVrlfzCcjLhf47I59T1jSNpmf311dHT5G60d1qKCE5pOJDDqIg4kDgdDtnofqrjUqP0
JDpLQO9mDBgKtgO5IEAp1jRQCdaP1v9A12sCbrIa4GKdLebwzFGlvijdwgOeuq2siyAEz/7QrDTW
FZpnkxp/WpsRoLIu+nSCySRPa+WfZNW6VUUUj6kse1+9hU/7g/HYXNqxExKJ+jbPhXHNi+W3W+hX
+nyhVbEWehzfMDGW7AMj4qPDUejheXq0Im5SYsUYelSyYX2PvXNHVtMrBnnTlN2yqOQqBfxgHThs
3gDxBIZAFeLd/l80nKSEuJuzkWxQnB9x3mMQLU/DotbQsiN5Hp8dzUmpxC76QzOATGxQ+mevwPKm
o7kjG8xrpyFCl4SJ9UiEj3ofJ68qdsXG6VqOay2rpuWahRRiLpDqs3p73UlwrNgoXTJVul+Rll7K
CqGt7UUCu1PAQo7hkwRzjEcPc01umH1wtSvAn10C0hezyjh2Um2Bobof22+ufmpvvR///w84V98a
W3FLF9bE9YWG4O3rJXBLWrvGl8tHa9Jw0qyYe9HQKqR471MfDn9BEgE7jDTFplWLAPCCBYx0x2Zi
q6y1mNRAZ+IAjaYP/QLRBD3O4zM8TrHHT4xwcMoQLbc0FqzVy9pXybJ5mc6yGkvxsNNY0ulGovin
ltLjgruJiueWTbtVcAGwXqucYIRTbupTiVImArPWA7AdZd66bjQBsK+rfDXoyEfxrBSsmUVGo0VW
cpBKMBIlTbfA3OUMeyF2aYQyvz/M2zvnEkD9Fcm9Po+kxDPcbGTngqTieSNZVN2gEjDNrF5y9Jk7
I+/z5FCmrdPCFi7rNk9k5Px1V4Yl3yXxhO8ly9mDPYvpL6g77/zbC8pSDppUxV91r3jlW65ekbCj
+QEPymqSftt2xr8BdmLz6dj0PvOl8czc1GKxEeTvkXa4qZroou/uTQAETjpu8rJN7NgcCJlv4hYY
YKrGSgHo39r8XNIuZJFNDkjhUU/skXL19YppqaBBbYPzKSCSAHHvtTCWxAAtd97RSq465+SbgpqH
LNcScvSD2q8LK8KRywrn36F0zmAmNJG46QVNaMxJetZko+z5guugaRnEE3PeM7oXwBHRb7IfurJW
zQ/9AgKPnWglbtu9vn9DBlo1L9VuUY+YNeC00zXcAcKQgngOWuX3tCk6aUjWHFMbkZ3NN31wirEt
Gfw7Ct5J2BtyAwyqaaE2WJJvqfV5FTCQU+GANIMv8SFTvIHUJ2aer3UHxCSShDFlY5KloeDreEb2
CnXimM4m2l0vND0sq12oHH4TeCZS0vSKPMJn3QCDScqReFVeTloyGN/Rvu69X3Zf1ZGN4t4S4/xo
VnY/FX3BPmWHeUaYCkgmqPxqtzBXUVsrLf2U5MziIb7Mr2f//PkVpLXIs3MSCIBlyofabKhkfQ3D
KK2HdS3cdiAKDy9tYvLgFSaDnNtwE8na15AVEeHmbVv5kKejRzHbjaOKYAQgcJ0rcDWeMAYcSLT0
hEJCeis4HLiSCX0B6bqPP6U/2JGzpovs3UwZC7bvNk2YhiUxWo991h2n0hPVq31JrfGsZZOg6Tlh
W0lujxhwnNMPnKdZFfWXj0yPhAEmFHIRTlDpHzFjU9MbWSQyNFqA1H5zWb9+HFgzi+DJzToenI3j
gR+EkZti+eQJc1vkI/Qiw7Lh92g/L7eES/gI0vkCegfPEic257mTrLhusONHLlM53bb5qjmwufeu
Mstn0jmuTXEjWJfbPc50oxyHN210FQIbXxO6PLQJmGJSU90CCpnHoTJXp0Cg0F7o9Rh8IJpcP7aM
gSFlO9xxvQnqPh0udP37x4V+mCs4Nq+woOHHfbG3UbwlATcgbkNavIdsrrgCRtqjdNXIaEkeV6VK
rBu+rC1hN2FwaAJAf5IXJH7kslMYXzpwPVEGmVygOHtJj9cMUVCd0sY0Fu+g7JOV9ZmgUNvG44yX
d8u5mjUKh8Ay+DTBa0Z9w0NXlpFfq6n/RtiftlaYKDgZjo8450VH3eOR+CcBj8g8svFbDwF9Zdl8
yjYnpz732u5mwRjjbhmq7zBVa850mu7/tmF0tQlyJQQ8SXKEkutERodSO2wWb0SdYpf/ZA/JaR0Z
4Lu1a9v2ngiGgSsV7CufuQtrmvdf5h+zax0dwRBF313U3s9w92Wb6/1d7Uh0ZYYGSF4vmxF4wlyR
HZ9sdelyJrmsmP8LZAy0aK+aF0sDrFAnD4vWottYiIX7Ezv+KPvMYvD6QArghLxErHsGo25wGCa5
yp8YMLLdCLosHorGFbrzIT6j253iWM9W8Bf4qstDoHFJxryODFKzNXjBxQDM+2lCQYCGuRe/0nV+
814f1hcI97Rr8T+4ouZAuM7McgRPHWT5nuQWYDOc8cxg97EfdtFw0Q3X0INxX3zuW+GZxDjKyMT/
U3afTA0vJIrv747bloxqmhrCVc3caNLezjAvUjqc3IO1kqDMcLQObgfFu/2zQs0OVoIC+d5a501h
f37mWkaCrhVc/RXtaJN+MmVLyyD8iCFE+32G0CgB1fu+inIj+XYI9Q8HOlD9eAHWdhnmw7i5uRbI
bMYW9l2TU/UkUHryOfpmcqmk7BwAZ2uwnOKqFlNaxxg2Am3xcj49DNWkRe4Da6nnru4Z9GhaeEUh
e2QZJL6o7QRWD9sm6gl60gfCR5s8FpxqHk/G24D7ZopqSY3BbV3cczXideZLE78nikEWWKKW53jH
9I6CklaTiBmoZl1/MCAR7VCbzmEn6UYKrFDHqG4FFeAAiwrmgxcJ9tZUIj4PhdM0DVuZo8+XZZiC
/ljevEk0T6xM8oGaPyBgQxOVXAdT+uC94irZjeTLu8ldbSUAyGoW7BCh9Zj2/IXyO1Gan2pNLELl
3AN0FgoZsz+MNs10gHeEs/VDoWaxaLSghV016xqJmRGI9PQIo+D8FAZbVNvXlGOb0+8DI2KNgeP+
YaLWGNY6MiP1l6cZrRe0cBrRY8I9XnqvVW74EARNQ9LZnu7cDOOE+OBacoo2aC1lf5GYrLMo867C
hEjAn219IGo8vOR9BNPPIKM/TZDkr7qGfUXYctaoJfIkCiIeJTXLduW/gy7XAocGITVYx1Axpb5g
6HghV3RHmu5y8oB70ORJBOH9aSqVySfAfF0KJ8wV3HEVDZa3CjNYrRwrYwpHLtQEkkFMEogseAJn
5Qo3UZpAQtkOjAXRASzIgn9FTmPGVcPjd2gUB4wRbJ1Kx8CI5oIuQ3JBjSxu6u0AHSOFWltEHPE5
942DJgQ2Dxe5FyXXlOtixpLaaGU74DtxRwcdUfMQolqXDnfNHKkSKGSaefF+fvA/URqi0YpYhqHP
6S57ZJh6CDsPPj2KTkhs+MPSDVvzQoE0ncehUOU8Gnn7hfcCJRoSkA6FlRLRGSmoJOwn8gXs/Grr
W8Q4Refdz4MrQz3pXvPrw47BcJR1On41up1ZxgkKpDE+7qll9LAtPcgdkGhD8kywDPyerevQP2mP
NukCM4U4MFwwL0rKaL1eu0glkNoiPQdGJIM9DniBzHa0rbBmc1dBEN2dW4MnLaI760AmPsQBw550
0Ew4nYvnvSkAMu6t29O3wSmK+HUCc4CQDFJv7MqZpJxGDNeZJqNK+LSI+RyOJcaZMGG24enZMAuv
PtSUWDPWrSr3E8wYH0Tx/9hRpUy1Kn3vDTxoUUHrPf2n+A6C3NVt7DpEiexSu1AQiiu+hbFcYY9Y
t3eMxojElcdI3DuQwgppABxBm9wQWjeDM/1HY6BFiMUavY41t9J7p0iXwJZ9iQN956rbcAiAio9U
Gd2WLtjX5UxDVTsBkuAE9kvKMWWZ9Zg629l28iTMVFVnkXgYh1aRk9nX+KVq1lNMDrfSZov7OI4m
z0NHu5wIG99qoqCSZToS1GaXK38hBazVGGUWoM4CNc5dmULylg1HV6cpLd6zqd1YOa+GBxFAQCNH
rQiZ5OhfGAHfjjCK6PTLv2yFq48JSLpFm7JDhzTqvCRxlIZNrGMKt5zK5Te8IpFK8IqwWuIh6zW/
N9DpOOVJY8tjv1+cEw38MSYSAQqhcH5PVy2S9IxCybK9Gi0OvC8sdnEfoUjW08XCV26qb+Dmh8ka
5+E34/6GSnZHGVasZfDpTMwCjtXwEV1yERtqAB4oS8TDQX6wZEhaiewZltElfwtM23+gNUIEb1rc
B1u0ypuVEvy0oy98lLyOLJS9wbyZnLe5GeraRAa3ojP408bT3n42RAtWYkshu5g6p1oPIKOjKvNv
6U1gbw7IXR6F546h+AoWwSQkUmLWooNV5usysByBTtzsYL1PvvOpJMvjNBeBO6d4IxYYTSZE0zPV
7joB60dlcE/YWeglmHVMFCAw9K/wUPfyEG4Zbb9l8e+VDfa24jc1RTwfYYWnYipfuXXIA1WEhpHJ
wspV6epgqGCFrmZC2L8A1n5CDFyqB6KbypGfn/83F/+DQVLwDhKHimPAvB7LEvclXuHXijRXZzcd
tx4iTwO33ryWLYQyrDdmG30y2aVyxCGjjt2//v7WFBM2SJReXB0My8fpGPdF+2zKDXoNd/YdzvrM
T657BJFXI5A8h9cnC0zdHV8cweIiUTJGYrdDdPcZaMSEAI+qtnRvXrFdXE85yYIMt6peg6pwmi0E
Ba+Y+FTgdGS0Osjux8vVekPe8MvmDxHW3IjmYq0t+lHQkaPOgLWKcUNCH0H3SRrLUuTeSCloxegN
TxGl5JbBs9m9WNooBuPE0GhBfJ05X1wxPg6ti6xONW08SMylu+VGEdXCDJq25q/RQbg63UVYlAu5
gyclVN0kThief0jTwFizo/Vw4L8YIRviROf6Ej5bXZNlKURbyA70XySpx0dmZFgECgIGaLAmsrj0
rX7uYjcn7OushfF8yvj4ft7SeglZwOZg7VbXTmjhrgKo2kCpQUNsn+zpnsF4fySpuLXePRcXLdUC
Berd5ZOaPdUy3/AUaRpGFORfyGlRhxjPoqDADSuvYw9CysU/PURurfoOV1ysDQHB0SHxrEGRy0ym
VOxN+INSw7tSwCvN5Yc9aXOdPYDjHy1k+JWa/gJ/vAeDTi9Nzi+WZUn+AwAkd9zAjmT2pibfr9oC
NDWhRdkWQ/GD60YZnoFUPu9bGMnjqx7vTQG+xfN3AJ6RVckj3HlJfgw/h/EFT7Y6q6/LHz2kvrYT
RyF1UQAdqttc3Fgy87YQQ30ppLo165hzcbQSFTYiNQSFy52Mbo3DXmIIsPtfBMi9LErkhpxycfKH
ZrL7c70juLpLseYwx0hyxVJazSGOPC2831vp/iAn/Z49GvljylvJ56GVpNqNG9aPrd0GXxL18HgH
0Y5U4ad/p+mCnW3C4N+RRX+srH7Ao1revOK/+m9M7ty1+zrTEuO9BQ08wpYXLxC1uPdFMXWXM1R5
mG2K/EcNNAFq3vt9vtK3QJYcKK1Zh8o9+sLV3skRD8XkFqVBYCct+798EPhbQgfOrJrjx1IL1LYd
oYK8TKwm2Xynlani//Ys6n6GBVbT/d8pOT+qCTI6mXegbr9sx0Ogk22acHET4ZUV33VyimyqIrz+
gM7ZpNrLuvPOhl6cEY++PIn3zF+gm3P2gNqkeB+w0ELtaM7tULH6FB7a6r6VLCTsVzgvBnaygR60
Pg+AfcGA5HIsrDa/YRig3G/Hmsnz3KOej69D17KxNiFPLMm+kPP/wuZr/miCOE0tJgVPu0OZn6vN
3xg/Ma0PilY/BuPF8o+o4+zebt6GGJeEj3Esw+3oHgKQfeICljQjzY5dZENnP/ttIU5hlNmzt1oS
UGt1oPw9DG/CfRP8HmY07qUUd9AmibQqw+vJ9nBbBxlp95lnZq6KiFNQoYCXntBN7kfcb5ZKrhRE
kTTrHEZ93RTSoDS+Q9iVneXoU2iAoYMX6tNDv+mvxsFulyTeqMTymLX8TnmI3rMR5gaR34z6FnTL
rWfjPf2PG8PPyCb3pBLmG6jSWczbUywRjOHnqmdAHnUiZbahcantzgD9TUXD1uLvBM0/0Fi5MbsA
lD79oQdyP1d4YKrYhbpiaDoXpNoOTXz3ODe3SGafi52d39pijVPdXkVDhHBSsPSGAXfqFkWOFPqd
cHukIwhgabL48IsP7kAzXMxHhslafnqgYJTwF9IwQflFIGSNlO67/ItpTcQvPtboX13xXZHHr3OH
tt5KFfadmLhBPQEzg/3AxSLndIBBM3098Jl63i91iW5fE17DzAUBz35bpuqudW/1T7gm+qePh1x2
LHz8C2N17+ndaO/tCwBpndRrx8KeYdOQJOoBSxVMbTNX9tLzAevTJgpJpPDINqIYBvPOIysobBGs
1hLNCKeDU9cNJvhCr8oOSVXrcRPzxlz2dJ+YCCFwnwnsZHzCYj95r+AUQwjoGlvrMV6eNkqj4CPj
3gZE6793OYTRIVB6u4nA9w08+bP1u/9k6fhviN+TUaqswQswRX+eoyJaUiJ3myG0F/lKVaobv+lh
tj3LkMxQoxUtJoa2hdKyG2ayMIRwAtFqkgqz9vOKqtznLS6B8bNXc5UM3rachrGr4cUMbj4Pp37O
vUd1qdDntNHywgdsffK5sXBU2IAiBG3RL6wR7oKSB1GbHr6k285FBm3bY7Wfrg4aX3+8AxnXDN4n
j6aTpa7/KAVI/AvF2Ufemr4mJ4ZXWY2bPaB7iG5zlZTvPPZq1aFBrTJjpuIuqowbAzJz6ctebjrF
XZGuLm+364qFN6x0Mrg9uAURCx4XVCUB8K2ricHcbHSd203Ne9H17SQr2NYrIXlu9PCcx6PTD9vO
NN8rIn0CnMbsgg/IbIUBBiqow3SrkHzNa+beEwzhOy6hpHmziXp73zDHHcGO4RQhUCQrrx9xKndk
nAUEANsRK1egJnFyQ/OAS0oPlATEEnzX3w+qRp659zcH4daieCwM4/wVELdLODmYdgJfQczhGP7q
PB0NKVqpOs1S8c8ceN8OCxxiesfVmq6tVGe0xXLd/C1LNFSEPtT4Yl7X8VJKav4OwN8CS7X82hfj
tLIpoWE/h94PTqJDPNARwhR8ZejL0VaD172vSUdpGYjA5g+EPJzwFrLgQf/mLTIwkde05u0GWM6O
R8XJ59NR81540qntGzU9xpOp7g1KwNvqItS+IWzou5IUmlQ0ekH3ekQfyaawgLBynRyfXACK2pGp
x+t80z3f5wf0WLcD49CsWWaHfQ8jnBWQ263LAaJlD28ilW2uxo6N0rx3K7vmFf0X0UQKtJB839z5
GqhnU82D5NbDyxD9brrC4plUpfEPhYImf9g3vHfPPn48+D3VBPmYg0kv5OIZN4shCT3eCRNOvDWF
leJkCokpT+uTfJHKauw/o5cKqC5eoOdmYzccl7fSXFikLTZASEz3uIe3v/XyQtUWXbQCGN6b8Aum
K79yzfJrG9fO4KBEZbG5srxR7ssam5jjAyZtOE73EqQlnzQGXlbrQrxHyHgPgyUqD5cAfniqciAl
p+ADLVjqiqJB+K76t3mWNW3ICfyTcitRRVih7wX6IiUL0GElUNNZ1qA2BxZZ1clefW+qjoWzOIUZ
dXcpxu0m3ciRXwayNOmixJGxa2/6h8LFWv5sxBpyskaFQB6Em5YFxollBRD1Uvz/4otoW+2VjOVf
DtuRlEvsVL24wJnmCfKloYDBduBQ+DBoNSsiNQvigdsLAzzkxTf2BEOyGywOHdAzZV5Wsclau/E3
6JUjaKOIjXrGe+QTBovA75razGICzrAvYEzu9eMtmtJF8jxkZaVlTQwUQHmznbzQJb6kSqRKFxbQ
tg/x1jkB/WsUPd6yTh7/QH9Iq3WM6qzXU4j0BBdY5WzT1u0EJs6LNjpv7aRTplIHSmlkgZw5iNCW
3vGrJusx+g/fMpNBjeqrjNBwPtBzFD2wUNNkRpLsd3Tu0ZBTH8/L2goYW48qvneTq1kN1KERHOL9
hdVNAGjxvwquZST/PMKfI6fx3JlvUTKbFlK3uIjC5e6RxRUO/zqTFrQ8DZdW2C2g9Kh3LZaaVaIs
GkW7wRtMZrD4ruswd1TgdUK4Ju76Jpyhb/0R4AUJXMcVUditlJr9QSJ3t77RKKwo/0XLZRALldK7
gQ2l3m26GJSAT6Qfhnaj2Jlv74vkgkaV7Sm5JqJg+UT6b6LSsL2guu7ydIUnjopPwMsMipywjcvS
Gx4yUx5BsiQ21ywXwU7GuIVOZ7BVWv5zQMKuOjJbGVITm+ujy/9LsyXdbjhip/30X4F8fJDXCZIj
NpNULYiKwxcTpAZ71f86sswYE39SUpawzFkC9aTYLqhdIinuLOZxsuZFKnehGNQKA0ZV7i1U2gWn
Vcm0MkVIcjoz0l47uRVsf7RKngefSQH+qsk2+/geU8Pho/oVSMZcOSJGpXCdOB7CRCjJbTTSQseA
AvmcMezh0wKPhSTHvHtY8Pl5LDfRcTr6KNDA7oR34pWoZa7nSKsJBuVyVDL10cMlTQvzG2cxc9lC
0ldv5/jzkjcDKKdjc7EUgjO3ONGfKvzHFp+2K/L7Zn6zT3+Fz6gqXsDadyStbJu/iip4/mBmZM9F
zht+gxLut4gErYB0xU92b2F/xWqIwHS8U3UXCYZhgidM4GHtfPLYthi5vrixnvpcSANFQBKSb5pQ
sDuJ918/Z4UGy9oyio9slT9glKvJ/z3lyCm8GVgPILQlPChma3FYQXgKJnyewTGzb+HSWmrChQyy
QeZ12sK+Woxc02BQt/p60DyQR2lD97S11jaT12L7dhnd3uiwzblmSnGvRqbWQWzHh2ap5IQfqTPN
AA/Z44h+mqp/G9giz8b6C5qC9Aroz0tcUWo25vLvS4Z+aS7AFhQ8T0YsxuA9HHRSNfRbq4ptO4ce
UIdT1uJBhUN9+FIhQzKEDKGCZQlEje/yYxSa26AO1RIQNRPlG6WzZCbG4uwEEkfnrtiF7RMBQuNX
QDpRgL1vNqjOpDJfyLaiKfCPV45v0IBmDfk/I7NUrIGEpmoTJ9OwmmZ8yFiKQO7RrDZViPbsXFGd
OE2HHJYR6iNT1qQ4MDcMnaV3cMoPoyhKiXE85/YUC4IIOyoZOpksJAFK3baJCzwxf5X73SyA8fOH
YWBSwS267lWSlYnqSICxmDffe66QMz0iBGZ3oj4GGkytP6wkLbDA+AdJm4JWFU/mgfeVxea+ytax
db7ueiBdQ1T3E3HsEeky17T0htnqBvrqE/i29X5oGV/k6evHJNTLkG1g855YXgh/Ggf3ym2mTopS
hRGbY05F304J2xnbCf1qF3roSzqqMt9mMkWSbNLLhT8OrcZIuP/n4Q9p1iqZymGH6jkG3CUbkMH4
//NrhTCOnRjKjRbim8Vp2/k5cQsPdNm0Y7EtUB2q2Wa0npGaMhWMaMOcJKBQcmmvtFD7rUg71ZxT
xFaMbtcLppJq+8inMOIxrFIigqs2hrxXRBg/xTJzMb0Il3N0YFUlrwY/3Vamj0rAXrqMzfiqR7CY
Ok+sAiA+FEGUdC9G/epIcNhuFU63qureOHRPVpzd4jtxt8eFHiij8GR1WydEUN3Vhx/4wShpbDD7
awTGSu3njrNdb91yjGouutP8hcnXD9EvtSHPgcEYbKTE72EkiLEqoqzWVNap4kIXg4q13BWGsgOm
Duj4aHPmpLi+zAce1zetpvptMcnX3osEwH2xeJAQJtCmtkvtdWMmjX0P8wOR9QJ1RFYB90yCFGw0
uYGfbI2ZSFZwP1ArcsGVS6W13TiVNVb636NeqTVhyVMXGYn1WuH5hlignzTnTjIebZCjqgypLuKW
VsG3Mdu6ZJc0/GWP1EIF+ZDL/aFAKVtUR4AHKQ4kYTWay3cU89kwXFhz3rb20jBhEURfqWbI4Frz
SPQwuyWCKxwTqPysLV2j0Bp0V1P0vFn7xlY/sg540zAfIl6Nnt0jrODDjmL0WWbCLG6VBK6zjeUK
S+4ie+TgYiFkuCPV7CfcLa53k5tm2gIlYSmU6UyaH6suyeHXsal5//SADf6E8CLnuKq6+iAPtCkp
LuMSyhIW48hSyhNgpm1daYWRED//D4TaD+QW1shPYqjw8Bxju5541IcNJ5N9Vn4o1tEWA7HhBfkS
QxynEku9th+/YO/CgtOwYpN7bKAlgya37PjCjcmxZHFWPyRprxpeNzsedzqv/XQYvfok5FSLoLQA
A8efLMQH5T+tvd7KkpM7XHv9yXJrmz0ostlNoe90+588DnMmLMZPbk8YzRF+bhLw58xFcgwlzKpr
HDXndWtqu4cE7hWns7Jhl+1Ca703LgtnXzIgVMVACcmPYsnG4BqfmUDHbkLF5Ah5mRsoiNDP6gHE
wgp0TIRrqOXpZiFmUJzw7rNvgzwNoskerOlxmH2sgGOGay0kQERWatt+lNkW4LRKcvHt4sWyXwEi
WJVY8EBqcjJyV/hrOJf7R4cip3YYkXdi+pDpK9Pl3vmecZRcT+zxGrypLh1jV9Op/J5BYXOOUeMQ
TNACbDHd09F2Ca+w1nPRU9kbRukb0eITKWZZl7YQNMBaggpqAJ+wWoQgkgBXWykSxTHE4Rd+VpCB
T4ncDtq8hmGQ5V9JeH9z5ASHoO0XvmvgyCDlcwipJsSsT1vPWYW8qPUyRRADWepl5THisM+TBRn9
PLhfMNnwpcWDnSJyz5toLV3zwsrgtkf1JpFmUDUz0H5RlQKCtPo0n++SjBZZH4K+uR0i5V3Co3ra
ibAwlVU3Ii7rMaFBtuup9biluQ4JVFe7rtzEbchUW0+21YCl1sN3EqXuIzv2IcBdXqqk2EXykco7
JvfYeKGuHocNqiJ194YrQLXgOkGA88HOShigDxFbBzFAb+jqdX3diNNoGc+8iFmgkJTUbREMAURU
lxQcAzhlq+xEt+5XQ2mA6o33B1BGZdbVnzXC02lxNtjY4mbTgxfcdmMntxBB4zKfBcOBP241D9B9
RmTdN0+RWU/0XOzfVdIwL/+g4Rq6bD/4sbzIXvuqAZd2wrjFgO/20DcAaF1pW/rNWfZBcAU7PGuS
BKWHA1jPqMoQmACRxpkrbXIHZGcwqpdh6j7+APzNH/+gEcYPvr43TFY2uwZBaieI00WFD2PGlczn
IxU3kxaHHotNkAMMLdPp/GnliXfej0KxoC8cOurqomCP96wDLqikuvkllpy2tzzz7ydRKaHGzi0v
ilFZOh6DObvzCz+AcRwPxA3dtnuqYqbZ5eZQJMmJS5JEXmYE4ugS5jbuuOhnB9tdv6hGwtS1ZUr6
Rd3L0dRGepiiFxqGNhvQRhvqkNH7KpDetVrlkj5PMcRuy8kA8k9CF9YNTDz27WSnNKq0m0PU1DAE
Fb+k9mymS0DEiYPoehC0zp/AOTo8P7ry7TXFNDZaTE49zLtI7PIjXhUl/XfF7MO4iiWvnNmaD+YM
XrIw4V6c2ZRuG9oZeOG1ObFvMarGq06PDBfgcM0N08iKpgackWFdwWxbBypZYJZecoYkBj/nWJt9
BopwrSrgUv5NxKl1ZlcvlvPNyowoBlni9NcZOlZ5sbgjhmBZoRsPaP+kEj64qQGV95MJ8u8GWDkb
HfXIzTBayRAV1J7ITMXne02LjuM6XojuAiT0ZBbPSgGO+ksKHGfF5yUxMCrPy/d5qUUWzcWg9nEW
PGhLNTqKhh2ykD0TEZCrSembCDcpFfDIgtXfvtuB+x6YIfu+0Y1U6JrfCEapNJpkjKz0mIN2tb7b
ceM9JHBrV3oApJnCDN3dW57Bg7ejjJ+iB7+MvAd+LXqM1bcH4G17WIGhklZ+Gujn8RiVUbrmUxGT
XAsTfxRD/LgAKRC5upCqrB4mw5dEnACF4Apvd9w2gmZnC+Xbyesw94P4NyD7Cq7hwFeu3YSl+t18
+fWSiK6Xrihl1EPaL/BYFvNVSHbjlEg6nsM25EIlAd7M1sH9RptvoP/wjoGz+c4Kgc2kCL7cQuHn
ram0U+3A67f/51dlWMvJTj6njQmvyAnErg+BjYtRwjlMqQFUiloVOVxqZwqVEaltP1ERooDQK2JP
JViJY3nmxesErDwPYYkSSvElebrcu0OszeWCzGOkfaokPPw2FWu5gnqHg2+dcJ1+CaaD9F8xPZwG
Hh+3sNcN6VQMIr40alTyNyTYpQZaS9KE35MbT/W0RGg0LgW9ashw+oOXXIurY7kzrXRJbrHP739K
j5J//i+1cm5MgnBeVuIe+nLY0TfwDJBDRpG4MMT0T2hQxsMH9zzIfMSckx5p8XjD+A8xzNkuDhM+
t54EIVkA1dHbLv0L0j2OKB0XhRR0VV3/xM4KPt8gXB+rsI/v+8QJ8B7jban5khz62Yp/50A7ORd6
vjwcfdPXbwmZzzb5XAG3WVL1PJ1nE6qfbDyaCQfCeCRPQVZ24D3Nx5/Q1cDOQR598ELFBQitd7VR
wotjSZRzlg84Ib0WddQXHC+k0rW5FUCyRdwprNKJxUoxXNSLNvtPTSyLEmOhthkFOyBmSp/bCD1Q
Se0wCPtKIfpWrEYdApD/bWMyIbIyVSKZ0pNsYr9otaPWeVPcIqGkmk2psrTUy7z4CpPsL1x2LHEZ
u0W02VUpUxWKnPY5pWVFuv/t971rx/jfleixXB5yYltmsLvXunZxXP6pRIE7kNm6F5YOx9wTrUsK
Obpys8DIXowTLDpc0IFPJ1pABMs80RUZXALFZQmE2WwsI2pHayKdklBgqf5UwBsYHBft0nFyBJjO
ep+CTel26ilLKZP/BoeSuK/8e7fSghfVr07jgJ7pmUIHdx7NpJYUYzC/KTexdeF60oJc5DzDwyA1
iTj6OalAQ1Uy528vcgrwLyrwzLG7Xh2jd04pyIhH3n6Ha3a0KmoTuqS85Yc8EDSpB5gOjxb2KQZL
YwWIm+EKBvpLR3dD4HH1pPITtAFUZzDxrh46gAwqLDRfiLiPdMWCU8BeDbj0Y1R8G3LpdEmqJJ7S
NgfujhBem6yOfSIymEIB/XjoNj+m0qrp4DzXrw+ZokplVAQZDxaz0+xKkoAOu11FoOHg7ZpwY8Vt
FeyRIxbRrsH8KhGLWPU9VyI/j/CR+C7NV8whxx6kuvRHsHF8rtu4g1d2T30UEB9jrWep/JFS2Biu
/IPjF2ktx9eoEiHwFBUHb/VbGWvpZ6WW1g5U8ss4g14Jl++EUGiq/y19QEW1LuRmNJejCY101aXF
YGnkFKY36LHty3FNJLp5FPUcDmZ0fYXvGZkWH8z7IShABT6dQ/CgCltV8u4m0ZJ+jmt1UpNDnBWc
MJaa8ZTNcI3MZ0tXxKevcbdbZ8n03l1IVktg3N4V2O/JMgkZw79TGaG3gn18uvcQeRi8f/N2XH1h
2Sh5+1vMWshOcgKxuqmGTDV5VQC7FGYmysRfqDEbuVNG66x0IY6rDETYNMEEDw1b+ic1GWgvKkWI
6Ft9m/AJ1KYWhpQPgy7h3kEWz+ncN8oHRmH+e/ECp1llqYwl7iBQVo+azpUjzkqiz3aU51Ji1CDP
/50Pi4t3oL3mBWJyrcJGC4ondiqHEnWvRrYjxz0wIehQbJKbQPbKLh3TZwoTc43LHMzFpq/Pv7IM
GG4mZ31I3ERd5tNycv3WKZqfqm8aFNvu/KeplPMmRPm2sZSWuakmPcmZSXFEHGRzibC78b0KxcSG
U2rJRcur01J4WET0/Pl+l2O/I8hL+KyDDcsvIYAf69fgz0HcKXCFctbAB2adWn8QN0uUWD4TYC6J
Vu0JBDoTtbvHLKVGYPhu87ovQIbF3Qn21zQZL9HeieDp1P1SEtEBL1D8C7sLhQYh9NWvsyr/b+DW
EJJ5dL1RzWpCzasUgyv9u1W7eHRJZ/ySDKUwSFEcqI1AQLVG0tatVNN4p9eUy2qLqiulLIJXwynU
11M1ce3vUGtsMg6BymOqs4C5FdBODRNjQwa/6yRm2St3jLdbEMqAvwluqBgffNSZ4dtaOfz70HAb
6mVxnZFph964ncoux91wludoouPWC2OOAJ+gspJDDm3JUWd9bHykDwiYYI+IDm6FJyVCXDofpGTh
1fjhEh0hJeq1lcY0OWGaWYr9bSr94wbmvjM6b6RnKDBXJ3TC3xdtzM72gihKqtYdvjN9d7EBazDR
d//69alyHex72nWe0RN9aWD6+lrkZ3Jgf3Wznqq6xdixTglqLMVj90NCCNjVLfThfSEHBnDmsTlo
alok24Vs6YvWL0QVbGkRHF9NEchgK+Gv6jjKa7arKVqmgcnfmqAMNI4bV8xCFsThfVThx6iovj6R
+6D32lDPuueewQtDG9VUb6TUBmnxb59nOUXHrGxaAHGRAT6RLMVXRhcHA591ZNbsfYHkcVmqQ+Aq
rlrBf9tCBEh6iy7qZAXrYFrRRPCX2JTaOAn+VBcgL8B4/9wlx4rEQ5e8L89ShTt5zwXl1+f+x/Z+
aszIP+wtC/GYi888BR7C+6rtc7Eqi55gS69OkOd7nJ8W2fJ1eF6bq+Ru9k8MasDOpGib3FXeBh7h
Yjbdexjwf41qaPb14ElKJE0/ybV8EaDHcTxduLHN5v9atXx2f4M/JTEfuO93HcdXXpR4fY1Z+Oly
uhqEqGbueTMEHjQf+TRUwxK4isv9hrd8wiK9AgYAX64g2fdRxJABbm8CG6bQgtt4zAoQrFtXKcjG
AF4LMjpHetC0TnWaLTon0uPG1XA5OQhH1r0krEA2ssNW7t6d3tSq07D9Km4hZjD3HUD6WE1vh4ON
I5xMdrvoH+OhERU8h5MtuvXIp1LbUhpcydmln/D8GrPzTQC/FyerRL2qHlVL4ObOrdPi692JUFQW
dfFDK0n3erthWo8OydP8pdxmmL1ISpWhgmdSWdT4rdV0yXMxo03sflC5Xv1JCNaSFTEDo8OAlVV8
gn5OyBQLxuyA3telKsybU4llawUA89ih9b5VnHnbbEh70gxO52rq9BLDVO6+Xy6DIDWnow9dXW/V
Kh49i/uQtnMGiAywcdexncI3SkswDoHxKLk7YG5vPd8QGCEoBUNuTNDhXlIfkj5MicOS+UpSVZ0g
dWeHvaOGrs8htkmIcIjHtNz1n3ZBTyKGzEyjxk+bRzB+a7XqYx+xVSplj98ZHv5Fg8t7APS7T3Uc
8/lAGMxU0KnS1qDZW6oIUOYLN2+K04afOO2vNIeRT1PM8AIwdaGT6dGXWJ7xcM/90402KiKLZPnj
PTb3Qv/S7Ozx/8Qyexr5Obt2zsBRecMquZglp4XjH7hCN4Yu7OIod9Jdvgyf4qZucDJhyziqShP+
ZR5yMcqlf2U5x3s1s6ZamFPEu8uxJtNCr8u1aM9iydH9zyd++EwANYPPnVTytpohOELq16cM8grD
8ed2wRsSd5+705kIwQpy9rghuYVTJpcFE9KMCpgNUNwk5NgEySibfc/tFoOpqanIaIy1boremLgj
JgBonQQ5405H8TDs9Zg5Y58hCgWV0VtAA+rGwRhVtJ5ALMrJ7KGNG+CZU1wWQhpUdTGCxHomt7px
Nij2L49fb6VHRJmJi4dA8j7N8yNptc6KJHHAvC4jhYG2HUHqzPzWDRNmMjfUsEmcpgLrnlM7jVfo
PKD0tx2UljpmE3uWr1VcK4lCXkGt0he3tlITzFae9YKFtQ1ydhiuEDdN6mFQs4jC4UpD5zii6KoO
EzQdMh2Sc0EduhrO2geJfqO3/23toXQinN6veZ8bKeWtzuiWoywDfV9wT+uUTLn/ybMx8T0Uc6Vo
lLk4P8VwkzomAE0uz7TTN8bf4C+Uf/8Dt1hhfDcNshBUasZDFI4gjiyAtbO1vqdXbPZQ1upw0oaW
gIWWI+WHKhR9LDtW8nhlpdq3q/dAFOYzRHp1D4h/hcKLqJICx6ZAT1dD3rBUILo6wXevX2TQmy2z
MyWhESri1SxFboTgyHx5KdFOzjSzXcy2SPmPCxN4LQQ9spbuZccA0XFng7ZSq21OXxbKLIbFKPYq
DuNXYYdBqK1IowzI+CCR66WvQYUbKsCwSJYdSusRwc7wzJrimWmDcc7qVnHSYROkUnTFxiDhqsrX
6JbELBy23Y8r5Dsfu4S3pgYc7B+hcskGFDu5ZgmaxFOk4wquD8G/3gZ+Zx0OoMljNBdV9OlL+uEa
87cnrt/7YdHZ1Nysq77DpEtww4HO7mEM92S1yDTvQalRwzT08/lHjQLrf5Th0tjNPCaCWKGT41u1
tXVvTPldzOE6JSPPxZaJq3MmF3SoaY2qnxxORv1FrQYKzvt+JTxrclpG/HPuGfJS6+J/2fWPQPF1
m+MrH7kBfypCLVxrPEKpqqBVoFCWGKBjehRheepv0g4sUZtYBBckO0vVXyrPP2zQ/8Q5h98l+Dic
gdLkUvR7dTaiFA2zgVlALK4dElb/1dPMhvEey8gEwnxs3muzK/yM78Xr/X+VycG1Bm3+Gzq46F81
C1BoZiCxt3czqoXBAP2ZQgXTBSJwWzxzCwZ/E830xL0j1ttwM6sZ2XG51feMpEL4bcVDCCBeUlmE
0hSEOFBKSAEfwsRebOVohE2PaoqVW9LU2Sts8KnzdmTVl4aEgF+wRNEbnaLDNA12dq1cK6a4EKrW
D/vq4DDufdwqWfgQIX4EmtWnXbSAdHtm9RvXk4r78ASTq+BWiEb51ZwcjIarpwCaFA7MGfHxEomB
W2TUqSgowSTUUDG+9/O4RWaUBmLfsycE41zEKrgbM12b7XMUIyA9u1UKc8jv8ZJkSbzUzsy6CqFd
z0D67nfT5pqkBJtT0gvRBjnK4WKk2kY3v2FbDICo8jyFEPJ0ZFS+m/t/sjLw0uzz8Sj5dvS0Zlhp
7GIAAJi7A5uDOkxTzQ8qZ1/5MZocF160b8OZZBjJeZcfvfHFnYABuA7tcicZWRXEW+obn2pdrclN
r7ZICKaSn3B8iBdytWoVAoO+phhNbAKd7S07MoRoRddXWpPiJhboxuMCWM2hialVUsEL5vQKaQm8
lr5FdUOzeeJimFptLflb16GmFd5jXbYDrxJe2TBxurbb07iT6mdcj/Qi5+e8F1fBJphEVu44K+lc
SLsOlkpaodGgi6ueCdO0/Oaqfgiwqpto0t7q46v8+ohAI/zp4XpJsh9m3DISr8TEwjFbbiE1CkrM
GUnyBEYEJoTp6IYV8pc0WShjiP18LMGQsAJdBlBdFf/ezHqVqb4ReSiNNR7uEUfaSKrBhnhkMzlb
R55XJBf5YffGuuXL+fJtmKf/D+lxSXv5J88n75Hb7Lr4LeErt5XO7jU1DIryGfC53QZHeVaW7IDy
xpauQGzFMLe29eW3tPgNGRjb32Y69DxlmOxOKam+5seDbIFHbqUi1KEa1l04fVpaRdPXKaZdvYoc
x9rmUizBZkVaqKeL7o18spqq1icE6MC3Ng8O790lQXQBQJInPsHGCYxmTuThIkrQNzUg8CcNTcde
wLWcVFlbuhDpKlGuUsq9uCDmFiawZE4eZxqeeEtp1tjzj1J/5PinmM2eM69YWA1rZaV9PJ1L8jjD
en74JtT4ikaEqFEeCKowZksKle5zVVEqSdSo9jcNMMn8ZC5Pxbc5tIE4WJ2IDZQXyDfuTyspxkmT
vIVQKfDg+121oplpkPmBbJ3jgP2Lm0bKu8qVtrqkyyQmkS9G7nhR2DrX11bNOXu/Xx+xGEUDMjfu
w3HF6RrbvX4oxQRVl6E5byOYnehjhAbqSNpWdJuMHn6pEji5GN+Juqeg/qucKvCYV3kggnAzbrVu
6rnARoDoK1TNSYfrdaPllBy/F4p2yu0EXdak1+ltmMCji+jsV2I9QLuH0pQnZq8ExWjkZzAVbj/w
IbiZb/qmEWqeBTWSUEKLiAVyNVjadWLProJ7MUsRQVFwc4R6kYdxBldr+SMdHb7ICgCueWmVl0Uy
zQn9t06+ev8VJYvxiq8U8qfKViT/uRiO+NymtGYYV9Zu907Yhwv5Avb5SquR1/oWabM209pf3AIk
k7NfXGQ8yUbYnfexORR07yJPywtO9rqehF564hftpksQPdPCOGO/Xl7mcmGanJgwZpP+YEB8i/do
wjPM4qx1Q5lpnvaVX2sjz/erL4MsJ6vIOsRthN5wh39OZxltUEAoI7wDexLkUZoacPBaHapoasxe
QKbPI6QJnsgW0WsyVjxFn33/f18N0jEvZE+KqMkrX8fw2ZT5kTozdR8J6yMvO/HRrm9zjcDDg4xU
q/WVQH7vnIE6X2+JpYL/uMLvGf0rFBMPcNVfsg9xDtg5d0+nrAMHoehDF7dqABieT1TRRAlhIhqd
HtvAQVUV1xowNYDZoyDeYHAViyz6ZT0UUDxXzdldC3ZBT2Yo/N3xeOs6YzutilWXejr8PE9YpAda
4TuAyi6iy4kVLYj+SWCmKiiskBaI4LAsI76b2G8+wj1NAQjshCGPjEjgRkJOuETO71ZT4Hufu4b2
k6M0LswEwuwFXe1CJnkVc6GM3nnIX2ThevPJ7gkxsnPKOMI170HdX8x8zXZxMNLVW9Xhz4Eito9U
WAzsMi/jWxmZecfx0njJn4qwCcaxElJAg0SHcXTu3JlgN0/GxxG643pWXpx+tPDwNE0GSChsz744
W2wEu3RfA/p4UubPN3JbkLHBt4u/qUd1TLXojaohKLjUCe7kqDT+CtCTn8Fu97gvq45PAJgstUqR
wvStShn3CLvbGD9ASD7XUL7zF2/prbLFd1ZAPtW3c4D9Rg6nWC3H+ZAm8LfMKKmwjMX43Lxi9o1Z
xUQBPSNxXFU3IjsdSm4mCT4L9180tuBgmUWonkKpzaxe5Kp2bJb+JYCEFSAvQBSCV2208M6xvHGt
QWSpZm2tgNfscNERW+84NuyR2Hi+o1CE33OKCsAWcwG/nYq7NFGcm+RnOoZgR7bZcm2aEzvC3qnl
j9oVCQTwkE6OAXdsAOM7Ld+tw1JafphYpTRIhS4i4CxT3zYcrIsrsQXlUYqVCUTe6+tgnJRwMUGd
5JJ4c0IGP1ANJpYr0EGctONGzN0qOJ1P9hO5uBYDYRcJ03YGcObE9TjBhLlS19CMAORlbKQis09F
e8GlZCY5ds4/uIWbPfGx1MivvEZ8F4BFy0gOiON1Ojh/CAVSTyhY7+XNlTMQEybmMLkZPyuaKnaY
FhZOVR/w2CJz2ZEua4ELswdzsKt+VlpoObjsb7fHQnnj/4g3rxkVvPCrgb2Jq2m1BPVuT/1+xPWL
w0doUVaVw8VqJXpDwRFXosnqB0RxplWvP2MqyQ6Wiq3uI/pN6t7TsKOTKl3HTHy5HHEbb5luQAcn
NB4plTdP3gW8g34EL5LJOIBoTkreGFKBqrKJ/DNP0y2gIIdPuqdwNaOTxA40ly45v/dc2xGwAYA2
VL6W0z2H7uPnaCltrx4NBw7o8dW4dhC87or/X5p5Zwj0FHDA/YAQHbbEWJ7dZTOmvSILZKw2QjUY
QO3gdvLRYUb0A2z/WsIJDLmqnk2oEsENSov3eh5UEy3eaV8cmhaUu4/EgwkggbI/HQFVOGzwv3sf
WhEB5Xq52eXtraCpeVL5AKUjYSPSKW0uLdL4b4I2Nmq/UhHQbRC2TZX5neBgxEscMma/AAwwvbs4
7ySb4vputnYp/ZO2cB3z+ACIjmoRBIz+ASst86nS8dojkiM1albK/HTTw1VrLdck/jjjQomBnlJO
GuGB6hBFkjVJwCUeXVYhP6kEo43VlHgFR0xHrBDcCv/A4nUqao8GG1xucPVLKor4Zm6nVXOfutbf
wSQ5LT3ukGTtonLRFuu1vlJSWn3nIYghSl3PejXYZ9a6uHdXJsxUVE2fEU4DUZuYZpyN3Lrn6Val
7oIZF5ZqUB0xzKShDVxeIoVOqO0gZEadAmOU/5VuLpmt/ggxkNScN+geAlhgoaEftCRoxGT7FCL5
YGjEN/RASCsaPFmo0GwWuERTGxIL+aky8iV9mqrIl0XBj4Sw2XOqHmtuUyGRT8Efq2Rd4UiErHyt
lL/kZN46iP0jGrW/OksOUbAxm5twA3fvGvYQxU+8X3eSbW+qyHS1GyCZi6ItL7LBV7/vJfPMW22S
oZCebZxAIXo/HYJl1Q9yo8bZm9f8d0VpH9RGT5KflgfI/dFs6JYirUbtZaVV12aSAlsTVqKolku7
fBvoC/vMa1rtobUDTcC2rJc1pRRRk5EBVWjeWnhVWIOh9BL/rpwGJFQBtoaUhIZmTYJyvGl9PoB5
furpRpiFagcy/vvHTObqECdWQzy/+6N+zfo6R0XXJJgTPtJVI3zb/tHeg2hQJXTwURuAjCiruFHC
bHbHhhVUBlWBsHC9opDXoxG2406KNZl+rw5t5jiruutGu5QDJyIaQ9YITbdVNjkxBtF+LCtMtkM9
joTOEGMhFsdcmz3KyeSeE8KL+PwJX9rhBuwQMcfn+cCXtOKU69nj5e9xmojzIY/TaI6KIN51Fsc/
uofl1y/WBGNNnCN6pagZhbv3Sw4H4NnPH7j/xjIRJVCar2wiOTJF8QCQ4mteoNNNf+/rhHoK67Ky
mUdi4Mx3TDv/8/Y5jA2YuBcp0BQm3keUhNmw6mTGNdJCgzpN0sjq62WS+0oAME4TDmE5SswxdfTA
Cjgoblj23Y4q79bZWVu4oeSKzb+pLOy6gEqTQMagcF7ZwCAgHEkUnp2c8ogf0XwGkilcNIfUper7
FALwLg+HdJPASrai8H6k6n3JSml/EiYRELgufn/KFTm0lGisYewob1j9Qkuue3oSJCoBWmTmZE/k
Kuz6X47ntHV4RBiXLRrtTJwB/3PevwOARRIXF4qO5aMbNqrB6X5r/UBlD+U/JpoQM0RXCtSH8jjc
m/BAmSyiNFZhcu464L4/nQKp2t3SmSJHm40RLmELyD9U2g7IWREPS3QKUXGP77J02SyaO6dxBAs6
d0xWbRM9a6lWxyiy8HnSYLZKSPDgiac45Y292zr9cqdbQpOqy8VTyCZehk4C+BKC5Ol3rSrrF1aC
zzfFk0JCAqNVwJsUrPMUibR7B2nparL8j3XgTUEa4wqRfaFUy7PEGNKsMGjqNCOdjPCFin4kRDP8
+nX1GYptvEyLNIpXGXQadf2JY60hUMfkQDgjiLrc/sHQYqMUTEETfV6Kt5WW3YIvP9nD84yt2YjQ
6QhlFyMmgaIwKrLvsBxQsPre8zub/8nSc2RQkxPU80u2s7HT1NcF+xMFhfKlKOjSQeBN7U5zVOYB
b3ulq7uoroTG+UX45nDdYqAiv2XT9L0g4KjxtbZ569F3Uy5BJT70hZvlE8u65IaMNgWakZDXOMEk
WtdQER75x/PWXxTRjxCBSNe5CpxEHZZaeT9039jp/QYw3B678PHo5ckmx1b7F4O7wdD8dLUsNgaa
ds0FtBk9stFP4ZbsRZTVN70eAsTc6+eENPi3H8X7cYBQvJ73+vHkcU0M8fq6f2lYuzzFdbShVK6r
k0XE1ddmcJlC5SJirKVcMPIOsP5KuldJ3YtAMKqeW6vlNCC2bxkv0koYB87Bzg7fuilIupsJJRx9
lVX7nbNd0QIOMrKBtrOEVih7JIUKwOfkQVCdwGBCVb4SQyk2xSTKw5KraXP6fTkHZQdiYShUhXyB
JYlpLAzQcSf/QomvtfazhWlQiIJFKqWnCu3A2+Ax1I0fMwM9wEdfmGbZQVKMi020j73N4J0ONsED
ddZu9thN3t3f0NPrGiKEKbvmCRiJKXTd0CPthEQ5gv+golRT/XQLC3rtBtkfZyfMfh4Hj2CmkjtI
7bgUmVfFqv/4+5h+d4Uo1sBy+V5KtAxHcXPrRdhvspI69VuvOwIXHemjMytRcUbnEQYk8ZSE+bQp
Da8PLBwyMh1KPXHhUsnrwMuH7+krxciJR1PKJLP8nIUbYGkxQEqG2zvoqeEtTS9CKBYqpHGyCSWy
pz9CbRrHymQk85dzqdvitNspfJmZxYwOMaNN8CnCD+DkhbMvjJShCfgaPCW9xWPyrhd9q1ZfGfrD
fVTfFUIlvFpvSAzaS2ATh4oDmDV0p1K1jRLG1rroNQMJUkURgcUbonNJ8KwprIgslmuiMkA4d7uP
Cc8QWW1Y5lDHYzJmBxYUyNj7g+yhJXX4Tj6HNObrpCYS7CqVixjKGSqQDdrIMxhk6P84vRvUDT8k
HdZrJu95czCPR4h4VsmSqsvSB4L/Wu8BR8GZmOax5QMrJLaoMgvse4y9evN3MrQDAYWgzNiAHdTN
+4cB4yt2kwsicehNAj5E78fxpMu+MTiN7aT1xPHkqBwVt5Harwz5ZN/xuCtQhPFE/wm/5uULQ0JO
wV6izvrpJediLy7kD6QYA10aCO6LYdae+3yjEgkEPb26gz0+9TvQrZkWAxMsyow0jlD9w7ZrjFYH
nfZXx18mxqrwo8r5jDsG9qr2GiHRmaw1/MantWZIXG6TGv0ECvKh/5g4RhQqefJ1LJT/mYsqT3ZB
ISpKfGwkUMOKZQJN2FPi0ibmKw4jYpr/W0PatuKlPym0XlU7t8M2NtLmJVF5yCMUGjwkyRddQLme
Cz0C2evvbSyAfrOGknNvJfiB/vVW1L9KG7EMivL051qIU4rDoMJVz8BXu35RpprdKj+4eNJbsUzm
htqHy77kEOSStENl+iCy7a1zmSRrL7EBnCi/QBIQLGuN/TgtnQiIe5EPIsCzfYaUDMzYvBMqY8xH
gjIn4cN3UoEa8vIlSqqxKTjP3R/N5ZcC854G+ucwAlVYCKCCgQ+XoYo/UkdC+T/nnwsKYe0PGjJp
SAsVDmvVmphyRNVtttcJlR9WW2/eAbxT5jwN37zHIx9hFUteEAd7sAF/P7wuwPliOqnoJJzWUuYZ
7CCuYwBQjoX/1OYNGiiKn+4i4onqNMU1o+2M9dMwcyR3xw9flm83VtrQs4HBAjNpz8L6vc/y+NcA
2Brhhb4SkLIuLC+MYP9wJDWr/BC2EHMmHaiPUgq3WsfxKz2A0PQoZMvDTiQiTb2+Ey99w4JrP0jY
MMitqKmUBXQNHX9ZJZq72PkGCXisQQfnvBdga1U60YPk0iy4/2mE0/rTk4a+ehrLQ2oAILjBDtZ9
CRf2/wQrAZX6yYHR38dAVxNTBZscVBJkh9gc46Te/n/mGgqsEUi1B+kJCbm9lfYOz0NTVvYlB7Z8
eR1sjkyjKHdX1HkvZovLu7PkB8giO8hxr6BG4efQsr1y5p/rVdVYj5MATTj1A2WI39nkbgiXYhhm
Vt522Tyv1dKB2QqcVc/fbRLnWzHodB/Iv3m+Cbq32sMS1F2Hg0b/eM/9ZjCVZ89dbN5PZW6fLZam
cQq+HjqF1CQj597nf2eXuhhbUMZvTmfeTg6mCv0+QbFr/2lU//5PDf/PkSaSC0mQa+wYxs7SdZ32
TWxyjg/6QsOJECbk7NEG1jdzTXTnrf5nGvixR5kNQSgN128FGeNXJM1L6a39pUVygllEo4UbxTtc
MZcf6Gakp4J5cZJPfDxFUNVeZCmAn3emMPsghAqCp9s13x39G5x4239Ao/4uWdPLuOQPyfSw3RDp
mmMMhOLiSW6Z/kCi4HKHvO1a6kbwEQqYh5o4HBoLY45amz5TZeAXA/+hwZQl8uv4mUtAzfhj+w6v
J7tjLL+nBiy+tE+rk16SdnrjnZ9Z6xPwkPWyzlCQTNIpT3Nit7pDy0XJFMVL5GFUYgPJRuzxcoza
uVGBQzLjAAzfMMqMFt4VGU4Q9sdKJA7opgRADYHBRoT6Ai5fs04SF9wDBLiDhhycMNPoW4MXXDIs
io8z0aj3v2qbkLwfPehFZdY1jd2hYbdrEIQhhoaWMP/LrkWVWCZe+xASA9kGT/ztD9suRf6luRrm
6lq8Rj3ktUwajn0cssuygeEKIL0F0idDs06CrzMOwNAaHEkGwoWFaATtBD3Ayn2PeyA987nfZbwb
EvZ/w1bOoogvlsSKzPhQdWQGSP6qSc0aei+WfJi3p7puTtdDlFgvy7MhpGkP9bH/8M3WA344XLAa
Cs2W3GeilllQL7fIqH2YHByvz9ByWj4rbJPAjQvZcwgyQHsiONnD4LFcT9kCrbKByooQj/nvfZtY
52mEAPQ7uKqZERzRHKogPfNDB/rDRjeJd5nXsPYpwz6NzzCCU1EoFuRNkCdHoF9rIXlilJmp3+nW
qSeR7UcmGjk0vsIL6jL0nKjSb2qe0SAtyvMHcIsH4ROaUB7EadID8N1akQ/MiYU1stJDlWYQGXGU
cKewJx3uFq1K1cydViChlXoO7TlqWENPZCX3XdeDbbmZn2q+Jn6/qsGyZrCgj+TBeFbx3ZF9YxHp
dj0UwB5v80IpRdzsrDMIQSgCAmzatZVBji/D9kHNGZH/PqM4UF4yhJGlX/J4oe4A8jB/tCndQ3gv
vaQToBWGe/PdNMKXxyjv2hmvlUK6KFbfU5PgX4n8DQRHGXCQd1eIYSU/KSWijkLfYOujBrNd+esv
dP0p8bg/LGpIe4EXgfts9TXdaE8JIT1Qbvn3B2Rj1z0QnqEXDx0c1zX/WfqDYwjggTu+Yr8QFxxc
16jUjhaGMhnhdr8tRFhRSDrLVarHrwsbrCVBDbdESOPegLfNEa7S9Sg5y7T6mol8kEgQhjbh5TGV
jxTGv9WlW1ii6kkS2kiR3YR1zpOF3AnIbmcKI0NFN245dh10kyU7RqFewndmnAuOPcxUj9FGJocu
S+m8yG2iCsRlMscHmREtcgjQ6lVLdk2KNBFTLO9s/3ahJQ2rZ39RGPZfrc9B6F9faxJMwb0zc8Hn
6IaRPdUu0EEH5oS3g1rR9eii7krtwWSoGQsYJ4vdPhiSCAkQYROJlVD5G9Lv4MJiUwtxLIiNW7iS
OKVGcnNGsw/Jk+LkEd0EddHC/PC93QRTHiAXdQccmBAsJN3ZSohwGFJOcnQ9K6pTtlRGMYFEGJj+
M2UwbMbqHl3RikX1w3BWqkCtCFs0y8GQCMZP08vxMsr0I0QpTfHR07T21tW/AQAh/Dp5YmUhueNC
S+cdEzHBsKkNmhCgkuQWG9w9HJhlC3wzE+R49jpmEni5YYKB3JtbZ4bnONSY+YYbA/fkISetg3Vl
/2WvzZPQAVGsAR6UVmiScEt5EOEX/k02GvEJ69c7V2/e/dR695ahqGV+PvBGT4bmbbgoJgK0wqp9
pkMyCWbfm00wPXl/0N5kLZxpx19XoRuHxsNvSRRWhp4+4XABJcDn4s+6k2siPzqkrUYlIenhA5NL
+pX/UtC/XVbyNXluX/y1I4Aij1I7PPgaBmys8rdIGVa7eWZCFn77bedgzJcWiLA5qPL5kEdLFQRl
+3j+1crnW96JTZA8D4ZH36br/Pf1fJbWptV8Ifcps4/GhIkaMuyX8uGftlv58E/5pHI17OTttbXP
ceyzgQ6UWZF6tE8zeKf/rZwtDvl0JLlKXv3waeC/+KmDUc9IMHgy/IjyI2cVC6xqfjngp+SCoQQu
LRRDKd115R6hTLOwzpLT07+gokdDuf7R1zyGjRg9Y1/IUmT+j8Av/SeSv858/AjrfNl3BCabdetj
9wWVXhwM53Y6/MMrQq7VJ+gjWZ9a8ntyczqdphfgJoWvvHPfiGspxyDwBF6v1P5B+9wCGO4ekCFs
JLrAmHAKsU+kmG1vYA9EDloqqQXJHDr+zTHYEIO51jd0XAoY7r2G8ng43fAMVrWMjWf9mHfYiAGE
glZJf5HsfYMJLUQ3lJ4yoocwJB+bMt7XrriOSwMYQNXowaR908l8L/JdfLJdhPEy5Ma1JF23KsjP
HpSGe3n+f3ASWIiWzc6xcx35f2p2U1ijdVS30UJBUMFMVSFtdTnmWxviETQhgyOV15meCTqsDMud
JDB9Zg+prPG7Q0lvYitccz05scqtMU9CUXdRN5AAhodh/E97MOw9Ti9fQGE1xX3bVyLuzpfkHIap
7LVab3+7u3m8+ViMTMjzO58K0CbEaf+QM8m4cgyxIPSqY2KsYsbJh8TtCEhGnSysTTA8aPG161MZ
3xvJ0BYazcM9pA0EPEHEQdymKXvhIqJaPyONnyg4I3QHokHrrZAHA8VhWc+rqO1hnLBtieuiEK0A
qRaeB+75ohVcyJ0HOcPGufytfwUjWsbNUS6exsh08YJGb4SkxJxp0YMqPLHO1ZmSCS0VrTmRHrES
4GlANtcqlJPKSUAxL9RBOjSqOxpItfQDCSXRxnKTUtf89U25j2iPgahSw5vdC3QWmGE0dMlPXbYf
FHDeomZWY1VgGNl3deX3/aRysWLK0+4p+jxQNrlXnhKnNnx1Qf2IEFhesQv3VJ+NexTQpAbrhNhx
HvquDrUPys4muW/bOZeHAiPGjEeQfDdOTQt09z7GbX2XQWSfDT7p7leHF59AR/idPp6e8RmjRwJK
GKDRECnZf1ba2O4Zx5unxcH6GB31Y9RsX+jR0cWMfF9LaWI3rZFvEVpNNlUVs8QNuIGW6wdRtl/C
Jjh/2L75X3Ovad3eRRrvBLOc24MxJv8Kn8N9fjTDVZHbV9mxtFBqKl5qORT9DSffcnuHZ3EQ7ll3
FeyRJXLYRrzst1536X18L7Lq+LefJsnDpBtlF1nOG3c9IlCP1i1xbNchbsP+Qb2RDMP+guRtF2g2
TVUs/Im4AaCmPW/F3HRHf25zCupz6Xycp3LmzhKp4Yd0T5IRcLcTgrdqJWcuW6FSBYps/2pPgg/A
pnJ8+u+aehwW2DNNWZJL2iT7/ACgO12wR0vmEl5MRSUN+kR0bBW0YL/709c/jNhY6Fk2M37tULDp
CGAkvZ3jjadW91iM0HBm0Hp4lMrp9WH6EV1u5YIpqM1EDtA91RNkHI5vLYjrug2jes1Rf4cWLZYI
bEZ9Z7D3hRg4izCmeMUP3L944S+kP7vOi9CZ7A4FKcoCQuTG+Z7aGxI5q2jutOyV3SwtOzpva7XR
ZJRXjiT6iR7Cfye8oFjunxnZ4AzvVi0mQFOgbhmWc+JNtPh1spEL1sLeuKLzKGH23bODOSUIBjPn
j4p/tFZAqBTxcCHZbFSIw7xt9zMbyOoYoo5OMJsCtjIdAgw6+dSZYStZCCdgIaHzcSqaPGUQqr5i
RAoJofhPS/rUPcV/sScoFyrAQ6TR1ykhdsiNMYk2cZ8Eol0WAmAH+hJjmxmo+Wgo9CAU/R578A/1
Pqhc+IMdRPjSqqPjNj2Toh29BLYjYRfei5Q7f7F9lnejkOvo+xLp5Z/iWsfxdj+1lkb19YTSFqft
hDuHCGFY7o6lRetOn1eu36Ab+KDjPI/LHsVv40tPPOne/LkGZptUCSZ9FiGDiLpb3wIgu6Ca56lm
h6fwAiCJGhdeSUfgY3b02ocrZoR2xtYS8mZm2P4qHG5wc66y3VY4+MZx5BBCfkjiWvw/WP9brYSs
QVjzQLOhWgBpntUqL37lnBC5mFmlPT+v5iJN6bZvKjsF5KzBTZnRYTSv1rJquBnVo0IbZRflfezg
sIfy14e1Ipzw0pVtqOiNwKjiY2f8PWgYv0YwZGMd7HJTWZSMFI0NMTVh5aO5BiQYpWFdRsCz8Hv8
Syvd+vNjOglR1hPnoINWPjKRDwpTgullSefXkTv8I7AAm2I6qiOlpj3ddYG8XxGjp60XaU0sNnaJ
vhu5FC12nxA2b5VgP37py0GdkUGfzOKgSWOGxOB6ebji+hrQgyUMTzHgE9OnvyXQ1oxc5jU3Syg/
9cJwqlsK9/kiM31HoKUunyOmkUH2hRbQCEJmp1nWOYuVpxTkK60VcgCzyVDqDb16W+o1WF45UOoq
BXiJSjkIyousrKfmP95guhPki44tdIJTtDRIFNrZmnLONT2pzVZJodXk7ZjJXWFKOry5qHKj9l7o
7nbezf+Vd4NeyEpZ3JAg9fFlEZfx7ocx9opdQBRQfNI4QEwoYBE/1iidijYcvUjqlE4BJvZmXQxN
clW+Le+j0uUJCOCGdZ95ZOmz7TBPbfeYW4L/wOnDVjEsEkz6Y1ligd5vkRiOGipLV5FC/md2A6cB
rXlcXl7rySy/fjk6pYcEC7f0Jyn7psQZMXsqCLI9987sNmJOC2KO3OkfKF/fdvz/SoxpTH5qQG2K
Bm/mgGzEZB1cwKndbalppUpChO43/hu0tiSPmuRjS+9ZtfZg6nJCda536ENB5JkcoyqWHvnFFFOX
ea5O9iq3G+rPHfezCGut1Zdaim8KwvPIh5MKXQ3jV8dUxKNaU5ijCAvRZmK7mhSqGws/MRyC+2vH
JbJ/uvTajSWuSHLwkn6AaCU5zp+o4E+NFMecg9ZwPyt4tTB482FKtLli+V4iRpk2i3WkHWnJP8hw
26Yo4FTEbf4o38RDY1G64JjgZAhuCEJc2DGXjKnz87CoVZmdQ47+NwZN7fmbqg30c6sirTK+G30c
tnetnWMPGyWzHqf61Ia+NGDWjkQ7N5pjN6iumvc0hwHtYgWH+3E3Y6A0YKcSxNkzHiXQ8PZWsegZ
GaspESr1Fsh9uUrdBqTl/g+0MDtZxYN9G2d4qx6FunXauZFFshIMG3pjfM4sdDhlLY04FVt6kjqG
V7BRfXv/VQ2S2QlAkgNJhupZ+NwS2FSORHAccmpw9MwRA/Yk033lEq1dasiFjEd0SS9iYOkZyf79
Z9kAg8m7kKSo/j/Zm+4tjTWqwXrMHM0vP0i2Jx0VUud4Smv3Eq9urRBKaKwwmsOr0i+oM7Xuf0bL
U2/fWEjajjN5XMPnEYfK5vS6p5wF7vno+WAujx5lbBGD2i2UgJsB7ZaA1/VUndccydSe7KxT9ylN
jCigLLR9wp0RiuUlnVEeSOxX04ieY+fjURRYYGVCsVAxrhSx1ITYdKvxiCj7i8p0g7cJ0bBtwHk6
o7Qfuf0YC8ojixdZTy6aGpUll3gEwrAXYqkcMiPqeQNdmsRSRqhny2PJ2b4I/ShGybrp5Qq56fNC
GQKpQ8KBO/bd5cq+B0ZfOhhJGyAweYnpTveZVJxhjvel+bbD49OPZ37alUofb8lvPzHyhZ09lFPm
5IAebkKPHJjX7vwM7SxHRXvwHMBgNc6Xk1YdMncBe89E+3f8LDCP1TRxVSOvD1KyHN2OXRyMMLHQ
5qg8GG2kOY3SbscAhsn1Qk102fPyrG8q7rSEH0Ba469KNXeCTXEd7cb6+OmkxLKGnli9AQeg3SAP
uTkSzA2tfRPG7z64C+N1oE4Yb0u8M5JRbNCh/lcxzlTYJ9ZUxmjK14pce+r+PZKumQdAApMD8Xdl
NG8AUsY8OF0G8Em1g/5dai2mkoLPzOxlTfyrNPhOfuXWYIylCshk1q3opI8Iriho5uxR6CnxiWor
j5CAwF5TRQ5S3KCqoJMMMhxd55LxjRXFOIB8O5igJN237bCPwHMHt7DtxCfhYzecVh74681pMTGJ
LFTixQ/l6gpRa3aIUffoLuy3MR6QO/vhXJ5TCSIDEWD97ggNt8miLjeBCbBS9CLEB/CHUxfkf9wB
rrJN13OJd/ZjgFAOTXf36di8YVu27fzNIGzl5p5HiOfS2ugvonKxFNEvI2ZoAJav0VzPJzG7a7sn
EpE1bQuitBUMFjNpz5XVuqYG0/TFF62G7lfOMr6N4q8obSB/Rq0734pncy8+bRZ/MNQ8sajob1Px
n386MzcfRXIfpv4cWtH7iQBnEvgrEbKlp9Kksjs+j7Un0cymBSbpBRW0fFwhoaO49livcVuOxLuW
eEbHbjJnZdB6XJrrxitYofbAIpBWPlZtw4mN+VUAMupPXhpLCnNwlxrv7RI4IqyQ+5JaAceojaHf
a+ODfsgw37IDnHEiu8IdVETtzhU9JSQO6ObNqcP2+cZ7FYU70YfhQqq04fFyy0WaqfhUtt8abrCI
TVOQaS9YlUixeXod1n605U5V+R4D0wE3PLmuRzA1inClHyXsA8cJE30SmfE0uyOdr0OrS98AX5zl
7xj//RiMw7WUUTbn0gZkOT/BUNYgFlkcOKtVVfPSunweP9L64i9tQGhlcBlQ3QQYea8a2nwk820n
Ko60gw5YFgWgb99TtXM9pycJoc0M2aPphlpWie7Wjs/+0kEvK8D7eSk09n8PDUitwrq42MPtWoqU
qcqf0Li8N3RqT8dEE/2ukPAGxphN4+tlT1qbKc2S5D1BIn7Mdd1PY0uGdGNJ9o1D0DsQb2/shzeE
8zZeOZkkKEe4T5WLX1lobD4VbKWn4k5qak02hzzckfZzQZcqZW9mOStcaQ5FddpIpsWbCwdFH7LA
cyRrjqaJTMDC4YDNXtw42JCs6k40sjYLa4kIP+at58hE68bbq1UjFcMvrgxmGZJVqf+GNAGpKER1
jxtvfjkVGchnB4rpO/0gIyqlaxxLolVNCjs+xPxNDt4kwqfkkLp31zhpLwGuONPRwG8B04taJZqy
5sOgd4viuPXkljCj5QcZ0dUyepgsDho3K9rXXAG7QPx+uhSwjlLIJsmsSyCBHfY+SEJamoEQUq1i
Ae9g6s7dgOn92lzvKHtagpgENUSPJ12fxrKWbFNGD9yOl5d+GOCZelwBEd9XiBoePFBJdvxyuApa
n5JU8tRu//N00CYD4MLWwr3lI41u4/Qj9hMxX6Us4Q1AGQO2vl+Ui5DAx0pUQGSHbLTUqx04YLaZ
hmwAIJ/gheSgtdX3pgrcl19vAM4lCoN0PHPjBv+xdPF1umA+r24DVmXMuoAlBx3sHnapaH0AaT6t
jZEgpSON7LjIo9Fr6LbPNhzXnalYo41EcAA6l9qkv+0IMKOAvedKQt7WBPLnZ1+c9lEPt7OjmcXT
BU2wORSLZgcrZrLvqy+sx9n1KXkwOs7GuaypHCtCJ39cC6j6rDx1867R84jDVDkF7Nqb7Id9Yxm5
mTN2MvZB9MTvHw3UY2xOtN0EJPQeyTBjzqu4PQVwZEl6noeEmnuf88U8ggCVwnLsBSIWxlagOHdU
SuwgSWviadeMwqwVaf50F6ytI70qNY5pt/pvHRqKnvwxOM/ga5Adk1xjyJH9Q2JYfxtlKrzqNcQc
ITxMOUZ/JVY7MeQ0O7ZLolvN/JitYlTkbr8WhPRREwuIEKLY/l/YAUE0AH/fV4gX/36KaKY/3yG9
BVnr2jWaEEPCIueNjzBhCPJRDdLQ0hgw5iGEgGZKUyhZ5FS61R5qti2EpR7ErYce2QYJFC5IKyaS
R4hO+8/TFR0vhD0P8R84q+VqmdhnH95TgsNcqn1iFOzJQnjeoAXGgB52b8fQ55XBResAjaln9eRZ
LJJ9Kq/IBVbpll4eNJG8jJGC44T8ikOTWyD8jHnYatvRJQfsprCNaJvUW5MB5AAPrMwMenJ7n3M7
0wM3WiyeGmHG2/r+zlHa7ydMV0GbAZzxuCTQJ8XpLJchIMt/nlw7fMcwiVk8D/llngAbk49wnTQ/
Yl3YePjK0fG1822pwX8K01pUZJMycNukVU6cIgrkeIgtOag+IIjMRJq1q+G3L3Hs4avuPHvA0JjQ
akNAyyGKMvfAXbdzRRxrXKsuuWraq1B1medFZrbOxh/Ws7/7TMvWgX0PBP/LcC6r14ZAw2rU3EmC
nldMAb3JTbAglfLui9EP3P1N59pFqUjkOJLFF4rvsDhtgeFgtxYGbTrbMdANct+2TyuOppi6X2XN
yO3Y6mghx5ySB3wwif9vbBGUi9xG7SUc7jMuKfcd0jW1jA5qj12Q76P7ZNnOMgafxPMap5dtw8CN
3VB8qJ5AM7bW6WWFY4GZZryF0ILyn+zhkcnOcYjeJzDBLeSgyg9g6oDS6ytWExhvx4dDNk8eEOuV
c/yqOFrEK8VzGIAoXdi362Q7tSCm+0VT9eV5ZUdBK1zQjPqdW9rG/YtoFvScZ8jltl4Ekyw8Xt52
GqUkxafjLV93CeFPPW3mg/d41uiN9KhWoYkSBW88zNVlB/Kt2Kk6PeY1tGZpJDEN/1iloOwKvCoh
TpU+8aVkW1Fk5UsJlfAUwSq6IHf0h2w08uY/rRCgtRv1IZaTn2I8uThkjFnJZtKC1DFm6Qh42Oc8
5PHa7oigT9is+2HpzagzLVdXYTiDUAXSiDGXFH8+KBVtmJmq0KhoVr59cHjGfDvdFPzokLyU/u83
GQS0gcf3sVu5OjHQAtmBHCvABJRsDYz3Pj2oJVty+RNu0qYN4TThr81uls14xSsqrtBSzyV6xa6V
oH5f5ZHrWx2JsMhx6EbMcL/j5UJN+0SOKPtAabO1EbHv8cpjVEQLhx1TJmecChWgkOOcZyU9nIrK
j0TPT5s6J66Xl5dN4D3vLuBpmIcxweH8IqL7iqeE5TkZO3RDrwt4mKT4uFhuTQxrL8zkGuh7fpe5
EOeu+WRnzq70FkkK6jo5A0qru119u9j2mi/Vz3haA46s7h3FOhI3TyXVm20IOA1UX+q3NRBRxhCN
YZZ1cjkAMjgTbryhIRCXxNsR3q+g1HhrRK6tJIVhf410JkelZGHOMIPfjO9Voizi3mjbhQR+yJJV
adeN2Vvh6FqYUFTTa+vFKeaV6C3st5b7a0FcSfaS2LrYtqMrbnj1zuApcVRzWNUNxJdrg64ZA51n
VJ6iJIGjOdiQ/rDZGSrPcOHO7fL/9eb4vw0QOyQiIDggl/sDnGkWPMSNcHEf767H7ikkfKVThbNv
5gw6YAmo1V4XYQNy45q4FtoUpmgZdFWFDae3vkgipb+MYzmB5ccVNYjdTSeh6XO3OLJspMXOdna4
GY9i/Y5PP+shMbcpvX6QuW7qP+vYBugsPRrChfQLCgPezc04BqSTnHQpHNz1/s6Rb+5Y9rdY9Xzt
4Q4X5kRhyF5GLTp+sGwWEtoviXNGG/Q9qLFn+xRJ4N0S1Pp7gdJVQb10vOZX1M45UcK4WvnLk6Kh
sgVdMgoJn1nPXulfOwKwdPoBmrVBckcpuW75EnNf8DeotT7ldntfEhk/8MsC/N5Jg09mU13HHFu9
S76AzO2ggbj951wOAFfb5TzEPW519SdCvjAR8fpd/TDiYdTGxWF+m8W2TCU/WkUzPk+s8Rv/6DC/
PrD44KKw+8aUbpOk20HvRq4N8+higWt/JhaDsdCX4F9REMjpS64rMhNcd9eY8J3dkFG1ltZA4Yre
HJieZv5oDmE4GW78gFLoqqIkCcGWH43o1rqF7i2vPv8vxMYQkF8RteXyn0NjoqTWf87idEJsGKrT
Hx30ehiDF8Izwrw21dcURRkjgmaTAriksn40M4YQZWdH0fPqB89CZMA7HwxgGypRaft79rgT5kxz
JtihLMpo23w9Mu34JUm4wug47M/huc21HJArIf4idDHzxYnnkSHXht7pFF7mznR2gAa+iBPt6Jod
viIdn5DLcfbfk7Rerj8E2BFeG476s3TcZh3ulS/YzWTcSk4kh4jsNhW7y9hHAXrsAbfclk8xPv1S
TVS1I6izmA24MDe4wN3HWkHQNp5yh33t59KhQD7JEgSLaornNz2JfWVvfafiZGE/AaNFfqUfSOZ0
FnWCM92FJCQy/jcLsDQ5mXQv1F1aNLKYrOdst77NNv336J+JENRa813CWI4DlHnrY2GeCD9mKD4j
/VBJpa8I0X0uPvPPFKe+tkj+SDlgGGshA6D6YAVjJrDchOwleKz8OK8rcODZUPqGaPSfuXO54KN9
cpFoSn6BHmurw9wZcQSiICJwQXOnZpJrFemRr3T25TwrRsQADFcDot1N8tPSUGmSYFTMKa063Pju
u0WVKtCP+o7AowBdu7VOXp7VjgLYIx4/S0RcryxotJxmJZkHwcgp7Y+vGRCiHhP5G/eNyKPOW7br
nWaI3wv+J9AIcqM3F6ejD4qML/+cSoTMsOrY3fAAl8aUhuzOU7pxKtyeqQlYnUpBg0ydelUutxbM
dF5KXmZIKHsysid+dox/KrtZMnQa/jbNHNncdDn2QQ8M0Xfu+eKQSHjKXMnHC+Ku+M7ZkaJXWCQq
TBwqVfSV7u9v2mWEbxE7PNafCaGKdWJAp0UTMFMS57iR8EuTentYo+K+CCDKV14M2v2Muiam7T0a
U1S5cqdOJauFHcJqiYqjGrc0FofpZXXWRiTmKoFwq6cgChJldWFCTplJAkxQpOM42mBQ0UFaK95b
AFJMyxX87eNgzG09iE6xEr3sjMMVSYJRbA4fl9olXY3kVlsXWjaopbgcdq9OVGNFVzmpvZXJEPXY
X02nBQws9+6MTs/AGOhDtWWm30D/mhVdRFH4U+EJCWaGkQvpzTTKTFcbDyUuiu6bCCJYPWWWkPDA
jz6Lr769ndENni9M29XxVZoN3T5IfdQPr+/BRomKfBrUv5oQiB9sZGMEx0HPCn8hpJYQ9Hi5ZiTW
ENbHS/AnZZW9abVS/vobaJToIURrqCJWqGuZ21mwALxsehnNQ3zvKCSJWk+U2pX80lqx+XlS09AR
1SOILYbZAO/eYJWPXaowR+znISIkL3sK5HepeqQlnvdci/CK9BidUJZgUM8+Zg+Thdnr/7IUURox
I5PLQ5EJWoQaoSWKjb8tVeYw2vXS5kK/ImIzBKKGmJufhvaVQKS0Lsdn3pp1cAk+wXEGW3N24UM6
nCXgYHVMZlg6p3UVwN/BYZEo2F95LT6T4X2TFpIG//0Ume4BTgPui98hkVMVO34xlULdEdJSlOwH
tGdR4XS64ze4bafsiqgm0Ne9d2oX7zjwsEZVnuQ210DCtu6ShoBKrb+JvpelLR1/pcbxe6fL2N3i
LmRe9GJr2SfNX/cLbm5nOLEBv3TGBWZ3GjUC9KVKUalWh6GYgNYCUxfYTF33TOQAwIu3prYkZPDu
cZXUJqJBX70YRztOoqX8xbsvqvkn08+KqpV4Des1E61XdZQQv2V/YUqbmQ2Sxgdf20IuxLp8GlIG
AZTAvZhkkfaSGvdF+TfB0owBtPg83mtziSg0EB8MlmLnYGQb2ABD12c+BREEXvAxTmzag4/zyk+x
xC4YgZZ60NAqTD2j1x8tGF3hdHgQmvKENULlmb0lH9AzCoUDEjXKgLLfjSXFMZyxiTMeiLrOWwrL
1CBQyRq9ATietu00reAsk8NG3mnXu6LGQDDLT5XbjwKAHdYBfcjZFKOwf6m0b/OdHvczILbf6BTB
rQBFBugJ3EWq3Mwsa/+yGUsGg7iOyWvLO6jy1vLlcGwmrqw2FQdapALTM4fA4lYrSYYT6pP+ruNY
x8c1iTe2ykG5DeWBsZ7963CH79iYi7QptlAJh4VRou6mXoTsZl0x6oqHS1n5Lb0xlHccc4UqYGsv
5CJ7tOV2CwgW5Yzz0w035FhnqvIb7bEH0PAKL6eGaaWP5lxO0kh+fW1hsQBDwPdDvomdurLA6ptK
cPUovvNOgPQWUu+53X9ugsPN8ZDR1D7EPshZOvdH3zwq5cj+gByT1D49SeZH4W+ZEKWd0oIY4Mep
APq9cMX/Ao31EUhcJzShz/d0DmSBglKzpg2zBV7Myld+a+Si6nEQX6Jy0aWyo2qhQiAnCz/LCNz9
KgqkBkh2e9uUA7U4M0eWCFJHEokXn8ki5yLoT7Q0DTQwOZ8QDvwHdWU6Hx1JHfXx3dLhUJXI2WCU
4fFWY44aS84nRnLESFxDylVJerlalpDoPYAV1tFCY5SPRFVgC7NikGYeh6rmcxdOGzmq8amGK39y
AO2Q3mGdo+NM9nKNaI/lIS6wo0Y59Z0JZ9GACS8IxXIBjiDq80rAdP5HyksF36UQa5yi49xBvxsM
CmRwcht2GIWXS7vnfMQZi7quV24iIPLc0kzQKGn+/hOJFWGxyQTS8G8vAUhQDRrL4+5AQx5/TyuA
7nkrdoo48PHQItsmX8WC+bDLRpXSDlOwFgcCt2cKnT/UnhWYJRzIFwoIoSe7ZNGt8KDW3SkZxvhd
eOzL/jTH3p5ul6glWdT97+QI+aBIonAnaqzdC/jzgtQuabfJKW98spEmFFqosUTimchhDXfZ1XM6
P/s48BphTac1/+a3vrJ87D9c0CarVQJVwPQQzRbpTiU1EXUFa1eI9hIUytqq1nVvDw078KtTwOcu
p+mfVRMImxgGYtlEi4A/7ABs20koLsfLulNeo/oANFJx38CygSjomkOJyGrZQgmYPzxHOj7dWRDC
0yWhN/i2fFkcUB2QHQUHJwUOtpQz5rC5WnhWUOAx/QutOe+QctGXPS3Y8b8Y+yYJPiXh8NP3LSth
RBYX713mdT2wZgQBz1fVv5u+D6z8nuRlpXexaLG95pfZsls1gzhRmlKLvaP7ZpGLe8xrJ3qEUKkc
CoTdhHHyNlJWX4l0T/FwpWfqrykriL8yYECQh6VKIZn4cWTxExnMqcDXvQj4oLYyYRAh+7WnwS4J
IbBsPXPAqWIQu+JkutJ0QknBgejB37N+2FYBvJ34zowPmR7p+2gHWPhGDVGwLVBWh0xPnF33BPW2
HGaKevRFLipXHa1IDaK9p6HCDl8HznIJLgjXKbHVQ89TlrzIApBMaf6x5S1X2TfoCJOQMYMLPAmB
I9EwUWXKC3ewu03PQx3xkxdRkj8pDqQIckvoZHb8lTtYPhwN6RasiufKYmDIxtCsSgZCjKpzJjF6
m3ynx9FMNHFoLxQvrL2Ao86oXuL0jKOO2xx1MMO8OGgAOczPWx40Hz+6tpkatR8+Ev8/0rfVIPeO
DPkAxaPHyc+FPKZT+o1Hv/Hopaeli+VuUzKK9ps3upvvpUoU7HvOPJVaH0zkCq0YwlNfQgKkVdtV
HhnRpu23jUxhdc3tdT9CQqbUFg1XR0EJ/om/I+t+B3TOK/2bpVdU0s85cJntG/MywOim59/t0B64
/oMG4ywf+HYfD+PbRRCVNcoopu1zZnsErokgUJc6NGhkKMW1PDV1NW0w+ZWLvQbdbXl4zemM75+q
Mqx9WbqBLwzow3Vca7ADxai0nAXePjD48WfLjQIS/ofUev2gRKdDvowgRDIR7ahnWyID5N8NuSNR
w8qfBmIiQoyi5lKdjOPUQhtu0adAih9Zimrj88mj4y7jx71DhQuwEWpkQ0PnCpPfNbyVtBmC7Ptt
zQOF/G0T5RJkM3O/Y/u4tYHdZH0Gpo+3yMW9V8yRdmtQe3fw3jYo5Mq6LYDzRTT4DPczi/kEArLk
N/XXsuFvEVP6XtNM5n6UbLVkTl+7XNySp+1EyYc9Lsuy75Xf11bH5Iv3ZO2ofzfMiuc03ImVxSar
4iHhM1XSqcGbqzF2sFDeWFsx1MEnQW6DwDA4mF4Z84JJ+ngG75W+NICMj+0EoGxYJdWdjgn4yUNc
8SVU0pJ422qU6L9o3pUPS1PLNX2kOQpSOoDQuWXa8144LVq7UDyjI2Gw/JUb//SP+pekKbtiLYPt
mRIc7hyLBDWyWjJ1IaMuLPRZ+dSsC1KazhvaSeQHoGkIFOzTGgPvlIHDamny1DILOqRnMiUFDJSR
Ml6lGGtXgm71nU343J/ZepT2Ym7Nrq8nk1wnVQl+spyhsrkDq+fymDFrxPYdyx0PC4gSqNwNCzT6
28BEEexNNxHJorTkp265YDSCYRT7FRPRfzfHcAdm0VxNxB+/+lM+jjzHPJhFZKmkyWQdDCQLmD3k
qMPnGDfAlw8j8/DGq+a6RpPwINoAQZNS/59hMZ3dWaGvBFS6aNU6gQPCEA1v2YJrjkUXm5DXkjr5
DCYerbJFCIPgiw9DL1nh6MZ5Kb+cMH3Pum1B4qGqDBpEcxm4FJLnx/v5aWQwYXwPBPsktu0oOinc
I3Ooagm3mAU8DEgpajDbT5CxiXhFVVAV6UfHlsZWIZC+sKzAwwFE8Ue06Hl/Ifh+vnEHBnB/ZF9I
rFiEMzoGp31CMd7Hfg3hXYi+Zo+D02tAgpj/8JzV6SBvXl4bsV6uk0QUUUrYNbytap8gZzjOfxEI
e79Wfzfc4n7OeeL5qrxKRW29oy/Gdu1uOo/XD2+3ATF2/8BQzHXwAiW8PVgnMKi7x6pl7iBC8rok
cBgz5lNdY1K4TBvrwH9OY3s2uRnwBkyq+Gc64Arz/xCQtd9s3zHfoGk/SnWTZ2h6mHUe38t2FUaa
exZXWLoAdMBNXSpW9gvzb+jS/FfWl4x5Fu9BRY0U61HXb6p5Qa1pUDxgVPXlXykRcZCG6aGNHGVT
c7uvS02mlUWg1k8y4uAcGA01p7EvhZFjfARK5FicEgwOR+OxUVHx/wP4dqYHH4p33c+XeDwFG8Yj
5KfdcvD72jN9PHDTSeXYTpKT4ylr928NQA83r4X2VHJq3WYHDgBLipYepWjs5kXUO6ezUnK5kRXW
M6/OJK3W1ApWyHzPSvEY+FBeJWgliwhHbk4JhdqOrtHOVBVZqBUu09NIVMwpsvU3TfaGZbVfY+n4
dJ37WwxhVLu+IAeAGC1BAWiCTBur0S3Bh59tulyriqK0KK8YL3jiSJOunZ2ZpJc6kPmiRKj89kQ4
QjoyEhHfKhCG/F8DInb2Sci0rgKAGenfPB/lU7oQ2yINHM7CrvdXIp4lqQHkM4XCEzlnSdOCehOf
gALKJvhfzZuDGWOVUfAAIJcrayrUGit8256akAdaUOQJv+yEBDUU3dRdZwAiX6+XUNl/wSlWk4XD
tGc6KjfIlDbfpRuoSgsx0buwdvZPGBX7U2CfSaqd69fZY+v5VkApyMax25djc/jjnfWQ1niTM3LU
zrM6PbnyEKlR7eEkGgVw4ukweQSWYdV6yXgIH8wgcHZJLBbvZ8CzC7vxkupoqOudbg/S0av09UFP
hnFmto6DyeIBMSszWRYyHTxz7wYZFK405TGDR2KQYJnnkEJuAIrOKymM4pdXdZ0hc+gcosJ1ayPY
mwBYtFyHGxQErFzTV3ii1doL+K1FctCaXCrOidELQG7ejpDzC01nt33Ndbz9GyhZc+wVrsaAZPKH
Kw5gkJwF7zy/N7G/4YSLlG9RJyzmmqMfOtPA8EcG10HmBesIhweQZy0m2MG8equxT2uu3cIXOnP7
JYFpGEXwVda4OTQIQMLGMiO1yMttuc/Weube2hPlmGijljSdS5VlO9stJbDvbRuopLbEvEfTEa89
XMVoue0iJOIZGgseCkhZwrYvcWsGGXMCj2QrN+R3zSsNIkroQFkPSeCbLrB1iLPj1jM1ttNnWttc
7iWGvogWrq3Vu9s87M3/HlaGW9i59dGOeC+NM9eIIPMfy3NyVWUdX7cFbSJrc9Sr1gx39Vw0+wui
6MocQGkoBgXHoos4h8ua14bqruvvwHd0qMhYH4LKor3w1l1///jmQiihvs8Zl4LCVub+dG8cucPQ
UuxCGKFB2s368P9/3yFshadwPjHhq6nevZ/Hvihm4aU3rWRriM2wc1LTUQmWlUaPZ9bKxJ/r3xnr
zNPewqzd+WegeXZK07YRu/NPdy32fZ/rko+/jiT2xqQfOuDQp3HWwKQtI8U70TVgWRBB0poNg4z6
f1eD+4EI8YrgW3NFJeYijHYUu6pSrxqYSSHaXVrVNiVFojCt290bGtXhHCE2ZUakULHUGBQJapto
Mp4hacoNlnk1dmJ5oAdl9V8q2kJQ+HMSEI8zNXjqKYjIOwwNihNXf77a0b8uhGSoD6nFlW/T1OxS
/QsS21mU6+oz6W6abE7kIrotMFSzrYmiJtA5Q7dw+2VXkpv199z+BG7ZP47tf8xDYMjAtLjVt3kr
68qjsnOECTdKHMn8VIRjZsUGNeZfjIVhZbNcPNLYDqLffAcl0TJ/HJIHbut77eirQHuc2WC/zPtW
/4W6cHezV63LoN36Cvfgc89rS+TcIa7dO16bHgkrQoc4DxuUzroTteLBpJyg/ycRazyF+pf3W30b
iWDsJ+fFM0RMbwxbN5QZousemBGPA/BpT5Kycrz4EFLra1pAUV6Vf8WATvWwj/vcOv235Jb9xDWu
3tVNNje5edjtXU5+d/x6UD7sgQhZfA25GyRr0O37T3vJBVJ0kcVPwAEKLxRacv6EMBsGIrVEq9ik
2hKrtfTG8Q5v0CwuzKT7He0fcow3pATz05SEyK6A5etxciFfagXXLMWyotSkHUmEkYkbOSHWhDpd
/25ocm7hpEZMRrk7N0RpmxRTHBjK0bmCgyw2u7qnSOeG6fLjskQ9rmhs+vw+gPl7WAHtgJ3U7Ias
fAWcQOzxC4Fjuqldtm13y10f5U82jEXP3sHmW9w1suZVvpko081/Abz2SLuCjp7bnagyXq/DJd7F
5tyvNomZyR0pX5ffskab/8Tmpr/KwDpT6cSgaTJECVFNHGI6qzAZWdrql6SDyiU9sexJmzuT0f5/
yq7paSdNySwatYXKxGZDjlrphChS9kEZKFGqfqSk9Fe9hu07MOmheogpbT3yv5fUf9V26yBwX/Ce
CP8c7xY2mooSFHIcQ5Q41ndj+/OarbhwPDsSnNQu5gz+lBkF9PWvDWi91X6ueZDJechNpf+4zsNh
3o3rZtHbCreTy5Q0zl+iSNj6gPhH1fHkh7np9LoVEMzpESGxlImu3laHqRApzOlvR4mp5isnL/V0
TnC+PGZoSR76LFIeev1nv26DsVfo39TVa9SaLcoEz3JgJPlU2bS/Jgp49LT8vvCSZn+azIEEcC5L
GAA6Rnx5rz6eI7tCXXvUx2pjrKsEQGN0d1QraYjSLVnImotqwDYJ0d/YhiHc7GvFbibQI+l4c5tZ
N/73skGrgPI5tIKQatNgqiNc0Mf9RjUf5CO7t9OxT6OR80UZQZ8k2PeIrXerAm4qqd6bHMPZGWp3
Q6rNCTSCm3B5E2YRkCysSWlStSugLJexU1F6tuS4CQoFcIK9wc9WmrG4bPAPzya1PA3fwNsNd3Aj
RXunkkK4InE5mpRCZOBrEu79ivCULPR5Yp66WRH9+4mdsinppF6K7sVkTlMz7icJJ7bEivLcJ/yp
2hEMdfjJGGxoK56U7eBYMQHj+gAvvkZYVJV0BhSmBxk8ZYvYpb81Q5x1jRCeunTnNfTBgMXm8gZD
K30P6nYss+dQ/Ve1IV8+ltl5oSNUCCX8TdvPPO7yKFIh4DYuPImaIZA2vm1DC8W49DTf0Yu/kcX7
fKJgql8x+e3sVaKmogiTpy0GUdzrdL9z6JRsSsKsPYgwdHibSZ6kL/WJwNoDraEjNPglhSFbA31Z
5Bg9Alquju2wxYnT7Hu0iNbV3o6q3QyjD4/aSI31msPVeYLgY0gpZkij167UkU/B4HWf8zByRqsN
7u8M9QNEZaQTwKRYZJ1QKW/ooVphs5/qAafYQIKqNLOcFOzXH0aOKi5O2b/uk7exiSirZE2SCeUZ
sBp9uFDDCp/uz10JQcGe6r2Vx89j0jp800dDo6F9s+SHSal+CcqT5pakr6pTOeLb0CUsc8loUTUm
EXpwMoYCAFK1v1lthzsRQvqZXIV3jNwKl6dZyCAMvZPkzs9D/vFcVlaM/t8QCMgQZJ08hj0aQ7AX
htvosE1xFMI7N1syC752ACibejwEYbizxcemMNLopVhPpgosY3wmE3Np0f+KmUFUOnJ73/0mQ9ra
AUCt05U0ABDsT6avO6ExtLHM5vp+gp1TSW0g6tyCkBauTIm+3XRYcc58QoHq8JVw8WMlcK2fLmXY
WjAv1dtuqwpvVTTj0CrCOnygB3/IykWMb5IsfL8hxcwfy4OiDwRA3XeLuRfCfsuMpX7JxwzVuB/U
S5OxTQT+xc0gw3NttYiqMGgu0vvdofHRkcIfRnSz82e6L1BOWf07q+P/Y/rO0LPzEP72lB9U7ktN
q/oXJFMMi1TlGhxV/mXDTlskooC9b1pPoL7nySoAru3PTMs9T81rQZ7+ObNGaVVm0WzAlYjgCTAH
qY8PfZ/TBrMxDcp1RTpkyU7IhKgRwGP0PZvm74IYrqv8etzzBJF4ZaMZkHe8QF+9SeL2tPD4wSnr
oZ+V8m/7u68J8BWInD8nZVuR7LkCSdxI5RGVxn2LagiQIwyOSYNwu6Mt+cI1rnofZmTJ3vqXQket
5EVwYXlmpe2JTm3r98jOlc/iV15k941e8PFIxOkSLQv3+D4i4hsHUExzqyWbYTRtbexBYStKBJ2U
jITY/qNqzoaSyXgF8J5df1s8GYa4efh0iVegoJ+jT7v/FAQglIHeUio+ebqN+wVp3yjeo7cLOuwP
/q6p/id6vxH4m1yKNA7sIEsKwQjFQTEVm/B40L/P+jWEi+6QMQYnu5RFpK6E3t6mTv9hMzit3VnU
Kec1kOTdXwPNXKqFrUPKW855BGuGYw2qTXtWyN4fjg9EJwiBU2pry3cG28rs6WQrljxxqg6pleVe
q5yTdMUh5H5eR2wn6Xdq/dR3kt5LMeP1IPzPmhnsaEa1g/g7bO169v/TmS4JdmqxUQqgzltc1Yp+
2q7cE+z/XpUqw+P5jPxQJT4P/WEIo/JZCRx7vu4Hhk+Q9yozBM9ceJnIEkrR1JU9dKX3BLvhKJU+
WEUURrI5kGhM5OSX0VjozuGogSZ6dZ5hcddneYHckoE6xkwRrAFdjVRy6CDSRiaxjCTtC2G6Mp8o
SNBGG44TpkT2i8cWg0hCOkDXqUB7zL/RG2AFah712wMUPJIRuMtFfg0RhK1ZRrYJEEJ/tBaAfZsU
rdz0FQ5yWLivYToDeQQwP2ke61pGk5Ro+w7qnxsaoV2RJkrDNABvnA7I2dDgB8RDhx8Xg4RRoJGA
kLzdOQgil8t4BU/MKR2oQeESWastqahszLWovRJEC1T/duXxAiSGEU1x6MGB7Pbl86Kl5G0lohRC
FriUFSMmmC6UOdcN/Fqq4CIanyh4g8ampVw2lkUuBcwPvIifvIIMF4ugMlTZABOOBkP3K5YPOFPR
kj4gh7I4BlueHDE0pzV63jANSPurQy3+PrMegEdoaURFsuHhaCNHmZ08Kj39KUV+OXRusHQJm15z
MGB9vO+4rNBJcQh79RiQGcms94g4LrvADdwTXuHzYliW8NiS1UjnS4MSeRmpoRWIXMBvcVcx+ig/
MGZNkvCre2vIdI7XpKCBZWTWP4+b0frdHWAMXRs08yA8IzbykM0O7gQbjMVCVVgKYrGpyZhFfevV
i0pvyQ5/IvFd0Ln0zQ3mymYfIAdc/JXycqnG5VV4UXhhtqwVWDXJhHUbR76Uaja3UfRsTOUzkJAd
IV+eS5qLwl8VGRa0RM2im4RWOb7GCm+2/NnDcON6+7vCDbc29U7Bvc4yKyABUHS0jM6dGDsr7g2z
pQnLNtd4o4tNGSbhieTTTry3Y4DvOlKMGfTAMqmHiMg17ZAesekQdG3XouNMmAGYm66JB21eURNf
dUEZVs1CDLN9o3lxdmtrAPME1V3RjvupR+W02KiyY7Wkjf8zKm5Gyz0v/Xr80F7G+Z49/1p8mLTB
aXhtghhIjIfxOJajjvMjbg0uSAtjDmoSVs0Z6aAbxReKsBqT36bz5n85ithkXtnfEeXu1LIDlav/
lOhoP0jNbWOMOUipJDlu9qev/vEebtyvnFLenTFmCP42iMTvMPBqNx7INTrl7JWQwHziHaD6b6uf
tFDmGEJAloraCaQP6SXxJmExeeqmx29mSzxMcf4Kb+oSF/4yU3SvYogXXatXSV7hAr3RToaazEAD
vawQbLwdX1kPoVC4oKMVZ5DGMT17lnWLo4mZ/wv6QUVX+f+HiP1byYmqBGpRkmt9kpEubvw5NnTr
7nc1wSMrgVlTwSRdlk27o3UE2Q5hJRMEDeZeLZCn09gmusnp7Rx64zzZz+OkMpkVe48eH9D9xZEe
Cm7jd3L1kcBMRt5k/dNzx7ssOcZLGU7kFVRQ1ugQMJTIVaoVi9R0qvvMhzKQJ9hiqiWf7emNBeWk
j8EUGMXaVgvihXIi6HZng2ABTIxSvMDkEY9VVHODXuhZYqWcy1V5RQKIDMyBUBeInyegZOpWgWIq
BXvlDOayTJEABpzYd4AoysO520qcOqexSe0t8ktly8yOJ19T0jmZ7RaOBIvJQve/06MZuqPg5pU9
+SVVZxBul+HmcmuSwLszwRNVY+xUrEaO8FVjiArM6GSHMgfK3CAZC5YQvZzeH3pjjDiOEldkbKH8
T874yB0aaX7vsvUipHTQ24anZiJiK4zhwEBEry2GI5v9I+4FZlV0H7R2Cj7ERs/fvd9lczNZ3LY3
4DmY0i29Kwp7afoyu5u9BDsKPGtQLGv1OkvSgHZECSJi2BtdDdweT8+gb6NjYPmKriC6SzecUTn4
KaLUYfWfHWkQeuiH1HCe7LzOkd7xuhtXAeWVdnGt4ln4t7epvHlETZOUkjGNMe5953mqzDcJ2xsq
QfaRu1rwQLczfhMQBI9t8k8svczyadWdDkjuz+DnZdPS8ZcJzFHPknuZ9NWEa5DY4I3H3O4eTZ+G
64C/uT1/b5TDFFxMzPn4RGJjgJW/KzIwpBxukqh3BDdQ+ZL80YE/wtXfR7H2iqw6lFR9mA60yGRP
ntjnOUBBSiA142eCMGz8cM0w8GTDpJYmDP2QPd0ykJJtMPcd8dX2Yx2IFu1p7r15/hq5na5cjK2j
3uksqp7cp9JCklLl9bukuXuTnccuiD6n6ZMBOi8Z3sgh5+LUow489r207G3EL9k2I8Gj68dMyuIE
sB9flIHkNTZNI9gx90gG6mKVDfQJh+GvvGFn4FNAmHRBfyrRYiEDGKtwQpLl76a4WggNM/RKIPnk
jM/yDVw8NNuU8QgIjFI+NeQQ+QkhWtJ0VXOT6jlF37MS/jnSe8PxsPq/5A7mAQGDM2D8TJ2qEh5R
TXcBSVOYqme7b5hBh2R0jNz276f8LqKmbLnLwUUwTQ/iU+/9QfcmAyEVhCZCbZx5yzFFtYKTTqEL
GNsyYElzF2RHZMPn3i7h64w431U1XGRyHqN+tDkaYnJ9n3IzQBYKfJHhuSsn6CwyWpT3bMUT+gq8
vq+75/+yYf7x+sYM+doHIZ3Y3TIrLTPN+oQXPpgSpiO9s/aFyKLjqxcDmrYfIzMOWg/5tOOB2Pd7
FKL9xEOypypED9msiTZFn9tKuLjJWRLql37rcqPrpKvybrI4Wgl4xdVGdS9BECaLmYc0QgqFAqTU
t2f7e0VCugXuz/sb3mrZ8de3Y6XdPGn0dih1lVlhkCH8Ro0P+oGwEQECK/eG9jSQWz2W4QLpQR9+
wW/JdoEMJ/ILyWEoh+FedCFLXKiug7sV4fZR3muYC65FGpix5TqZIufKEnytkp1AKnrK65E8BJG1
AM+m/ParficPYCcMfw4kGmm0+dNQQsmvcWfAq/7t2xqbC+Hxky3sCfPbFQa+dq6nRoubC/Zn+R2n
KfYB4HQ1/E3ZxLGgz1Q3BDVZKYgAbjRe4X6cg7cU6K2d3+CRbnTH/kj9q5HiFKpe3SIQjFgVey4o
5cEs9zxn1ka1F7fF71YPbYlXcJiZZdU+oZWB8cLg3QZQ+yayBzuxOB/gMOkCoQyw077QNYzu6iwo
0VwYbO6gbn9k9NH7KQXKoWIgu0nb5hbproVHD9OVdfjgwEn+tEymI1/rY0jFh3GCJ+C2yqy1aCP2
qRkeH8HODBrZKAsWDxvLLiwIsjtkULOjx37nPBvf7KkgTCde4pQ6FYhqjvI+qSUi6R0uLyVEZp+0
QpvHDvj17Sf+pD+r6/m4VPESPd8uQYvOaSZnuRwzaLuIiee7TEqER2eL6wFEozI7KjWD4e/k01rL
KOHhhu6/xXSGrg58Xqq44AFVPsBQ2Z5YrqF5jqD62t0MK6/YvGPAHkIvR0+/yoa08p+GWtRHQXxn
/SRiyGCq9Tr1ATW33N7GeoLzgJmJJvnbCId4J0Nq3IhRBZPHHRoBv5t9LGOQOoJ3u8p/BLfXlWVq
LUX76gSWq5J1mEw7nFDBxrDbappPr3thRQ7IZPZdM+iRBFNVaZNFOl+w/wR61aORpvzYsAVm+7mY
qDp9jvLK3cG77KAIt5q9CERE97Vo4b6+kSBiqruW0yrtr5bMUNPkrGw8GdaTYjELWtgrA3Qs6jpR
opwjfCn51ZkZ/CsRXCewvdpJwkDSGLDRSfp9nT9eEdohqsG3kxfncDiQrXRnn7l5R88SRqWu32bT
6pLgUx5oV9kTODNfiVx9kxrxLxwPIgZrYslNOvUjulEgd94apGwN+bunZAdr491lYq5gNrwLc2Pr
XKI7x6hGbVRwa3o2mj2WBdPWwUeLW8ITxZRc2Bg+C0LChSL0T3Sjk2eTdtscTB5IbBlxod/orsri
wQeuqfMQcrKgZ3RQhgHcqL2G+/sZtIY7liUhOv/z1q2q5d4oIX+VvNRl7C8iMowTM7mZhH8niO4M
qGNn3syfqCKxw9TA0SDxslR3x49jJGBHz82P6cz9ldGfla/+GPrIw+RpeXdO9UaZGjKeQCqNhSqd
vcuEvziXkZAXNKfHf6p20L0rsfYxsP3Qd6sIMz0osFYVdbTpP144/uo9To41Rwbl9bMZDw1L+5Gh
pwfHSqLrpNCKORkselUBmLowP6sErJp89Zyv0DT7wmE4Ru8iAs0MWFg8paraRy5QMn6/Tm6Zdf+g
X/Llp8/bsCTzCzCra3lLYuS3lz0437CPVVC7V2rnZ1lx0sAyonjwoUHIu8qLXpGisWJLHKa+pP2f
04eEEbdsiEXLQpDmuQrZit6quwYNgllsIs6GbRELjZVKQp/sceIUQYNSEPfR3ujvf/T2q9mbB6PS
cFj/8x3RE13Ro/Y27TWHIKRNYoI7rPxSrNJb0n+uNRZfandMy4PSJz2qEJfJ5Vw7yxncw3mBwBFl
ZIj6lCXHWT874nsBEWpIdDmiYwbfDnk67loeOkahv1BBYwkCGn6Flal/7+oaA6KU86DD+toLX0Fx
YGNHe3ARMs6+17JRAYj3HQUiOMPYg3w/E3pWqXx890n65qLyajvUBGSepmTVVlZIvguatOjHYRn/
9Edo23YgPjqZUJR87y8O8yl/5s3IOr07ZTRUUH57XRV9e6J3UZNrhJHozeJsR/3Xu6GT3tHhrlGV
C0XLb3ZPd7ug2ooi9NCzA+VkEYGQQX19Ic9ejtcPtjraTOWkuY6RehG2L8NrVYut4BPK9Y1yVjZ0
vZrlPFNqvq+yc7xNVjn9mxiInzIfzRbx1345GD+DboHZ4PpPyfmjgcRGL43W7DG2Y/bGD1fyyFLt
4dui8lCLaGhblYMRQK7EDGzr0ng+YwnKtF6OfBXldwHGO8lLg+uan71ALEffzxN9PB2EAK9W1kNY
TQjUwf0bP8KP3JRoXhox9b8CrpiMP6PTATpOeVLDwbk8gQCKUktvA2D8sdARR5NQzjl8plZajOv3
+ubhZp3+cZtbMOJQrc++JtaOGo8z5YKvixkv+ZRQabggVicxQDwAWknirvoUnMdB3pGZouuhiilS
+iTc6GZtAEN4JTiKeQK9gA0yS4mVpwcQQ90eat/6cxOsyUfzcvjQ7b6SRRAXOyJZlApkrpivDLDY
9HuUI2t0RjHYHOJ7Wpfy7fEbUcy69USzcFqlRlSm619Tszi7ILNATp35mNIoEGpnf58b+waQcQRG
Fk0yPtowb7jTClmZ3ZIbbU5J33YNtDaUYynws7ofgPzN47XyssgkacZzetEMzNaTz9ASy8NbZMrm
D1Z+JP2YcPvPlEcrcsTSGNQUnhRJSWMBjFz88vBYXu0kgcHCbszBvbOwqj4xl1Vpv7i1TScqvYmG
SqfjFhFPxuCQiAsQIVRCewklmDB4BH06PlzWygZaOLTO1uc8lr59FrbsJQ2ov7/KAVJ5UmvaHVT2
sMZ8AEFKww8Av3cCnl7ahMe5xVxccr0fF6PvsJXkdGARzuzRWrs8hU/bOdfYBEInsFo2jNoaZSMo
vRcJvafI8QR0VJnt6YsCAPtqzEnl9Kw8JsX/TCxtI6XwIIUCgnG0REczsuNxbGhy80X/ZMSokCk+
Qj7zFA7M3JiQ5ZSxp4PZ90jtmXmyGyyiAnXTHRKSykWFmpIH0y+Lf3jysp1swcFKM3LNEfR8qGWY
68boX/kTDTrEjJK3EiYh5QoVH0yuUdr9cOK8nEas9mHgbeurjEKlmuqCQzCovKuUvnfOhD/OTjpH
Uw52GqsEQOrjFvQK85ogveNSIb0NE3+JODQmpVxyrtAm01Kgz0bLHxUJNU53GfJ7Y57XZi+FVwRB
XsxPSPh6tMq3D12EOM/DYY0SF+K1YTUgiYrYgZgOrbGiCyMrLH30RLa3mQ6JPlEhj5wBO+mdWMZc
Lqrz96fGjkJmt4ne9gIjgAcVR7ZYCT8MHz2Nv08QBzT3Sl6JMy0+kgF9GpXNCuXrQVSiTd/Triun
VqPP8MXQmnvO05I82v/+N/UBerH0K1FXvmlBT47fbUna7/gHR/csu+59TI35481ELEUPaEZhh+6U
idZ5qK1hLJ19O85ge8jw8ytO40QUlC7O4q1V3h3p/Fy7sCmwVWkPdjxLm4+bkEc9ZgS7XZ5UsCBi
6kVTMWC6siuoCo2sygu4DMcUtNrkc2tG65AN76ArGYIYXZoq0Po56g1dL6EfQlS075B65oJ5x3YT
i9IHTsAzxJJKeJ2bDjGSyNnsw4k2jD6waJnj7rLs/8D4ah5rnHIFogJ2WBKnrU38tggJhht56cx+
yeCt8qz5kv61SMETHfVhpHWy8fpg8CrIhzI46WTShzmGFaN3arzMeuCaitB45dZVwr9gg/KtCyr5
i6smk5DIThaZg9AjDMI/lNEYk92cevshGZrMNhB21ipC0SxWILbVXYEUJ4c8n+2GN5MJ1OJGJ8PG
q8+C99hTJXm2dAYD2MuQislasX8m9dVIuJYxgRuxm8JaW7yiCJxk9RKz19MaEFIaurQE44+xni6p
Sf6wB1SIo9bd5hy03HwWL90GMAywlm9atCWeWIFbfXLznuQuC9gCPBp0jEd/8QCYYT78XUYvwunc
VSVE5z/g4qBzG4/jxr3/vLn8GEhQEWw2ahuZUlnPaOJySyL23cVBaqj3SSwZMGnqluoQWEAKU0tw
a4tuga2WXl9Q9dArQN+bNnqNt9NwAZ3JQNmq7LE2Y6zW7Ssr8WtY2ehmOc/OccvJyarHLp0y2XxD
0bao0oeblNk91Gee4x4NCDUkbJHRCazz07IN51HEw5kEOgLqVqsJE99C+jonIrM4QeKXNlCP8htm
J9kVj+IYF3jnLANlpsyt9MR0UlIsRER5zn4Kkqfj7O8NBs8Yqm3GE9R8QR2s
`protect end_protected
