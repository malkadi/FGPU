../../../../../RTL/rd_cache_fifo.vhd