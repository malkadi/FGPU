`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
cQDd3XIPPlgRDhqULvYHvwCty2ZrVwzfefmANvx1dZIylIMC/SlAcj88wfYJOEUSOPC1U3p3rRJH
cF/G+RPdfg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
hcwXqOGXIKp1yMXglvtwKNDD2csTguI/218BbAfP1Qe5YaY7t7J14bh3PN4/sY8v5SUfs5PPhYYF
AVoQ7+Y8KyIAkFOjVjl8Q3cizlaMAyaX6UCc4wmflvCCOjy7mkT0VJKPELyiFH5OE1gTiKu4NfqY
cLpas2QiSAVn/xZw83g=

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
JJiSVarYWytdLFzHp3wkrD5+jxEb6zxCxwIxMuHES7X4vO/81ppoMZmSB67P59pBX5Chyu0EswKT
bCRha6XDZljqkcBWrrqj3cLRE57UCaEr1RVpDNBMw7hjNrwCb9eTELEwb3X0mZPKBqVrRNroBMN5
Mb9o7SPJ2GKhIDEDF5Q=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
x9rjekK3vn0E248BFQkRU8rm2REs1XV6NiMfscimCVnt3moe1QOgVJzTLPCcPYvThLcZJXwVyFUX
J1k2lVxuHKaC3FNNToKLX7girUcVANbS6jS2AjaAfdpYmQXF6epSjXy+KOWM7AfrGv2r7XNIcV6T
P4He3ZDDIABlWanBaDiVD6NYtB9SspFXaifjJ2faT9Et8gWmYJogYQ4BjXl960BUcxWS5faBudWm
MidcfsfVFpzH5bJ9L+thBkdIh/P3Rjr9ssCSzEagp+1l0DsZGX583KqMaKiaZiIsR+KyQ8Hrld0H
vh5k+kh3k9z7ewkJNwM0LCpa2Y0qGSJOxIauzg==

`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
bMGW+/GNxe7XIGxZQsPwYg9NhBUySelE4d3DawPwcsMkcAefxMJ1JdlslSvSp+VjxIobQhkauqfs
plGQEEjRkhr+3m8iz7uiwT6s+TtBZQ509t+m12KAHsziCshi0m7JEPgqnpkYUxS5ZbKQCRgudms0
J1TIIpIIdBJiHjiJWPFKhl2FSk46olekE0MQ/LvS36IE6UC8sP+H2MLZpAxpzqHuZ9TNFvVcyr9C
pc7viw1i7pElJF0USsLWRjDFrkLdXdznJwKPhjmDvq2WWhH0UZss4B7FZEDrUrjB/HO8EjVy2Hj1
fpw3eQ84VC/StEBHWhh2/ovbE1xsoAsXeBE8Tw==

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
pp8HZNaXt/evJqKzoiOa8A1cmkUh/1mQf/2Vkpam3N+hCoX7wAAqGU/zZVMPYP16RpMjeC5zeSin
YvUeVcdgv5x+e+joKUcjexTi2LwQorDqPIl0bCwYx4LccUexnWG6I9/pSM85Q6QNP03F3dTfZ+nY
q8I48HLVTNxhG5xD9+JTBp8D7rjXe9TJGi+hVikOsYhuY2PrwtvuAWhuicAfJnsIE23LJrp0i1cL
6oyVsfKsx+68L6qOWniySUGZ5yDe5zDF3WoQ1oHIZl8/tfnTJcGPsIRyeo3fpk/6/w5zWnz1pHuZ
HvGPaU9zIF3KNoE/3qKTDNhAcVbvP4+ohJfKxw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 69472)
`protect data_block
nXe51dT9MNW1tnj96BZVcZiRAr+xmqUYgYv3L9IGG/LJTocQzRj11ryTuh6Xk9p9pyCm0SzteE/p
yK5PPeK3Jeg5iBUTG2N8pd9v2pORD/MIPWjolcAfLQPmyAOOaeFKuoX9qDgEC/9ngUJj4JIwEjRb
E/PK3khKeH9KizCbnQ3K9x56IGWYWAlERKNDMEl8DquopVWUVAYGvXSTD4X8qZQrKzmzDg0Jg3vG
9SC7nnuJcQDjwlH2fwIrv6xu+ftUS5j+zVUKHIjQFSpdvuKu9U7Bu5N10u+fczdNye1eS9xqD/8K
VdR02aR8jkveTHDAHzO9fS8Fc/loYyZGAZ/YfLhKjHVhGty8uxNUuM6VF/xE2Bp0sBi1QY5XaJsx
qlx7hetVFX6JO1D+eiTfb3L8rXzF89szVD17Od/GZqz2+wqLAFBJ0YEBWF3bD+xNm7XUIey280XH
UibDYuaBwp9uBHgEhfmKAn1U9ic0eXZMwUAZMc+z3CXe/GXxSLyKTglHTFcfMmtVJDgWZv1KTQ/L
fBWYvZA+eTV36bw4XUEP/ghgZBXnrMKxEOMvkoRlRiQw4bNHjJoirICn2L92RylGNXOxDc2Zd6VZ
s2R7hkjNMWIPGsiOSUg9/7cjnE9gBlBIyR6i/PtWmgtSwlwkQ8DdS1m2e+avqAPFCx/OGpq+LYMW
Nz2NTxKE+9+QWDEGt+r+TMqGOv5vL2e5VKRKAdPYIqCn17tdM1xfcA2mu1FkBP/uKCtllke4gr51
t+z82jz9j6JLIa6dnJYPxsz1699X78cgAZb0QR43fT96v5w1Hd/4p6H5XVyXo7nSDJQ8mZ5wqCFP
xIYvQtc0lQD2WxLbhXAYBmadUDsgKz9q8t7CgifiddX6kiyMSDBs/n3905HtdtYGzTcJAi6K3oQG
zQS2NMiAlAHpPK6+LZEvhTUXvrmofvED/+QYp5ddwJyYrvNRfIwAkj00DUCkqig34vq9QfQcImBY
PZFaTwUB6afcMG49EHGatrAvh3egwe/0BHKA4EfTNH9i8vJEwZ7q+Yj/zGpYHtvur7RxsBUp81gI
1Bm85I8H/a80GDMx8E/egFKD0qs8/iqOSqWEaif4C0fZiHlnB/bHFLLddg4cVOmm4UgYGvg63/N7
+bGVrMbBX0JK8iiM3yQbR5FXzFz5Ka/akB+jKJ5M6LM+PtxT0vTz0qtQN26OlFBDd1PNPrSWgjMo
VJmrmUlGBwffd8vSlUYd/PoTxHMLJ+B69gTDw/1t/oO0ARdyqIJvjkE/I05AxqNVKvGKN/r4cl10
1H5HPDjTxUH2YXLMxx2a9SA39wCXncC7+DeEPqGesWrNDEwSdKtYpKIeV9kcfX1EwaRN48V/uFln
hsAluutZIlFBxozY0NQ7Efv9+48Stm1Hssnct0B+zHaYDiS2uNeDwTYIYXjPgmoHhbcz33Tk0a+Y
R2PEiwkH5T3jP67MkJS3BzouCQu7tdrN3OX+zlu6juFLyPmvz6LLueKCyKbW3N66X02MPvWhhZah
wyecxsuPZfabr9g8wo7Ur/hSZ0FhwJsHCTaPysl908D0ySa1FVL0YVzb4TqYPTbXmfyEALNyP+jR
9gFqYe4GKwyb+b2HudSwEHxHn6TP4GEKAe3UxP/XaQaS4gDjwZX2OCpGrrXwgilenlllGc6d3yB5
XLyYEUprYGIol/M+9lfsUjqAwRSQNfx7UTnOV2xFdQm/2AJ/WYpwcQBS46ogXzw3MGgpF8LH0tKZ
9XP91gkcIeBcKaD3aQQPH6DQfCgik8HJxqlyvDXKxcA5tCDp68LcASSlyzUzWIxGKTDyldc+UVRn
vbIpN2JYwkinR5fdOZ08kvo6eTmooOHp5KVus6/DthmS1kQ2lbrijtNYVG1Qlo1bBVc7crt8+pwG
TI0jACj1P1HT/qTbHGARDJnLqa79dZ6ccYK2ICKIjZwWlcRf1/Odw4vq8MI5qqFdSMDzAHaJR8aB
LUgPtLtjcuMJffLWdJSdkgRH8WUSgkqYeEa6Ms3Uko0RBpCLVWksZxBFfTH59XMxSSHOLrg0vs3F
sicz3kvXaRHZgwyKcKQe2udwrME9I7H5pJ4Q31faP7rdCrBCrJ4bIkVlSUULMiKpuZA+hQGAcqv7
OEuEn8GpilMIdnYsAuDZa243s1ocbGyNn43q5tIAF0+L3ZeqecH1T/VVk9cIZrV9Dy3loMJ/3C7q
tmTsgdCuP+tBHEKZsp5HzWdKrUsGCcw8BxebHkL++4VFDC9+e4emUYXpi8OMmqwZ8yemtw6/PF94
PjyTxcyJleEMh/ltYmx2USbe+STBKIxkQROEXbaDh7MX1HMD/URWL2fCcqitywHEfMLQiEsRWDZA
eXyPcuo36mO4Z6Nt7mI0+1czysde3M7SAsNroQfzlLkQpdWCF30JHbCyM+Za236p/s1drcvUFnxj
eofYvc+NdgNzSuvjM2EPKCLQlda7k9N3DU0yGzs2+6wKg1j6eE3AWRf9Al3A1pOrpxIDIHkk/+t9
ck/PR7j6l9E8Rv64x034bZBfd4wS1tO9wo8GUEulzJIqPX1AhTOHx15DsQdESdEnGJjrIaEIDkzV
h/riKmut4DC3Qb+SAbLNxivc4d+HCDTdx5FXPGb4XGo6gMomuBk6jDY+dx45h+ZsxAnVSicicYhc
UJ4EqfZhIx1Ig3kl7LsrhQbr1tOLLGdU2UWnl1I07pnGSU1D7zU1xZ2VLN8cjPKCo4OLCAsdkupn
0+0niw0bFSumLsU3ZlxxatGjr/hUkhBy0JPk5Y1QUIFPgc0bnRGQkW7J/LnomI3vJtSVcatxJ/QZ
ttJa1qRosAbApI7gCYgewW1pI5VTPYk5TYV/Dz8ry5izyPUwjAerXMig34zpv5dR94i2fBUur6N3
kZt1BS2wiadyr5CgHr9OCND53xBvRDzh0UhM8LgkH7SLHi0jQiUmJ3Nml05oeXhm2y3oy1rlV2ie
X4R7XJXsonsmAXqThaHSARdL3km0O/jRuCmK33+LRAHx2cZNVZRs/QwwaxeF/vAbhb8HOtsuTmrx
fC8yn0t5PhRSqApOFu9gpNLcMOki6W66HhIR0Xam7roTJRtdsfFSeRcUY26FYbhDn0/q8T7XIdyJ
II1/AS0vIYI71BC9DHriZdjFSlYK15e2XiP5XCFLkM0jy3rwmUz1A1T2f7M76Kc/3eCpWxqNAAzE
/BRqY97MUyGLkFyB3fhvr4gVY2hcx8GpmxvrrzjTRQQViWUwc8+krBV+WuLwttVL8oUOQu+Tyk6L
XtVO2dSA6N9jfCNi9oAFSDbfaFnoe5lb4f3xY/gulSRdVtu/HJKyoWepS9VwaXYeYXzjBzsWMVHd
RX5o/N9py1jBw619QzKCZEUpvsrsRBZwm/550OsxjCM11M1Kn6KgoXu2DCA9v8wWvnBaYYC+3pHk
Tbi2MuEeGPbGwvGKNDHIPmL9A/yeqw0kjKWoSA/P4cu3BDh9a0J3b44gsQLl9AXmUhC+HGEFodGR
OhRnhakI3BE4xNE7inAu2cTsJ9lMVD5vcC+27TFP+MGHThSMngNG+YdjnGVhKiwWr3D1fHWhiAdP
skX+LxvbOPGgubQCXteURtsnXuJ9KQJVmwYl7DVtZzJ9QNdNwcejmAcUpUMp7t+3HeSZhQBavVZI
DvNU7k44K6Rhpyw+IkclWyBdWR0Ht+DkHwLSwpYxLOGne7uXQbjc6Jo3pbujRCh8f7lXO3YcqUfX
r0GQRNCahHNaO1a5z3X+HCuGM68BNlh8p9Phvsn/BoCJpt3E3aCuSVL/0Z4ogQnibNWMGJ5aHw2w
JMpCiBg4OP4A6wRuhknb6VfaXxIKEO/XlKQsYWXLCOuBv+vBtsoNpS2NAzXWAj2yxDdWtJZl4YEc
+J9urFZhB6MQRTi7i36pgTOwKZnECglF1Now+T5dMNtJ2AeO9lLCf3taw65Fw+GhDT24LJZykwyi
iO10VxP3ipM4725sj2ZVzGv3LCg8oZU6B+g+qQttovp/4k0G71ESf7ZWpOXDz1HUDw3hFtD1Kib5
kCKw7DIdduzyG2B7gTBRo4SQjQ5X8RE+d1DDqETJ8QXtyp8RurfHmDfLdJL5LpMnqH/fFcgjoKxt
WPoJWwEOim7tO1bT0n0oV3ISOggm2tG11Bjuin+iuD1JBDlG9zttSTbegrHsHbOGsBwGQKXSD+7t
uxQ3wsnqBPJz0vcn1wX8oJS6SQ0n34cdUEXtWe6/XX5BV+cUDsHN14p9vJW/s/qEPmXf0M5hrKFw
IDfUVits9DdkVmkpNyJi3XbqXmDNHhcnLg27jJI8zxPoax3nIPhiYBajiev5WcT1Pcb6NkZVrgCg
9sCb5C332Pb0bt3yvbpaZswYDzhNNBxzXHT/NZ70sx7lDHIv9INAdy2Qzl7CoR8UY1TZk4qMl5IH
V3jdHUzRmCFCMg6fd4IUlGdBSom7wdKr3mnobroAP7EpPuHn71yPLjmbIgrSlHLrzYNz+7ec19PE
/YXQr4wHubciOh1+WScFzoEDsNpRf6HpsSLWfSQGOHY2Pq481Jh5YgajEeBx8xQ88MPTjMQkybfq
NnaxcG2MMiNF7ze9Il0pnfMNtyQBsKRN+mYBSvbwTX4/hoNOkGSEoskPWwnhaTM1hFc3nyY2SY2G
Kp0jXSeK1pRO0cqwpG9EFkjYy1d1je4K2BruftiOcLaM+m0RD6yBZu78eEM3A6WXY6CwdYBky0JG
l6b3GJPvdY3tGgTBHJ1BOzpRAIw5zjZ2Y+P2iCDDU6Ekzj6H1ttUNSMydshRh7jRRajpkUTUuC/7
NlXrmHVOUUMRuRhIRyXY8NjrKvftaMNfquclsLrniskpc3CiGM0HI5yM/bxoXv+m5/B9ka1LwXFt
96BZmhaoDbhoZDYgz39umKreix8TxtUHnERGd2FKpEzbM8PGWHPUNB3TfCjqbcYNucpH+p0S0Jaz
dwXqAAzUN/eQR5ftqAXkS0o2vFavFVpiKcwbO85HV3SzFS1GUNhnhHqpLVEoPPyPo8alEDl0GDc5
NDHVK1Qa8VnR3ChC0xyBqk0jWln1LoTtQHvOV6s4383zdYn0CB/KOmK6bHJng+xYE+e8JIsHrSa0
lIhnPWNyJ06EXHc+4A1aJIhy4QnVVHwLNAstbHbioaPVSBJW0D8JTgACAso+egHXD9OU1sgBINHG
jl94Vv8h1bdvvGsK4SvtIrKH096GtmtxbdI8ftvuCnSm02deyIxXBCp8IdSDWffHu4TH8XkBISNC
IM6N3uFOi1MMLPkkERGSyyY1QUH5+Z2d6oSQd78tiMHMNBCY1DodbV5JWkqy7tCTycxCKYeNxS/Q
NU8fqrEVaY5VIcuHlevDVaqwM49ef+YBvZtmRBDNpN6T0QFGe0/HTLi1s/82jHKO372AMtKE6I2n
teZnsUtAAiioofu2sCCKpjqfiGuzfdQuHGFhhuOLdVxCWgXHjAZNRQiLtbEnu+uiOPhFkBADgxiC
/eZfxZxR8Un/6gu1h1M1oJ7maay0z+tXwU9TsU4VWJY7DXEfCVwlVSbYhL29Pk590d200Rv593lb
I66eK5+qr1JcZAW0wkpkjrHqDXBz+3Oqpjf3tH/Q7LkpvxbRqsqxIp/33JoyI/s8NeQquotX3Osa
DmD50A3iqobxhXyiUorOOJMVFAS8e4JS3CTN+2eoyLTRRq+TG7XbZUTRrmtl0YeAcf1EoKm+zsEq
29nsfYVGQ40N7o9Sjl6/bw1kIrGoqBzC7e30f1BjtcN44tVBKHNTScjTL4AMZ2ctZp5saejlh4YF
4VffKMTEy1Pc9IqHvg37n5nGZSJTeeP0RAICvfi/Kxwp8bshyviTj2EWw+p+dZc5hxWLpEqa4XK4
wdxl9KRgSg9sfOqZ0hPEdvef2Haw8721X8HBwbJsv43MwibpIF+ZBf/R8G/Cwz5S7prkSrgIxWI5
sqsApzv3l/Ng83ISNp+vfHu5bK/gumazRARm041lqDxtRYNM36vuzblflrfvOoBEt/L/enRAFCC1
RtUnpapkw9ffkh9pf0MMOiyMnY3DyvW/hfv2Pt0+iK+Ei3WtXXnQSkYlwG+3mGoky2ZHpU2pgwob
VJtWI2DdmA1LNuXlB6moZj12sg7hUcEZGgNPS0Gjl1pjYbSnzbO10/s34xK8t98YU/Q0kjMDXw8I
vSOYx+yjXX9+jYc0iYo+BiZdYCsPQiZUqVfdbR31LWBuVWl7JCuVPi2ni67bMmifU09shX+wFHCw
V+n9677zEJeGtqIAOOfMPFokouc5dWsZst5JohMU7g04x8kSBINxKhtWQ7h6rEv67UZ+urwT7dwF
ZDJfjhclE5NJSW8FbBg0b3QvsrAKQJygg4dST+YlCagWWxpfD+Qop6sOYfIjnjeL3Bze6KZxhk5S
L8uUSHjFUEyQMbc3elMsxC+HFesy9YmfwvIuqLDmamUxyKXQe81C1bmT8wdfgIU9b3T2FsGUXWJa
uPuAJ7+ZQGX0xcInuHP4dof/46MDPKWq2hF5bt8GuRTFkkWqUG8sB3y9v7JLXY/mELx1pzperI1n
VjGyaCNVwpAdvhsRW9+OPGb+4QJLN4B4/TfOjUT/5FWBaRcY+jRoVb1Hic7dMJa9D6pODN8Ew3b5
f7l1pFJ49Ov8ucV7zj6M5WQ3XxzTWv5FJ8wkq++GK5qG2kFbbFAhQjSoSWUds+FUvyhjNW9OyaWV
hInn1HIR2xYskruNIOMN37BYKIuNd44DDsJ0Xd9rvWUHV/aZUzzk1BrV1go1YEchmcpnD+yYs1Pg
5n2SSN498D1I3L8DTUhieFsoT55yxCVQ4gORoY1p0NM8tHfzv2sYXPL21dOlZaK82K6gVYlzELYo
lb13LRKqv3Snz/JtTNWGT5jMwUYsEEQT5hUbxSq90qBpaoToFWocUR/z3ZaW8YgSv28XpIrDEkSb
EGQigVQ7XI2+qmApTMCFBtjf3ytQHK0ppjBa5+iC8DQ4SbnTMXd5R1h7AT2BJy9ghIhoHPtwEXZq
zEsCAzJ3sNXLq68y42orX86HPX74O8x1WL5f145rwMZZtjQ4KUlcG6kbxW2ak7p9jwsN+WEYXvss
5He7nCJ1tOqCTXvr1AR951TKtuURbv7673afUcEOlxLaSYeHgeAVLLKBBYi7QQvhy/n4jq3eat4R
EWnwNKETWp5wFFLtoP6NXwPdqvU0ZTshrqIshQS0xxCXW2w31/qdAkkDdvFEAXwtggPpphJWs8I7
0+0maBMuBAlwkDHycGs50iYEGjDxvmR83uM47I6GsUfVGtHaSCSfFvXP9salx5yeb48MeQx51+GY
X8vIB/NorBo2ukrqyPwlwXBpRQDG15pPfnGuHwhQe9D4dE7/8JowPE4XYS6QsN6uFYPorNoTyhNe
phhJhpQJh3VBSINulZV6ZZ5KuE1gCcZKXO3aGArXQTeJaYfUso1FuSV3tx9iPppBvee5k912bsRn
HqIdBl2Nz5ilcHc4hfO0jEwNPC/02lifeyJuPcnsv33ntdFd3DjPO/JHT0ymIT0GV9ATWGgzsZaw
RYaHLyS18kl570SjC4APZHA+cg5hSD2qZ2AnRlO6c8GnBEdW0M0HDmXYcNHBWoQHP79Ga7t2+8hk
H+IvZ8QM8b0K84q2/bJ50bvcyzR9V1Fy6A7UgYhp38cveVk6kKyk8mq6T8oFyoeDXUSzjUGo9WHl
ByTAojIlPPN6IvFmvhYWDYGwTDojMfPIjC5rUJAp9v7/iu6nf9JJpUe0M77JR/hS48J6lqxOo2H9
ciCmfFTiH3veFIEQGAGH6W83THNZ9Ug3pMczMAWuYBFecwCEucmOjG+3xDYhKqBCR9NyMq6fHlVu
RgbA0dtVmpMmgepY7dmUKBD5gWMYH0dRJ1IPf/5EK/0LqGSRnnCddurSd24V/QemxR7IRD/uYoho
AwDaEegZHAy+im6zo2Uxz1wjQ+de37aDhVRXxeiHVSGqVQitBzJT9KgfkGA7+jN1415k6kbcTtSB
KWAIuAMC7MYWR8NFlefdTc4GYSsFrSzHkKmKKbeEvXwomsPqyiRu3BpzKav6suF35TqtE8REnLY0
Gy9Z1arcKL+yai1r3O7U5BlH2CQh9R7b+wBRpdwMO5IC65p4FeAOKIwha9nhq5stAsyP3QyKM6F2
nvq6Zmp5j58k3BroNvW7dvEWSO3Sge0cFKpO+e2uzHwbQAW6wEh+tWc8kUHhzklnxpBxBk7Q8w9k
F9ihZF1X6GQ+uiN0fL4ChEYeyl7ZTG0giIBfGH58ttXPZSXvNdDdsisVexHZHLzGOsoQ59yUDAd/
wYf1oi4eaa5GsQY8VF42rivaKZXmnfATSfcqXmvQkIVfakUSFYHEH6VQ6Ai7BlpcofJjYBe/KuJg
8zH5iTNBc3j7RBIDOd773059eY+oLEwN5mdOS9JbRRpQWe+HYtVyQIDpspWKZihrJwpgxEYNAja8
mDJ9KjWMvEI3R2f9ysYswPKa3wrE3KSsXnff6TvvyJZiEylHPVa6Qk+yWDtJ55i0F+MV875ALpok
Sv25uZGSFoZ7i+LDYNjQ3GfJCo0k7u6AxSYZsQXYEqltU70dknL0xyF1FY8O2FfPJe48AlLO32ZY
9UXjtziy4NFJIb1ZWYjJiGedRuuYshvdpBNNILzR1HbQuNbcczvCn5Iw3S/PEhiVDB2eoxyB3KPd
pXK+8UDQboZhLkldT0q5Mmuk6QG7w2CCbJXSyD1Z63KirrLxgaTmK92J8GwDB1xW1VcNm/nr4BrU
kgbSWZvAn53ORkYZCXAMNSCzWBs79Ve9G4XRr1hvj8F4M2bWPTdeeJT4D9DmqdWC4herDc6eon/S
OP/1MAWJCwr4fHIiqB2P7/6twnBl+NcrcOMiktiVBCvbHc2YFR7cSVT8jSr45Bo6W/hOPmOYgJII
hdNgZIazXBART72nWnJtm/ZgWzNroAsVILCNzJCXWeUwFIq7tHiqzqNYGjLa46LioqcirSn0awb5
L33dDgndN6Ivxorc8gosG4r5K/0ZqEHlEG9USNP6AJFh9SIaViFHYeRt7UANPdhjpiht5g97ZUTx
VNPA/sA633ZKafz7V8FN9UrWuYbq97A7RLM0TYSAze1I3259PJnXu/d8AIX1Vx8G0ryytBQJbynQ
vb01XnJxAVGhbXDTafahJ/T8sZ+ZJOomwa8O5e/qJnLBZgTvryK4xdUry7yFy8yxV2etEbDQDrSA
k2ZiZhte5kFrkBVO8Ybv+WsIfCc+4rV8pEgrd49X7Xk9LUh9Rf/A1C+xmb8l6ZfBII/MQ3QOPhUb
7pUsvPKY/ZF4DQjUiRPgKDaAfcmdOpvHIWN83Fh1FU+4MmciI0THnls1VG8hTJxFSglI56b7jSus
Ooss06Ylgp9ks/QsTZpkIuVNv9DMRlyHpkzXjjGMA94aGw5BT8Ylk5ih2QHRfx2mYWovWphg0V2J
pxK63YZger0KFMD+NEIuJHz38WqmaXjRryClpmXhX0WKw77c1CDW31m+HsZHzWk7F2q7IdWI9hp5
Aj67Jf5eiRqGe/f2WTfnde6DvBfR8rSxjwN7he5yU762rYbC1wRWU3L1HfYmfKicr9fim4TGskfZ
SmDfv9mIictnm38/2wJ27G1b1ZHdCPVH5DNGlgpusBsU5/dUrQXAedlh+uOWjGpPjpI/TXsWGPyg
AK0bHqTNdltu/q4YkbHziZKaPycNvdJaOcsXcyC6xErQay8yejE2n9afToo0tDynJayd+DwBcq4K
9YqZOcTNCqnOuBqs7gR5KIPSmfR9ZwYhZo0qiw5Zb2iEmlb3AXxOhSk2n/kPnVxfBHxmo+21ddBj
0E92aBwqiLsTZhkTAZv01uAGvMFvfya6OMmXuX312HVgL+J/HEGHHe0N15dAZk9S0SbeDYlOO0aL
PJVbm00lT+hq/cPxz4TtmmdzClYB1iaYqrlXDFZLNNF2kupAAhK50WXfdsPtVHYCBLGbjEMnwtIv
qNwMhtZyEHZS6FnqCA8CyJk4xn8v90YEmHm6fKoZMfF8yeBiR2hpq/JAkE/KBzwOL66ijiJQWPQX
n0yA105XXk6EakcYbbfw0Kah2aHGfo3GkJFHDoIDdryLRigRAxw1jHIOLbS2BNrTj4eJhtlyCiVj
vH6WfKET2krwILXWRuSKTeOR9KwUbJXK/9mcHDbXJ5J1RxhgDWRvC7HW7xNUPOaHOjkTELKOzHEw
JU/PgjJZG9b7hVQMAnqHj3QoS85jWqN8YMjl2ssaaGz+idmuLRji41Dk642TaHQ3ixs5siK4pI9R
NPCaurjA6Fi8w0O84VDPbBTPV2yoG8fH2deQ71Icj+mLqZAKSdJGo/cq7bNf3AeBIBfCna7aj+cD
RCBsi+8Tb4pgmtK9FlLqE8drd+3q32w+qACy8jsURzLkme6qVguw1fY6m5hYqjnhoO8IJjGtpnb0
SBn2cmLP4GfjH4RM7jWOIignJr3v6mCqXbJggJZUXn145G87vGlMHmq2w1QtFFm9w/i7hmttfW7d
0unyA+yuDXKTqgTX5PuaB4t/jMKFmYkmbFta4G2STI36iQNWMMXelpoocICalJIHCTeaCphQ+Dag
jC/QlK3ZXko8fEsHp7dgDiOfrHRFvzvuyLhyS76jXHI8PY896exJMU0OCsGQMJkFo7ILQeM2jC1L
vPdU+vHV0cPYmFv+7Z1G5iOeEgdALZmVBzhAWwomQnk7rUAaOwOBXQz95PXno9sbdIxHjxG4gc1t
SpFGzO6kCZswRzMg5k2oOOup3ldxx4B9hfhrGoOLHkO9KAofXHYcqnRhjf6w8xx6L5GXP28/expG
h2JUSQEJWU8ZUu+TSffqWKZYGqDaBy6/M6h6yCjYfDpzJKrwR1+jqCFBvj37M6dQ2F31e72hShuG
tVqmCdxKu1o+lM2uw9tCPS75WLx+WLZdZ1WcPwS7aChQsbB+ZcpMNTNeSJCEkA2hjrm2WQY79Bw6
OO7xzi3FHfuouMrX6yZZIAftAD9r5wswzgWgQ15JGb4Q8OCMA+EPdVXnyVK1puaF392n0sLE8ZgF
DfePNb0R/iG4lv/xroUteog5KWF60OCMjHHaalVD6UtLXGs6o78wCS0nKCRRqkp4hQQ2d82vNTvC
JUsMq+mMgc/+1s/ddemT0nMoKXICAPAfL8K0m4IhHj4ah4b0E6Kmass8fq40bMpmFPujJ5xvu0ti
6xxGVdfJ/LiwdiKyNMfW2cdKjcKtWUr3HQOBvYjl1GuQ9vEg8lipp/RWVGDmqNKTHLI22MePz3Jw
k/ZrMlwAbcLHHhe3lfAkHGPGzirVESB8AwBczMOeu1e4Q6UCe293QWpk3mmDnHaGLNKEC5aEpyzE
rmqR+pyx9icysBJh4NBn4zd4rdXh9acP8+UwtE2g0eSLqHnVLPOoV9rSN4uq/lAQ9PHRdnqPdFHY
RjwHC8tMDZXegnZLFybleaSGrFXCu1dKaS0SVeYHKM9RqDyRFQORQo5S9kLMwixXNlMpbO+YYjaK
3T4Jht1DJ+11xPJzun30O+QhfSv/7p0txkKkVceLcoVrCA7dPVWzkvshKl5SPYovUFEIirt4nWY3
Q0gDb9D5wSwnXiDhhvd2IMNFSUUey2sAT0vpWaH+4zIcVd5lpPYHxlXv3CrJ8deHqhUPOxsfpOTM
d0HobmIJwtFifNgHCvqytdZ+/bRbG2bA+rXId35UhXiN789dD9+H4kwPFcx92fq8i/7ru1DkpHqQ
j59Abw/1Eicn+kRl3cVbTAsZN+y49dpwZWcCpCHxGThkfYcG+9cuvhDXTqdwm6vxBEed017Wclrj
J3K1NI0iqQ45A7d1jkoymYcoqxap4qpHw13yboBTZ/zajtEGMBFdh3yYWNfGkXqNPgjhwVbOd/dg
7RliMWN2lMCTNxCy9L0zwhWF/yVZxwpWC9jUDKt6uHAPsViKB3bpxciVS2p2xC+uynWEKJ5Ju304
nOpeXTjWucRHqAX2jXWG/R9dhR5Ab+a1Lshdj1IBG680uxSlNYPdyByhP7BbpfUeN9M9Gw30iDT7
6vXhmqytxqZvhbNQ2A+ZPv1jAUZMOEXeNGVo1XIxU+d14NkUwZv9+g6oAm1Nu+TK5fb21ZEotF47
rqzctRSk3BFJbBrkMKn76hudkjDadUpzPiyu4GVXTz5HDQEwFP04gBrBy+mwU5hjfaIlO9K3Y7Zk
oGmhXRfdLsmayKxhvUN/K9fzNWm8eT/INUjLwcCE9fdLcroNIEXRVOZN2173D1WCcRPFjZVQHC2Z
k4+gfiLZKEx9RpnFSWlQ/GngpeDSvQMdUBAlPWsBgl9lRi3HXE0RofwsnUR9OxRDug6SuAK2jcvi
pga0NftT8PdU//ePzj/R4o5sPdZDFkFrAoG1CxwhrPOG+zRRpWKdb45GejR4z9g1lGam7g9sqc2V
KADbvAR8NepdTCKI7NMMsWpaCfbXQceysqvxw0uipdqtlMn+5309lbbkX/EN1I55xhNqufA5cUg2
Oka6bWmAeHMz1EZo3y/9BnjMvVirGNo8Hd1BBW4F0LBWtVZUi9Uym3EE26DZ6TnlOpAPCqBarTj+
MhaardmTeW1QgYUO9cdOMNrT7+qUsziMBaLoBCm9BTKGPXDZeAaKpYmCm9p5ZONi5J9mhS5mU67g
7QHCPEEHmNXXH+86AYzLZ8fB2dEqn+Dx8MGFeOXhP7MRQwyQPOSUWEbZglXwBM3b4CN9t0RZBRYK
jUrFAptpcfynYmFHUH3z8u/HBGKtNsytlGNPWFjUsOv5jwP/UaO1DTcAPagFx9YUAMN48S49UuZo
TeK07LL94Xpt+qTTi/JMcksdl1hJSkb/zzG7IEsIQayzNdXDZgBKipBRQXalSSblsBFHR4gSCQkz
K2MTNzrythZzoPH2AGSr7hxaTAWXKTDpAvqeiQCG1ApsXZtV8pY3aETA8J2oPrUbr0BLe3VAc860
cmBRqMIaDwYwnswU7JxVYAjYbo6FjLRQ28PQRJg2o5ESEgcdD3psnvessl6ngV4Suw68X9QmtLPK
+JJlxeuHlBgZYyVuC2nizH9D/GDvmT4JLM6oFJsCp9y5mwIf/pd9JPrmstb5ijeB4YVqX0O0+bRn
bz6wnMqwrSmvzDG5rUP/wNt6LdC0o+HCQERSVKC7wYdns5/T22wpIq/HZcg2QZNQLyNM7ghJC/a+
lg9sVcb04h6sSa02L9aTJ4hFJYghnXsJJtgHJMWsJrSiWWATbuI/4ftt8/qwUXJ0YEVNIp/zGSDI
xrRX2+J1UmUgA0XNjyfQAO9nPCcZ1KTky4xH3JpxzAiT+gJyjgHzbneQkW1//wExEpveXzBCZwOf
mbtsL1yInI3aEyNk5Ed0nhYwHcY9IxDQA5vh4fJZQr5/7btMGShygE28z4uPvP0fmV1iTGIOpXlM
/3D9yVzw/BDgr9mtYMOB/+PgrI2o94WPAwBrCMWIIC4Qx2SZEmpiEthl928p1qCHVeDVFRxxOZEQ
OzsoZM6tM1vNRBAco+35/BReXPQMS9sbn+7EJ5HD0B1HuPZeXeSrwdsIFqg9X6Jd8tf7k34I3cA4
K99pOAEjbHKV2pjF2oOSRwUvgbZeIlDLxqQcLFTOloLGADdf6mZaZV6BfJxDUYqsH4npRsfcIMGR
zph5G9IQtuB2SOLHuZKNha9Vc7Ph0Bec0QrtPGgUbEMUdW+QXBC5NpS0BeWpXSUMRyFzc4buBJCe
0pdOP0jCViaNMt3j0868+OR2ix1lpUgJ0UER41MkIFkdkr1+fNv1OoLO2U0vQSrZ2TC462OrVVTW
0WzpRuL0d4MoWgroZ0TrJfLaqVGqS07S0aXBP0IrXl6GfaGQoKsoUYmgejY7hEllYUfMXtF5rbmO
jRUtkbRgluLZa49XMutOLh1u1o/58dKB0mImCXhcZ/yXj6GNemC7YQyGXwY8Dhn8IiqDO8xWBfju
V0AUj4VmsdqcH5sZvTaUrSfgPEGvaaMw/p79skz5F9faAXk1fRdNfpHeAivDfy9OYUD/KIhQ3p3o
z5DjLTgCBkYcNY0bYDqitbvRwoPqnjafnTynpnA2Om4uK5ItLegd3AVZGwTiHrqXMtkj8LyrUuJF
TA8X+ToKgFaGNhmbasFxW2NTsy6ZbB1yzs+EDGyt67vRso75fwwH0QS6+CDC1cROlWVylFhee0Xt
DDTmo45DU/+T6qOEpB9kfK81TyMhNgBLRvSW9gZKT649QSfPwpLGjlcvcmri/337EvHL0+OrOBDq
ifIIhb0IqiYrWWS81kMsUVorvROY3BoBVAe7j8tewVlNe1WgkZGd867uFep2FS6yPWXauywX0DNY
o+UjBLoAvUUVQFlNWq6nHREGRloUfq23p/skPqmIX+J3l3oXIT5vrg251ia9f0VejK5pVB039pQi
cAexqQHxTiorZVXAlQ7D8LqTxNcPjtd8XGAc+XogC4mEhGPcAYJsFTNJPfbIPglaIiVBPbF+Vr9K
oa774UIbi1pGWPRbVFkOZZl3qpX8YX8YDA2lkVGxamFCwttDMoJ0ie5I+3PYLaeUEfpmD5If9qgJ
fyjjo7ej0MzLHKan9wYSioAuaOfauOlzGlkQxKBbZe1ojbwoEVY6+YBIbm+DhCSuF4Ip+qZr0f9y
aJOy4qXSsNhLAKEnIWgUWFJz/kR/c9YqEQ5ZDCmYnoUHy1PvL8EiTIpHJrcpG6oOtgQdRqRLLb3D
+/pCkH3b8ro6PsZKOlBV0AMLZJszBcX4+py5gdXhOcJxclkanTpuWy5d1JRhvjkkw+vHciTLWyva
lCwWVWzurQ0m5h2cnWX428HH331d8qUuHNlWFKTpANF7d6jvcxe6lEQRIOORnvi1k5aSiZZDt0JB
eyPXFvoDBvDrk6SnnHuAPoIOE8aSAsF7P+IXvhbxBBww+gckIAS+c3wAjkRZh4Xmg/XOwI/DUBhJ
paVsADzWXk+A3xgy/OdtkKY2QeE2arqqftd0AcIqWSjU5x/uv4Ns88gyKcljjIfO+LH4VLGSlTad
1ZcxS/TackLr8KYAGPF6T6AZzS5MRkQX+toQS8J3M62pmbdwPWj+Qo9270cuCBUcwSKi4A9bAWqM
jpfSuvWeELIpbFaeLTSIylY9xtVoIPXMLvIJYpWSczcBbVGg8f9ojJQcuF3MNUycZIEpmRD/CK0P
YjwFWIB6nDBaQZfS2Nr0NiMXJEsIEz+3iUFSt7m4Jo1vVZrd4tvpNZpb83mj0ZirLcGmioVx4Hcj
ca/bJKSt/jnySYZJXXH3HixRCROqt5wF3T1KRK3PbtkLQInMc6mnJtFqalmhufnSICm1Y/HDFC68
rMu1NRhSw65kS3LAnsD4zvCJuqoT4WxcmgfSfUcc70fpqTDwb0scBOIJGsF8W5UPBh+k+tixZncw
HEJ+B8Qd8geXgUAd/TSDB3tPSGedNvTcPbgPpsialJSk/pE8cxRLObBewWZ9HTgY5gIIAU403bV/
UuLXsaZcua4r8QluxZABSnNAz5KUtBOqedtT4+Mas11Tl1UeZsOpvKBgNV5gHuoM8Fp+Rv6wZK50
ONbLgrRIcKsNX454LndJx5OSlYrJakA++9CDDPSd+kPh9V/TBM8HNzFayDrsAT7+U3o5V91XX8Fh
ZrjRM6Yioss+YBVFTnUc1eSsQhu7tX7QWfBMHpxunkv/y1X+d0hibeTR8FqKsKLMqe3hOCaiB2TJ
l9WX10K7icJhNPAt0EvJCIaFw6VrmU65f7LIPNI32uqUpciSuFaGEppc0Chl+efA1Pw0oHYN5gOZ
7jsQdcvFr9xrWS0PJJgF55ngwsz1Ir/cHWyf+kDMxDdcXoWIJSvu2II6JYlFAkVOSMgq0E8zOB8c
Wsw4RhBi5rhPfqowC9Z1FCS4augOb0LFftjSYtWfajwwI6x6w8oyc/fe1OLqEaJBz8uj+OpXaqaF
YHf9ctQo7w1/ZiC+AScxqyeI1SadG8wsm/80o3UxxJO0rPmUGSyiMajWxyukKo5IPQbV0IqhxehB
a82fcoL0kSgBKrPZhmHzA/kdCo4qCyUo5cNH+otQtjuR/vl8OatHwyrIaCneoBt8usYqpyJmXEfm
gSkzf/vVTBZVHdLcCQXeaNqd7diBvUQ7VerOuV6f+d/i4pNJ5mH8EJdEwXMFmPCsBxdS1rrz0ixA
+pkTaNv2LC0vm2znAgKNngkff8xxMZoUdBO2Yp2FbLRpUX66ueIu4JhcpZPyvVnc8QO6TU/5ONWy
k1AI4Q3slS82yPTj1czuk/063fYLWw7mNPrlFgQBaLCmE1jP3hDzi6Pn0JxpafcqBVeSvHn9cIIL
kLjeqcm1vuvl37i3tLqDpDF4LPpXyr030ok0knKgYoFqkrguHOinzz76+3b5i/OmHYi6e5Bbi/FM
bafb9mZYEEUs8uLdGDbxXcKHjgn3qofVIyRL9OBg4gHjW7D3hKZGXHOVYVLVmw2XWbDSdffrcldK
fgXV/LoINok/MZ99DJG5pbSGb8zoL2quVqjFPwBh5fVsxtY/KNNzhbNZMiyDSgbg9OMshUmrPIYA
zfqGL8cCmnW+uazmQA8UQn6BdShR9Ij6NnVZNzg76XQMwU5YXeCI6nPkW4fErzsjUSAqeEKX4IkS
8u1+7ddi8eYnqvNQY8PaAQ7Xw0d6HfFFnhaBVwtqBg3CY4uPD0x+ZFkjNNNWNGqo4MKoHAv9ZkGy
pcaqy/mYLEr2S2kB6H3TMZa9XKNzqDZCKyjNYtfMlXrMvgbiWa849G7He4jn6WP3Exa8tswWqt6R
pM0gqZbRVGyh8kGUTXcyuYqqiwrcAcUI06rfeVM2uER9dtckoGMTsWDmGGHxSQZa9Wej9V36DJ8h
8hRrjm5jxMqq8/YF/iQWaFRm13nFac/peXSsf3WmGMPEishr6XkbrnKiB2CAUddmmHiPE9FSTc7r
jlmEen885GK9b1yw8dOyRqisNzao7ovKBHroK2J+ctFEFwX3/FFuR0ZgaXjK8tNnVls1udfWHAvS
aRAfhOFQmaf85H3eyaLoWKr2umb8a1ooLqXp2Cn+33QtR9+QEnsCPtfT8aC7AaYGLfMnFinVDbT5
aN9Etxk3TAsZXcQ80mbP318VeIetZl4u9lUegU/6i9XqrPN/jN2cBJBKHdxucziFZWHSeUoympJy
3RF9epxIX1Yu+1OYvj3xZcMG4fMg0Oh4Qmy4RH0sGMpE+uB2yxHFMvfPmFWDpaTM8OxE7+jTUOqz
xAYlYUPIlwSkgQ5p02nUg4CTN5/8WzIQzPJh0fpyukDSlJLq6jjVUwvHyKAO6vAF9sANjD5ZVlLY
Pfm/e6fCX4uxEXTCmMi0XVBf5gm3hTOpu97YVRZykt74n6SFBzGleX3MLVW7xJYFrxoGKgGCSLXz
2u0u4M8pAhGLoVoWzOn4KxwhgsqyFI5Dq3uPGXnEDKIwrd94LYOQMHXZUd93/V1t8yaMF6OyUf5J
X6FhVLgTvbRoc3IVT0gEnZT4kj9jjO3vfqWgsWIJ3aibJnwUzxeKE0b4nFyKniXJvLWHN83KJSLX
2XsntuuNr9Qo9FDbQdW3Tvb2XqrfRtefjVogcML6KJNY+ozxqK5ZxjMWK7EkUEcp/hITJDy80Nto
mX8DZBIJ7yfFyMTy34iAzIdhtMzc/2Y1JNuLm+ZbWBWzDNyvNJMMW1Y8wSwD7XXrqWt/7iK9GYkv
giOnIiRTuAznSlH+zFA6duSmCyy3X51YHeQLfDQ/mDrHvaA3VnYfjFXyVzMZc5vpS1lWkyi9WIKc
2nXnwkgMbzguuxfUGUgIA/W0+oo5FKXnXeEX9pbzfRkyo4LjrNzrLvkv09BtnuJfoXbU6WQ2zAOL
g6gfMpCHUpSg00oltqfcY/pDFDfi+/44FOollWVmbYsaVzSPHj0t5WQWqFfNrEpwC5WsFBaVCrna
pQNR5litN9onKQgATZvt5yCHSsO6rp0cHComIm+N0V5aQGiakPYTewSBXTyS9r8gj7afFqReIENB
k28/wUNi0oyqThqYaq1EKgp77yCCpnqg2PJpoN0vW+osSFRQYZovFop7BrcF46swPNqM1/VZg+6V
uMEAXxp5zLamRP6NshqDNrO1RWibR1OnNFLJVUCpAD0dJFMs21kyX/SJG8vH2Jt9hxvcbMkw+RzF
KxV5+1Ivh1hmwcb/SfghfqPXYpb8bECUEE1vOMmXiEN1AZ/6v4f4NvRkQQot7OrJl7pV/WN91jbO
nOWPDetNwYENcX/p2fg8pjE55Xx4v8vjDbXCMyX3/TMmueZWQjMzu++elyJxQh6PjaTilOAfKvYU
zyMjGuowLkFPwMN6CnAtLvkHLgmddxEvaHZWdzmt+iyn30cIxLJTvPNpEDYXRFvdrHvkWP4pOs40
vzp3ZJEOWSDoC3nQWVRwL9ldKRSB4kVD3BMkIhGGV/xtfe26Ir5qtPnVj/ddNA92UbKpmQqLQhPg
4O3Qgqomz8rSNclzNuGrAhlvVe4/gSKzOYRy6lgVFjK8FlbCk0BeLnwGfL77KmQUTcHKuDxcyMn1
sWTsa4XargGP5CLKVUEw9eg+SfiMbALuihVGZmhimIQFMXqLV9cDhQ88HTPopS5aEexyqQM546A0
aITZuIS2DRh4qz5aqdleQ2fFHtjNkrliU1udi//LK71BWhbUVwFJ/7VoW9VfwjcATHzwCclNmuC4
+jmfIo1U+ccRwm07u/JStwBNSnDQljTg0e1kIDg/DSNBJO/8LmeZqLO0KN1/BVP1GvreZsFw/IoS
Em2k9glo9k8Luwrztg83Tr67Qp/pcAaDqMUj0OmSfCv9M7ySbMLc5y+s8RP0nGv552jQ2QY7jfhG
qnJ3hdRhPsOAI35yIJFmvVqAnBkT/746WhHm9YaPwrllFWq2JRPyZcw66k4p8/HUAKXe7ndBwJSn
hf3zVnlEJD/L5Xz35E9lKfDpIyBvnEPoKqm7xitDDiHPXHUktWmzWvrX/oBX7L3LbV+MItETrmNs
iYxvFNmoMw7KFr7lXjqYJZNYfQNV7vvgYt03DIDHivuoTRD+bSWAMdi1l40CsHB96hxiilF0+ej/
kfUF2WnuAu1MuGU4bnR1fskPZgc+Lauf8vzQmKqVVfg+VVyF1HfTW/DDE5fZMPHC9jQ7qUEQl0RY
qebvVZqkl+ecI9i6CNbE6DpGqGbvB23X7ZkqcC/zWRkSAZaERti7A15FwAMq6ifOOI6SaIa09KnM
iElUeSANTA6dcvA6NdSIpE+Yv0VjmQRIxUxKK1EEeUCdtZQmuyyYcNOtWKHpzEzoGwA4p/JGtmvc
Uei6UGAp9EB6vmeUeI2j8UWu00RGBtuizCzvDu9vccaZxiiGsktb904wXOk8r7zrdCLwd+nlcmVp
Ec97eZX0nC4Eoxn4Wpt3I+tANOMkKDE1ugQGX69H6pbwoyhMXQPyB4akhrrgExK6EShQ/rmz57Ma
EZwxUvxFkWuDU3rOQvBUnwUPPMfiCy/wGqOMEhL253JG9OABte/NXLBwMLa4tqnJ2fPSkIcF5MRv
+6i9/GxZRORSp2JMbCgZ8Q2tRT/UeMXBuciwFsTcy3R7PvB7kJLy+V6p/pfJqoYlMzg6CZWDMuQ5
P8OpQJk/8yyHtoe3TsRkwVviTgQ8A+tuQJkLJQZ9aQOv7Vqwoqs6yifSQeZSNDuzB1ZIhY6+VKfc
HkmbqkvCxfFGdByGv38m1kbAUtXwiQ5UhP+MdwoMpHMPkR6YWuchTXE9WRBwKVu8AfnsVmAp7E28
5SwLLejrREVUvcUZH8EkEh+O3LHI00EWU+c3kbTxK7NzJK21esVlKJPaXFt+EFeX90EaY3XzFkEL
J/TMnB4uz3B2rB9auii/s4r88Da22AqiN6wThfmAvYVuHjFR3ShLe6mSR1NKDfpER6xpkd8LhDl7
YpQlrS0zA6IXeDdFh2Ahkh2IAlHBhoS3nYmdmOMah8tjqdgbVu+DzKmASleuqLe8Rqc2TsGgKAJr
0yRs2UFBh3CIZWAa5PjxUIYRUoYhnuGNpc0aCMoohPKFIVWgfaobSKB+wTdiq8E/cXr/1YILW8zW
7gaSXEe9c1BoUBUfkVkWyIIaBwnKkPAqyy71ZCf/Vp3pbEhqpJcTJVmcOfY1/RuxKRmGSysfhoHB
Gf9qvSNN1ZIF5SG/hNoc4QCQ/ab4J78jzH4TJCNtt46DNrvpncvDRNK5s4sJyLEHPZok8MRfxCQU
tUU/AarnFc6xEFYT7wMb/qAoIxYtoHd7xzBSKSqEHXlnLjG6tsv5WM3/VlNXoha+16Z/J2ggO68U
b7EzIoBPRhaWeczBG3axyJ5z8ghAF61MinWlxHiIAEEtUHyXmPBg+SAhyy9LOMz+gSe9SWdFvc++
JpfZLIjsCADPeaezYyXI1lulgAxnoLUV/bUWtpNe3WhX2oqqsG8uAtIZAMiYjEjhUhB7dZsH/7lS
Accs3ZK5FKPKrXm1vvuDt8w+uuQ7hzQiYDlx97QB8PtNKSD7mnfiiLtiWitD8+MxoNnhm+K0HoHB
Nivg68m5i6FLrMdqd2qOOM0jeqsDXg6k7Slz5RB+M1AYqw98dEvV5oKfwHx7eNunOYEIUJSbjKsY
/HR2S6C1hnkxlALXOLXhfVUDaIWKIGVB0PrZaqkr+Ev1uHwIpio3N831pAMs131hGtKBO6L15bOv
48TTLodDbXs8b7sBFt3lMYd189jGQL9P98az7LVyjlWjm60Xdkf38irnNN3Lb3kAoZeV/23eIdpk
kW7HJNs9hMT1oeigx4Ma7TCf0jLRjjVTQE+64AO2C/Mwi9cJ10VO1nzLUlnXFqxNe3elKdSpxOzE
9GB7gwL8EoGZifuI0+va65pW6F+qR/2RV/tmxeUJDUuFTj53gzHiqpOtHKEExpVQXMpTo+mjox3T
KrknGFM2rrqX6SaZXGOB9cvnJmDGuv2WcG2WsOK7l9oDwJ/H7QT9JSfO9GgsNiyuhyKd+3QwPktZ
TB/U6Hwe6+Sm8s/Gu09qN8P1Yp2mRwp4pHksEyAH/MYNlRdTg3dqfjskEHFTeDRwDto7DO0wgZRZ
2g1FZJidlBcIUtkF/xpZ4pTugDi12+DRKNxXF+dDIn8gsSHsvXi1ZbONTl5coGDtvUVRU0gnUvmV
ueqO/Gm9AFQLIOhBzLHMTqKxxqBHzVtifXAJdmoLY65nsk9AWR7WEJ4likuDsAjYJa8PO+Ijq0QW
RwvwbWJjUNLnOXwZ5mlKqtB+QrK02CFQTmctuC84ebhtnwMdrt22exhcJA34foq/m7PJx+WH+l75
PCUA/A3lzDoCAmAxKwWWhXT1HHEUjJwRn+UAmK8ZpO1Ij/f3oTlGbrYl3zE2p84qBsNGV5VN7Zug
pw+HkPV+k1ttfHHdfgDMGOcJ/v14xitmwe7rHryo1OeKfLBWsFLTqsSw54vEfi5iJ1NMXoZMF/6/
M1EWP1+cVz0l6qWqo6FEvCQgu+XqA3Ix/35q1WuCoq8UJjesmcI7MZMkWEAgaQT53dCYVs9g0K0x
RDAqn9lAg/mE8mYsHMP32w6HaLFWTgK4NC69/07aOZI215ZX7wIsG/80npk+Z2nDooS6fwMrmO82
tUBUQlRZByTbb/o1F3QjPzYjRJTu+yW4s6YCp2G+UgRVkKmDXyS37/+1i6MpndOxHf7/ZNFNhHWD
e2bf+pu5XcqwC5CE5DhTmVU8UvKCl3JCpOiZNHJDf2BYSHBW9+YBcNZv+hckTBc35FsIjFMfSSOA
XMFAiqATZWWopCqpj50lq8MRwh0Y6cTyeS41w4NfMsUh5gEEqkrHHIv3LRqsFyqe8I+jU+gZjFxY
0s3Lcxhktt6mSeJqcsgOKv590jt+sxLsQ3A6cFK6BeBZb9o0iwOdCbG34HQq7H+Jfbm/jI7eczAR
8Ux0Ly1DgzwlO6X7imBo3RED3Rkch5EMraWKG954qUBGSxVlw1UHWoirhYC+VhiQTZBqL1Q1wXCn
pVVii5XwkCqxsK3QwyoEnZTnuc862ac5RmWn1Wi1L2B42t1doVT+DOkLoChg72mVqjS0Voqe6Msx
xmUUtZUZ4PjwpYJywhDTv/UK24uyc8fuk8hVNUOowd3BRDhLtVhaBPBXrUtYvG/m+ZoJD/z0PGeC
O6J+yWoX83AXFxV/+SGQBdoD6eAiwLOni3WeHwZlFEi3SFRKXndDhg8k+Rp65PKhcJBfXS5vF2mQ
1Oa57C/hoiBLGxZJ60NnyhvageNMnxKMYXduE5Xl5x5Dk4WeHbfqHiWTJ5YBoXgDTNC0CHD7/ho2
44IwRa4q16xOISDyvUQHbEWSZccHPx/u3JR9pexvUbbKGOPyNybPRCuJCaBLb7fw5jFfwOTyVg7x
DFd7g80Z1n0IEcOCD362/xuSH/9SNO1ZxdoV+7QkKb/b+Z4TCPYkNBpONp1CbvdOqYFFd+WRPkq/
Ln4D0XtlGrqfBxzCRw9WTujAr187lZJaZhSkJRNo9sZu283IgzLSY0Wdw/s3kHBOJLhgAuqHDmcU
aCZkn7w95pjig7JWLSfm2YULHKSlNxxg/mswSJqlVONnreJyfvJ1i81kZcQ/QW/oU3jmYL1oko10
ZODFdt9Axx5PUE1AWvjWEhjUY5WH73Aadz51aFOGnHkvIt7bRg5Iv8wUKvlXeOSMEicnNVvspAdR
47kHI7gIYo4jZRvrPsGIebf12UI2nFcbU11VraAevBUtsZOOnUptWvSe0CvGQg4LsBaLmxL8GJev
Bfxl0KGdnp+Ut3Dsdy1gDJzYobutNPInZhILW52jkO5yrsHi7cEJD7Ib+2welC1m+XCd/DGMzlyf
yeZuQBAOA6T2Xg9rArj0p9L5Nliu5TeH4gWNO6I+mDIujtlzYy17VT6ndDZ6pR3e10/Q61DBDXWg
SFojqSib7Fww8a2jFP56Y+71HlcRTk7LP/QIUiFvG4zCRTn/9NViAYq/qxyaw3/lDQAJNIGwSO2m
tZhygRcot099s6asFXuBRSSSpouisXRkt5FYIzi+3rgtM3EJZoq3WKsYSwGqXZKUd0ZC45zxroBn
8X5NKsEwjlkq9OP3FG/RwKhbEUR0Llbg7AchbkKw7qUcbAb4Pc+MWFBgb5/RS0+DN/0Z4xXj8lgo
3UnFqn97RL2i3yLN5/FtDKDhKTxLFjp52XbG+OgoM8trW6kQvP0K75vQHMs+QvvmClqy9dChDKCb
1P9aOTsvtm+RL0g8N3k+pubWEUfk4BYngpXI57EGYXpkRZZhC4RPcobBbQqMFieQ+8j16zENwIes
Lvt5l3XraZom+SOQBXYjl1ldWJ7ERVNZ0CGpOKSi5ewyfMpMg18utkoWH0mkTS3O5qCLRFU6i8dC
h2xkl95U4T4MzXpfcE95TplaSZjqqQhf1924qXOw1ckJoEOb8noEH7Q3I+wQoWSMmg8Ixyuf0zRX
IcOqu1BJUHtRLk+vNbwIYtPgL/mkxtPmwYCIw5yN7ZkL1ehfQYuuGVwFRRgVhluJ0FNnpeUP23WH
q1HHC5pnn6o16Jjx5AGeaMxJLDhVMtu+yHXUCkleGjAkhMk9qtOjr6LYqZzJW/QxcPP2sxR0t0Bc
Bt84e3z80KDl5khOItmfNVcnwsa0IJxugGZeqTLLhHbluPpoi7HVQemRuxFDb+YxCb0n7iEjUK1C
aJFJ/e4ZExFyxrmvqoFNtRw5Cmig/Q0cNHG0d3DgzjHp095WEdJCGmy3wTNoS7gGgtmqFI/5ISEj
3jSpnFD1NxjyFuLNOeU1OP5ZDh22eIJtoDk9wOFJYU+/5GeQgLOTBTUbMU2hc1wYWWenHgoXiGl/
Vq9YITZwQ4WM2WnhzKp9A15VeA9wceqGB7C5JabzbrPWCS+C8BLoRyWA6oBUcVOA8jXcbapz1OjY
iuaQCjhBA8n82qb06D2M3a74EtXHHC+TKcEiMzM+hUsSipQNTE1zCidzJiFXmsPKbuX2YhvOFDbw
9UUlydKccLKU2NhjiRzOiT76upPBRE+uk69akCOJkYTa3id1VhiuHhzbYGZbA/lE1+SiwFSHrFMz
PoFAYi9R7Gx4S3XNUFbZjzQvPZHryvOSnaWC6d3xlX7lyBa/gIFy6I+lKqXBmLP4kJJjDpeokX01
bS9TUPswvpAbN5nA27zsH98zTfyt+Agf2XOS8noWxywsc46c4Bb6QnLOItFmhHBkC8MM5vfPSOCo
4yCrePRuWpNmMTgCKbNm0zsuTrn4wK0nCmpUa0isZ8A/CFCUzOgpTwXg1gtkuWScZwQ/xNnu5mU8
PWjseprP377TQMoZJ9hT0x3s7jGxEYrX7xMJVjDQRdNZiVvl+Pc76dWUYlLhvPYSxAMe/7iIQEys
ULeigJr4PJizjggGRGGmZ3R9qfuOdv2jaDxhxeRq742DAUUfZMW9pARsTC+Qm2pLx7FnDZm6N+vN
OAMnxOUBbwtNpcP8DNT4Kd2vWY6cEm4RcIU29nK9xqHCNIzo6f1OE3UfhBssYWfNkkLJ58BjWdql
TYCdzf8huHbd9PHw1SqOdy8z2ZymnCwpisZw1wVLNFpVgtWZYLmsWqbDsisnkzzoM0zZwMFTH5zr
0Cp5seujmxAImdjVbmSJUg0r0R6Q4yHAe8N4In61kfwzEEAxWFd50V5ZBl3y0qxeLDBKA91PORY2
ODu5dvXAiD0/TwN+D9KJNKd5gG6Csgr9retm8HRkbsrmjp7q+D85B2bbo8DD/dof6w5wvr/RBcna
RZAC5yNowqcA2MJe08SuOG7zDHmIntWbLKgs1MNRiykn83yuuGcH79H9HCSr9KyVuZcXPOnHYJRk
RmwIPxJM5AzX526txqbp/mKfy/ClPVhS8s8n82ET+KaeDfchlomY8+IDDWIL90ZqKf8hveBPQZ0P
y9GofNwyZ9RN9BoZwOXoNFhSU3+RU+kjdeeeFWBiAuOH7JJ3D8JN7v0S6xt6erZICfy6V6jUVGGs
ZwK3+qzsatKn/kWRb9uIKNRVnwLzEkf3mIXTGWvml3qlDre7+1SvQ9Vkh+sVT8gCegtXUUFo9b5n
iJG9/J5xe2dnRB0pikx3cp6gIeGQFi6HB18VIg2JfHOg13OxT27PlQBv27oS208dU3QsPpIVQ5+x
ah7Lj57+Rb06wEVq9zgxLNrKF55I5b+pj5YcqvZm8J1iy719AmaQZFRhcMB1ULezTl7lsWPDB/9/
1Kaotv+etWNYu8pKq34VJR5pWroY7ja8YC8D2jJSsnDCfsFTHYFItyGfwjm7XCoyeuCJdTM9bCKA
YBtX25ku50uaYGKTBy8Pkk9h/6sQdS7HtEfLg+VTOEWt5M0petv1IN7iCrCx5FEDGbZy6yUn2miU
sXsXStQocSafKM+7FX1VqbR0zvA9PXBQE3X3ROKi+RCTnYDOCWxGmh+HFiAM53U+AE4eDrBrBI3o
hwJbbcwpZmll5G6Nd5rwjXgRbyhjJ9rWCt93aIrBK8tJKRr+ue6/fm9Ktsb/V+Upp8UIyEGRTfx6
1OLj+IZX4CQ3xb0DkS/i45QgOWd5uF1wjfw3dN820bZtSdbTL7wQRnn6L3wYlCwAdkxKLK1RdJBb
rO+FcPCfcs7w/vprOGBd8+HfijvKsHufkzFTiNd1JzbvJFiTFu2Wz2t3uqnBiHGiplgGLU3hmuZU
NISZqRi8mmNLcggOp1gykAPL6kPgZuSmnChm9pnfTdwspZc7xIi6wj4xKtJydCro4QAiuQzVZkV5
dAumhi7lEC7zInpADY0q5NxUr8ksNFf6SKGX08KoWzfRViRbObLpU/QdBt5lMx6nJ1nsBu54wigK
wcEGaVPPezkf19jRQQEawRBzyHNNXZ4Df+vxDpgTxyP0iNDRNyiPPT/8j/xSFHBXwTmjoTmgrcYD
R+sZMH6dZM0Va8LTZObZWhIpxprdwRED5WqovnTh0nknT1n7LteVEwld4hMtrZPo+GiuP3LPoiZu
q+aqKz0kfNqc7BFrZR9JA1uLntSik9WDCcIkOJP/hh8f5Jq9CJIN3G6GdtME/8/qkGAXWA0kRaiq
IKW9GhU0nTULglsAgnlc2hSx5LXgkrJH8B5ovXmVnhT/MZY+UKbs7inCHjh7/NudO1Jq/G6Zti5T
cFCknVWi9DixvN80kGGQA5UJ2iFv0kvbpbjQcKJzVjY++WBc0OGTQYHMAha+zyLXR+/PtRAov75D
Jmz6YkwaTjsDwUZ5xwafLVk9Pn8wQyjui0IL8DELZwDu0osy3aF9kmGYrWI3YjmVqYv4LTabi/6L
n6eR/RpgP6G9CD62Gxc9HebkVFfNOKRWgIHGp2Lz5ZFhBhPoWgSnI79Bzg7jye+3E/AINQW3GCbT
+wkHdZuGrG4VERRA6uJgcesp/vBMKMgGDi77zWXD9em60JMKX4yHaTnEOdSpPJfzh9Akl2vLt3yS
yRYKWKWTzobNK66xS+r97rbDcQGO0+Z7yDWbQpti7IFmwdDrDJyJwBnxDIEMT1fQj1IspBVcbyOA
L3aQZU2H4k9Zw/ff/oyIm+9Q93QPZl1OQORZMjyozohJiKfjpiPB7LEHnE0bc+AXTf/fkt+6OWl4
6Vim//Jhy1XRe6bGTih51GgbPMM5pC9D7zLJlynr3gC6oXGew+GRwO1t1SkM3CNoKFntyHBDLMTC
2nVctbWc/yPZ3evq3TNx8itOfTaeoq6447YFI4C95Vz8lDKouq+MFJm5ei6lu9AWHvy2fXOhbcRS
JHBHB4GwkfCk2ai9iEILy9MMRamXGR39MgRQRYS/oBbuzsqp7blHsZv1IHxYh8ApTUDU9Sgg6cQ8
uLPrvmGHpdNF/Fnzb21JD/6wshSwcKtqhhCADom10RcMVPuHc0kW3HFG/ye0flfmp3tLrSn44oMD
YjQl0GEPf4sx50HmbXK4PtCI5anyL/+L1R4ZpgBSPOkOo3/B9QEstdt0kcjbg7lONMHkHGJtKB7p
lcj2AA8g0MGprum4IZHF6SpLpNUZ3bl7RT+DtjM7RZxJPnVcmg9d2CCro75abNLOsIlKTzwlQjB2
2rivpKKUV4NBiqYywUbXk5FIr7giA33oW66diL/aGbjMXgfUCveEn8yX4K1HzZvdHodMMOgHKKgo
mVZy0wLxx5km/xeRkT+6yFGPSWTjJ768j1FFEqvDNEcEigllyzyK7uDPuIs+H+c6VOeW3WzbjKHQ
ipGRImkhSe8dFTSgP7SgExhXeG9k7oEQOEX9V+zrmGljhaO2K6hdOZ2V4vGccHEpLAtTXUj6J3Gn
Sa+zxJxlmmQoZ5jaFcPWTztdOdvF0vc9lVlAPWsqiNnLJBKG57HdkixoquEinsFDlhqJuyoQKN/b
ACmeWlWxEw3cAIuRTZBTcO1Krq9LT1cseHKr4J0Kyolm/OTjBWoXkawFXPtxPQqE66XpbORYXy89
4/KZErfHIL9+vRkVie6nGPkX0P1YMDjNsDx0MqmUfz4JRh/ESu7+UV3doGzK7j/ir+tgR8dmqf4h
xLnLpwEstWG8z5es6UB+S0/wcVmpvIbj2mqibQDrO0hSLI8HtBULejCnEroX1x21J3YqxcMp18md
w1vcQNinmR4LQuKyX1qcFs5TgY7SB/cJc2gP6PFzT+HasB4owo4wYcNUo0Vdz/tT0BWR2dw7m4eb
aSuKzXBrKWC5F5CrrYV/uSoYCs61+n9nuqtSUViwjedjuJ9MqsDDb6HRxVvUq8ofrSPFO0qJBQVO
TUjVlGFNwRMyY4oHiyR9JdhhIaU7Mq6Q5st3C4NSxM52tHZm/E0+rXj7qb5hUWriWoe6+RyBPr0U
uQh1D5DOp2vuKQaBdT6cmbiuMZDJD4i6wV7SWvXpXk7vu/qdbLt8Pfpo9BUk05K973GtT1JJ5Qp4
kWqGISs/5RPPR8PCewOni3BNoM0qlPquTZ2r0+bpXN9AxvpiJSD0YlmYAtGPClpYe0ETd0jlZNKk
21b9Gpx4Esb/8EkPOJ74GBlpmz/dlAxj7eTfgnNGyOoQghYVI0in3NuklQZHYCmttw1pEVvQqVmo
UrL9TIJZaqqzgytxVVc/Btcq02oNptJxdxjKe6nF8mgjQ84t+tj375fSMCQCSYC7MSP3m8KMpY6C
gKQT6gbiO9TV7O7RAwX8CHfudpOTlgJaqBLFLrheEKe2wqSvl/UNxiz0zWyO0u4t7PfIN862+UXN
Z0mPF85ZLceu2YWMTYsYxcOhyfPUOw61F4q59pV7Qz1ZXbPlKEEBgE1Eea0HvKDgtu0hiyjHSUla
c7B7p4ixAdf8v6OT09+mcmLEZbb/gRbEAOBrf5dAc87SemYAQRxYAsr5nHHlZXZJ7m/pqEzgo/2q
Fe8Q7lujJvPPqzuZY8A27FT5QfmzDRC5RXlqp8vzb8GYl2MpRw5EBWlBrLCXd2InDKn5H2JwnHOP
02LhpbpWBHbi/yWe6kD9AGurU+uRI4i9cF4PQWH2IxWtlTlh/JPqWnANvqY5Bf226cfw3aNGz61L
XDIBJ0eA2+PMtR2Uug1xP5sDsKqawqox1NJ0NApPv4CEwqn9rVOKBu33+0rDOaR7YHBXRNC8q44Q
qZqCce4J9GrXKCApLNtQAlbP8Z5XYtd/V+f0p2WVXgqZZgellc8PwxDCBtadTMje63K1bdRHaIkb
HVrjeEpPLzd5aK2HjnVMuYHSITxd3vfCFMSq8B9qNeegMBI0IM+SJcr6Gi5y15edYK1tdCDd9ntg
bh8hbTPC0k3iuBJXUiVHLBP3YgX8fZDuTLYEwgeOgEwHmvCliR4DCbud5CC5qR2VXCyFSrZc0ZI6
9r5Pz0ExfIk7f/lSXwGnMNm5CEpJHCuOQrJ1mNTTNrBV7IfCM8rLbk0l37YwN7a4JTXRSGfnnRPu
w2ywk7e75osAReDDE6Fw13jOA7ksNO0f6XI5vILW9qT1MruGpYAstCVAgQ2SVDhSLzrlTRSz04K/
0I91Sjg0mkQ4EMCUg9CosWeResoHZy//mBjIgwvqEFdOsOYlDNrJY3ke+szJZ5naNXFTQSG1ciwo
lCBFyw8HDymf9NNTJqjNmFtcqFQ46NvrcOKtkTrtlDdfZWQys4yX0Mg2hn37E7g931QKtP/y6F8T
ZdCQoOoyQIzIpCcJzcoXdT1byS4PuNQLjLq3bBoFrTi4uFEwiOV76uZ9YKatfr1BslJF7Ln4gIYA
9ncQQ6y6iEGaCoqMBKWu5w+xqN38VKc92FrYVLQmcfs9GqFvqRudabEIdZyBQz1ti3Q0Kv8mHLOV
nz12JUm+egrss+b0RIs3mn0MqwOYiFJ/3/coBf69ttW7+Qd8XbGtL7axm1bfps/kFNo+eZ3bX2+f
YDvUEHg6zWXb5SYE2EkwQJROl+fujQ1m2LI7+/r2I76cCfogKh06DotSfnTPDolxo9m48MqcbzRL
DR+35uEiMJN5qfMN+0KcHy+7tSm4G7j8xfRMUPDXwxiR/2kApuMW0wjox2fWHzJb1FeugWDhFZNg
oflsLakMCttlLE0/oKrCUMECIYbpv0ehfp3b9N+YeEby2763TluAzK5Y7TQ/nR4uwu1bf07bevnu
tFokpcK/WkOY6gW1G8tKeCMyLif9eYf9AOZgpRvI9Jsh06kK5lyhUhi5DrKErEbRR25M7ErVMmFg
00AmzhFlL0uLIGIB4oFhrXFm89bQLPzH9+aUVPFR3PanIzer5PM3jZiruK6E7z/cPujJWe12vTU8
vx9B2qJEEJyLLcd970jjnOgXZIVuNCmyi7dKwlY3nW0hUF/dph/beXfqs6b1bo8y06HIC+L0UH+u
VsUwuUixcoG+GoTThzYpuQL/GiK8qnvWrpyQZta4jDdcePQSDbePloUnQSqKZ4Dn5HeRWy4NPhfn
J+fe1J7TkWWpCgeckeD1YROmlyyhcC5y6YAnNY5BZjg3LFRG17u2NQGmIoB28JWhjDu2vf7Gskd/
fbty/CzQsbowZioVd3IQQ6WtoiY5X5b24CfN2FnXeOM0TTBUI2rUCncFG0Jq72RaggwkGJDzMXWN
rqwfgMoo8LE3T9MarXwUARYrYYOXpx07F4u9p0uq3Z05t8KhS34N+uGyG55SAlwDIjwGVZeVU7aP
Y0Rrz4JMtzBhmj6D3Q32AeqJ/Y+7TBKXrRr20OAAwmE/qAZanZL+9xsYOhBAiitVLfTxBpsgM+0b
DFyvO+lDIDmAKr+jN+IgvsZiEM2yVT6V3QZ9Law5aYbFtUEP9lMn74A6fGHtV9dUFTLLR7MIpANR
WEVSKmykrHjG8Iba2Q/xDsjA+MY0Wm1uu4OjqhBNnCNPHSLw4A7fTWjaIqgnx824/yWdrNic65m+
2xJBiKDS1JztvKxhN6JXUSt5sd21XFRGmeLvndC1H96TZAfT6PwDr7rVHf81KvjMbg9lQ2Ernm85
kefQE8akvsfVFuYHIDicjDxFMCLUdaTdhRbN5/f2YbdXLvw3j4VChAxBEH8IsqRqs/9/imcJ3dmI
/kZBLmO+u8yuMUBgT3T3bG9Qp5we7vtIniQ04Ld5jBN1cUcU3Y3+fGcMY0Kk7epOnD64jA0jb4gD
jIB02EvEsRuUB2Nu5/Eo+BkT1gkr+yXKSApfB5RhTgmK0jCTUQzBrCjRnIvNEUbLR/zVBra7VaL7
hfssZM/+E/87UdkVANCgzq6d0WEMsKQQjCv0ouItXWzL4MEshggszrQqamZIDYXDZ+8ZJ6Vfi7pB
Udrh1OMkqszR360EQfq4ZHtCerStepnrXvLZdKUHnQXDD/y7gpizK7AVr0HpemkWB0PGPkFX1zL3
S7CyDKLLXNK53weIB3ziUpce8EzKWLOyzpQEIyHYK5+iuAaT72xql8JNZODzSqdNb41JE0bcGmil
k2zGefjCFOVF7Byv/fJIZ4kCDUxW3UWG+9dpGRRS+h0NPMp1sm6oFUH3CoYgHIqH7IzaOAl6d06Z
Oc49jrAqY89jQW+Z49VEQS2cRlBkPBEqnawwwiUCEEL4eUEtE6JhpWY2jVcbzeN2ArS2hYlyVaIf
j1SKf8F0sy1zKthIdJLSaAZE6kIdgv0nxv2+3aNxffQo2vbfNkmcY0lNM7dhZz8yWN0KvJ7hJ86R
AQHroLgnK+42vmsaDWQOkoPy1+CuPkbQAC7cu1wp1XUApKlDtNrIe2ViOyAX23Q+r8YFquZ4OLNe
bSHcp5/zBNX8CzD7OdnHyW+kY7g24WCjtVTCM6tFoz0rJOnQ//xF0el1Rs7Ho/FfIHL7TBupaamu
tHKktr6sbT1+VgMeeyHdvQBjoz+a59XM/JAvDOrbW5wS35+LZK5sdYgpt0ssd16YB7aCoe8I0RzG
XGPFS8cDM1kwKnIqMSs4NHA4nboDFcCpzYDfMeA72k5B3hFQfg4gG1Qmqqe3bXheT+XHP3ZPx/I3
a7nRgR0gWf4MI/TrinY85iD6voUi6sNoA7RanPOXODrmd5GM7qI34D5pleG14MXdqJ/1My/9fVCe
MFc+vTMl1VJSRXLfl3WcMQi//7L9r6rt3fN5KYw9H88I68C+kNsFbycraT3BujaPdCWVsVbWLGcF
UMcNRJMEEF/q50CD4hlESTOvvrTW7W2BfL1opI6GAqaLyPYCqYjTf8Fl4ofRRvfX1fwtmz+2MZxw
u6SyxykiA0C6vezjKCggBkv2yZj4CSG5jSM3/grGoTF/33LwjMCFEZ1Ar1d582QOaBwElFWPzZkg
fFv85uEx67BkkVuK4ZrtPScVyqUHNWJUb6kMstMoO4Dq9NG9A074AlXvhpmEIII1dHCxgIisv6Px
T5XjGZF/BAdL21IinnDg1A0JydceQ7mn5OwlpDpdW3BlGyOV2Z2lHENKxg90b/PhYOyekYQvA0t4
LoMXDaHdHRvqBwKhCOobAG5hVm3HxT5kHBjX0ggimSYO0MEYUKbWTRLaSV1lx+WAIHtIEOODjeDA
Nf6aFyxJBPXNRISS28VP8xLTqs1g/YYAvZcB8f6FFbK/+R9hdRzJXmJqp0P4/3obEKtWM/OOqmjr
e7hRE0VkD3F6wMPOBaCn/HrYwHX5rpeJBVx+T6M6TMM7DclUhIA9IetwnZY1CA0PG4MuHDUSYOij
4MzgivbQaI88ZvjAQjyeiiZgRrY2PwKT7ooi/SxqVp3SaV3B8wiadHS2nB7xOA115Pv32+OyY/Mw
t62Ps1BYT7lKDCWB8lBkbo8sSW5Np1zGiPnn58GyPVPnhb8USXS/AO4fCadm2tWjT7zUZoz8Cset
+MAH9uiEVUme2gdaxCZQn7BupE8F9UEgOflfLEVZQ1X1J/sKhwrgxeK8x94CMruB8SYfz3NM2oKj
l89p/29jgisWJtmD0JVVUU+NnzaqP0IGl+tMMFn9uuOPHm2GXp2sCNiZm1CJ0/XmK3gPUq7Yp13/
OA7PYPiAdVVIaNLpYMFYYJ8QBOdq0A5OPQWQTbrsq5ICB3QbPYLBgrmZ+JL0tHrDO0UOMDERJblf
zIijSmSxqKyEluZ7Vq48SgzpjNWurlc3/vBjCIkcgJp8oD9UtpjKTutGmlCUV9iO7+5EILUZMG+B
dbqDwfq6K2jRB+jJC0y9x+cK/9vyWacNkwNIAZsNp7t17Io4chK++cM1w9W2xofINy4JD0yUIzG9
ReDTj4y2VpSW5rms3kDMGBm0AFENWAyrK92BmxcRHRtdA3wB/cFqeR+NAPIcilK+RAa3CPjKSvMf
zJ7ibm0sdCGrV7cUM4zaiFFF7lwL5OL92syetW7/IvSazEnIOjSp/d7/2CvRxvsHoycFywtu22V2
RHVfxB6gvZMN3T2Ymr9tDJO5j+DM7ZS9HfnN8+ATjG5NSmvhvhejSsZVfHlE7yam+nlvkpWnOj0i
7ngCWfhqBph0wuE6AVYnq+Vnb3EiOV7mzu0TwCLf1iYKOSbJrBvFEPHVoF3irCTZK+VvQMhH5hYq
1H5NiuLRAGuTScmkOpbH5Wl24ZluSbPWCSuzYyNBpQpbybT7l25v8bb6wYD/AFyzIZlAYef9pl9v
AUCvZZJuTfMRotUqrXUrXRBYbWo/iPE8/i38QVnAnbQWXf2CghMgiYxHA5IngaK7Cqg/QeTrWy9A
bcF/nHK/Z/XXSxAyaxNMya3SnRUutns589Hokw9RFsxZgF4QN0gMhs/aFvLNesm6ePivBV8K5+ou
s+yRvLundaXjT6dQtqNZDK6wTgQwZvj/abCZqkLy50+TnOYIr3ggVGeZQ2V3UF0WX12bfwUT4cDn
UiWw7tD6Z3mZq12qUlVJuFrVroz9olN/ycgj1LQV92PcGMSUI/n8R5GtW4O76+VZCq8VY2RJPHWj
g68yXzFCX5rh6UuSauimgQgMH2GmxPrUFUbeM6Bd/EN1tv1MmCfgM+ra+I0/jX/nM4LPoc0JrQYw
bQO5J+4Fz57gJjI/kiS9v+cqxPiLXRso0gszdAvVYfdgwB+pmBC5obSlxg1rh1FsggfS3jr/5Owk
gq+dGWiZRbFKTB5eZIYpLAgyq3AOZUjzpP9oO+AKuwRB4PVfBNjSOIwG5yQuepLbTfnqC9wADS/U
MAq/+Nv6fi3Uab0FRbjBKLyUIQICegDMiagBPGT8/Y01hrLXJoN2dQMlQFGf9nVbMpw28KNyBhCQ
ouIbPgOVUVklRwdhtfUWLR4iCl3izJrSYbph6EO15ZlgOQXNW6QJMbjP5Twq7/dhzvZxfWKyr0l+
yx8rkCdEtknZpKR3DPS+oT1zCH2ub8c6pw/GCzsTUSn/Phl9bSIowH64TdPQNwQO9UWbyuIdcEhL
YJps9SntBwhAlbuz4SWyPl7+Et0cVIiWoEQW50ocAiNEbsERjS7GBC1ZDJ00wwEKoVcTxGOHhiEv
brjHENsmMHVa2r/QbQAunf4D1e/g5hhXyckgnvCx8FyGeLWIIb5wiJvOmZtWqSHQecWdIy+4WOeJ
i/FZ6N/KCEjICZQ52D7WoDa/IQuUr1jkYLHBFgUXjZsP4SK/bI9OnmkgtnBFkLbAJiKmF+ez7iCl
qeSudmkPpy2Nqi023qGvdnU7eTQJxRYEfK/IdgcFeJPFGQCRLP+zYdvw27XN3J3fS7cK/s9nqH2s
QwdhxnS8EZqabGNrD42hSeUDd/YvOeS+VZZUduLPOU2ZxKRguFS6mL78CunlGrebSXLpGdehhZth
bAXmxeC/sAj2aK8ETDpu0VB5ZEjou3G1KIp/RxpYV6ckgzEFs04u6BjH3RB+0aKj3EKrzrccG3Bd
CVkH+N3VrfkTdqySQwmQ3axDVBG/Vvs+FEeGRUKxfiiWRuw9R2kwxVrPmYxFeAf/ZVNq2SUL2ut6
24OQ8SdwU0fKgTjGmc6/4qar1QSyI4qn2M00tIl/BjSHkr1hhUKyS7j0ittk1JJST7NdECSxNibu
kNwzXLIjiWKxxGahlyK8WiQl4JYTzyTtjaNrS9gg6K8umIIOoe2A8OGJNU9V9egWC23n5bM5hkAQ
pVnPUqVJboJOqcCM6CcD9bP6neupeB5ssRqA3ONmu3JC8rkAGaPB1HmaDfCdgYBAr5vDKGsaVb6c
Xrf21DIQVcMb+vlFFYMrYT3EP7LsU1YV5N7dPxlWKTAXM3eIFhptoOgQxV7c6ImRYRMdwO+5u2GU
7sFEZJJL01v4oZOsfoCyCVVROujSKgO56Y9SjekX81zJ817bplTXcfvCnBZzkSBKuAj7euoPRKTI
ZGLMFsM1k2GV52Rdkxd4+ipOpAwGAJ42hKyeOeXvWqcKHq6MhTdu/GOpZqv11xmQOpwmXlrHQ8ld
EpEdC8XLnZ7OBIz+MTfDVFa76mrzK5HSjzrRX/Ho4rulXSMYUGGw3yh99UKBPcvhBx8JHUDRkePe
Xyf5jWbefl0rbPSg/1aoSEqhcoSiqy9FpjZZSTkwaFVclz86vGLUFKxsa0Nw3mUT5iYCj197ArLY
3Re2IHnAntVuxVHMFAQrlcJ40AEibomsPZPLy/aHoLcGV9NXGESacnpZGQQguriogXC+G+AwiWcV
DUY6kYFVd0XnkK9QSz9x/9tJn5MswvJ0RSvHk8etwBcBKM7VoziStj9RhBVgZIPXaMX8JjkYwQO3
1p0Pm9cPkM3Sc4oE9lcjOJPM47OR+ID4PAKc2tJ4vRqC3TS+XpQe4YBjyMLeUGr/2Tp8QOSGDhzc
6z9NFW/ESU41euGPUzr3WP3Y/OZrbRXPK2eyQazudjimFsfkIihw6cPvYra2IBtNNZN561j2adwO
f8SeFxZobW9suIYle72MA+fUnhbNZ983JEvuqZXkskQ7FwkpNec78oVv8sj7YKWmYXiSJ+G3uIDp
naUCBIE/AQljBgG6s7Cqw51zQru9Al0sm4DT9Zcu/O0ktSCahJ6Dopbxh+wmLW6Yu8cBQW2XNtQ1
2jrzcuSLYsqZaP9E+kXR+iMhOGUZ8xPZ5/QuDZLif6+4YWq4jrqxXN7idg5oAcszE3hAQwvjJhxs
6B95mVLBQ1hhNv41c2wwH5T2R+o/kmTeKhIgvexEt5M6dDJVlWXPcRMP+1l8QIU45yoZR1RhPUKN
xtKDpZmCQuoyYfbRe6TEs5FJ1zLOeUfqPpApTH8V3KKUuvtWkPG6BinG7vxrb9MHsBuEfXz1N/Mq
4vc8X78yiPMo96xyST6h4CfyxDXMKEak0Pmz0AOSXRWSXa7exJipvg1/L6YUeroT4jUSJ2yOmAyk
yRhFeepVMRy734ZP7MqrefN2l1WJxZbgrMOiG/sDqYJljes0nJwtvCOd44fhkV/gFEl934lIRKtf
R5vglE8WzonHVA3mIrgeDVJQ30xotH2of3CMgCjmEwv4/iRep+2FRj4p8GnOEZmGQ55FW8YV9LFh
nrQKTrayBSvpCNb9fxf0T/weYzL7wKzmDnDJ7T7uQ8OljJ8JKW5z7xQHpP9K9mz4/x2f7wCOT3Uv
C+FWL9J0sHFCr5rTDVnATne8uwl7gt0xmwEHca2pXfiINlP4I/UtOoCOxnpHDb1V0DF7I+5eq0dU
+o94NBP6ViKFPJZrFn1mWUNtzhHAtj4LfJaxR5QrSCcMtCk9URhaonfY5RfDZ4DZ4zCdrHbxSjog
hC6fJBgLK3C/wW4PuWFoJRUvbhFCEuNliGqpmp526hYbweovE4oHoG2BQ1Q3gd/Z2OK/8oGzeCq0
9u7gC7UZTmYuSDLEwFtMjl76Vs0N+44B5uhrBj5XSCKyKzCi92ESTOKGBpL1RIqMz9WGDUkL13Jx
xvfBWfGtfwibdN58B9aWUw+itmNq47J0ERi8g2H9sppIXV7xzWEIlsbCyUnVzMgrLRX14htIkmEF
C8dPXyrfe+HsXFmfX3UrhReDgfDhqvZRvFaIzF5Tl+FaHRfClt0EiaOp0Rnr2QSxq3QNY9/E9nUQ
oI9cuAna7mnf1BTh8V6X6y2u9DfB81tRE0/azctTZQ+noy0rMPLWBa4muES0k5a/d9gD6JV6C2MX
RIg/K3qUP85kTt/n4plEaBTpQVe9M0Y8Vl6vYCTZS2H2U2kvgZ38PeZI6GMUtJRxBCmVuTdcAFvy
Re6T/jeSa8NjDSGG87+YtqR+RPpv2eyKdlSKi5+rvXtFGR7altfoX4dXiF3ZUJZWYRqpYhq57dSJ
FXwaEprtYhZ/PsMKEkUCS0dzZDQc6gsf6y0/9x3ZotpCVJL2b22mg/kFw0iZfmvkVoeDwtfzT6Cv
wRDZAONh9gs1rKJbY0P6wd8q2ZwHAPOfppEVvfPo2oZlBz7IrE9WZ+h1EeiDGeiJY2S9Jg6GiTE9
FdCGyREoV2lnI509sIbq7Qk6BDWuNFvN5EWcE+HpZytjZqmb33wOau4LwTdMnUQZSlxYAoG2T21u
ZtkOAow/Ht1ug1m921fjv/uPdXJaEaW+/aifDS86BYhw1/id35wUtefSBf08cFBaG9TELt1HzZ1F
la5Lm6A6Xwaybt5VhN6KGy6gybkFNHxy6afg+T8gRKhHGBoITWerR0Dpkbo6VvB8sOvP1XUkp7cP
pOcAr/wnQNIkCxTHQSb9R7BrLzVMnrlc6T8YhzPJyaIysF5Qq8tYBulObLx2yhkUkg/7F3xU74eJ
DSZUr1xkBt4bhLXwLpcYQvUu+RV6DmEvHZ5USF0ZeyXb4VTWQyRLghfHm+CGN3Ar4+tlZspGFUlu
igwCgwGNeIXP+k4SQE0rVThbJEnblEGXVM6w+9IRTo58iEjBjXTgrjlRNUwgJMBC8PfI8m6ugjYJ
HTJuaeNTKRVxmnQ4l4GtFAzboEHNjtsthE8WdEBW6+U1s2S4fJgGtBW4xIQMSNc2hBFMKSQk/GMW
yYeLVNKVgklAdJRGvBvnJI3DYLIbL5cm4VUEeJDKDly8ATOuFf33hfZzd7dr+t2zsHXr4FVBR6SR
95MgzIgzNsirGWmDGUgTKgUyuhXHFQ6zVQcJ3rLIPNfVrOKK+a5NQz++VHEUP4NWfSZbqPW1XD4m
Q08ciuM8nY1+QmPlbxmKWZ1rURIPYc4PtAKPRoMeOY5QheViAJQ1rd/BtbCbFgZfbkvVr5mDzGv+
MS4VvdYxPztpFVOoYvf7sLJtsNnf9yyb0GE3/4MDJ/qXTEk1EOyuIeSTkpPEJw5cOgIoPyUEI1r+
RNStfqLeAhnyxkikljmRzZ6Svgfi6r0E4RgO2DZjeahoVyUwleH6+zEDfM+PViXwMXGhePsLbmv+
KnQ6XBzBa0BOv4A3EqcT1uxyKWSkofDmHGmh2h6mXdACZWkejKugiQqM/kfYG0wLCZAsv5pmd2l5
64z/ZfVaM4QfT7+g76ORhGIci/0sivHeSziV3P5P/WwrmkqMY7U5KwPvC2qFUKzgCtqSJMlhMy8K
x0FrzAqffvYDTkxin6zBn+3U87kmEbxCh3jPjNInEZCIR/hu08mttVh3U4hkHUBHqChKwOojaffv
dnrTi6QGyIVKJsDI0wb4wkXUl3xG7eIM77spXAQJkAwW9itQN1rpVJbdI1kVrZtUu68AfxYBDpxd
q8DOSztOTLNyYHlVuk+eX4HFnVqxAduhX5mDIwN8ooPA5WkbOcFRvWftjq8q1lKOEeROkXKzCvtH
LhdGtxA6L3VNz5IQc0OJbXmxyTRFUYS9zve21A9z/x9qRM+iX1iY60mDCMttfDKVR8czyymK54RF
SRH5shp2gJrI8+YCDOGBYRCM1TmE9PzyfkmpQIul54exjkk+1bn/uiB7714YASfhAdGIKhwCSCnz
C2SWEGJksxr2R9pTPxGOaGUHIuBPE3zmT0AE6PcMxze2KOA0iwn5wSasPenUczN02Cek17BDOnhm
kJ17mzKlKVopkkzjyOi8KwMFbv3QEBgSsdnuL8BmlAZoLFG4fiYGcKGMoAac5uTOMjZP2/wpQo8n
rY9uhI0egY+EbNmG8khlBMmdLTmD8sOpkaIwBsOi3uc4+Z158aLQWmoNpwB6aIbH229aALlXup4s
/5zMgN0AJJIAuwolZGW0gQLWYLcByOC8vM6biyqRw4bVXb17sYN3ho7mwMOIrd3MhhYHXtqRdLnq
3eYyMQudmiG5qIO0MsEO4Uz2y1XPgEV1WaBifDqErj1gdnTzQvq69yqvkJbHihXQ0n8FnaxKN568
1El4mGg9bwWh6Sw7+zw0IuxUjpHZu1qGW5xcQjmlaJcMZqCVbA3kpvIhNQ/+5MWiAW11kMMgmKae
4KYMt+SNq0U3G1YnMyk4uoS8DJMPirjVsU8t3A4eirShfovq0kiEEjDKXWhyK7zzIl46hegH+LPG
jOIp9hgOX2VrGvQ4lJukctFAesSNM0eGLtdbBK+gxPCrtRWSp2tIKWPyFNumn+ddGmx+X0VbOyWJ
CCtYe+6kEmtSeInO6ts2Ctk/g7hpLVt5lFev+d7AjFFcHhRot67wR9aLaJeaoWM04FuoeqmKWFhj
3olWjPdOZROV96NEsE8MQBmUwX9cX5WJQQG64nHyYmMVFXWOpx/89iBHyBTJyUB1OAWl0j1D/ou0
ICl5CH9dfwkfxcDbfYApMbSAY7j5ywl5iMI9gQTdL4Ce9lhlCET2e7X/xwuhfnO+dWqvkh5Xuv2G
YgFYxX7BKeQYC97l5KRso/dvtVAl120625CEJfRusbtkHdVfZIx4mzj4qK+2nqQpHViY/SNulZ3a
CNficq5y6HLWseBOTNMOeFNAnRSsQvmCEWptXItDy8m/AJ97PDlfg9cSrfQkmoq2FO2I1Y/JPbPb
jrBcAIHwC5/3PH9IxYTPVGQ7F/kvf7yxhR7k6wHSJ0JZR7uF5zY6oGKQpGqFTDfwE7DmMBahef32
rlA3iOJTTpOxqzsoIRvFynhxo72DftFlQ6Te5NlAK42wZ/CSf+PMDMJU2Tvw0k0Iuu8Q6zJW76oO
C1cDssvR6DyoVZf4jHPUhf9Y2r3Jvj4HHjuLPXZnftM8Ahm+o9odWY1BA7sf8j141TmtItPhQ3kY
6dPaCxnCTG8k0u54ssjhXROcKB3rqnxLsGKLbSgb3T+cq+gT1ToJe3F2ML7M/46x65kKgkA7jES6
7Dr9KKlerwIQydhQnJK0NiRuoV7E7fZWmJXR+MANkF6+8m1tL2DlRldsLlbMgLaeWUV/4lmpoxeq
dRegviChgSxbcNPlyZhuk7cpqHEOXPPokbcsTJtV4Q1WSeM7fYS2821t6UaUFPfqOZtt5+BdLHoJ
96WLgsnQ5xhh30bsh49Dyx4WZgidnpUnbjrcL8TuczVqyc3HA/hORNZJaQvhFgSHXCXos6MVXtQ1
2toaoJ3n9LbGzBCYIXAww56tFjxXbFnHzhqA0deg1qpbijl7hbuRZ5flBiQoD4h+BUFXl68dxNoP
SnYLYVjk262lxJHPsIuE2pm2Pi/NQdFjCqA9fIGkFpGxXUfxKEZRMqJuicvt4D4CFzTnUk8PzE98
7GDQCIhWaXs170xV9wOiDVUnkJdFxGnSEytsRHYbYbCEE4fs5rbeiuQYnPxnG+zmi6QUrbfoaIe6
eUYC1Kz+Fg1uYibH9rlU1HdvOYHBl3LhyQhXtinCjBecmzSH5AyXywExZxrPZpeZpQbe5zFI/7N7
HlVf1/8kVF9bzjYNNiMI3ehGJWKurfu3Ug5tL1s4YGi3LTx89T62l64EefyEDtdJea9H0FI6Xdpj
KOX9U9hAvxRwyZ9ii+Jy1cD7yz4Cu0FMKUI7zvocq/OhgDb3U50trvt1LhbFs32VTF3I+sm5FpE0
4w+HPWh+zf7tv77z6lQpt9TPMe6WrVJjyzT/WicuMv8wPfiC8tuMwL0Acay2E+umvht1zY8T8DW8
N6K8kbN2xZNCAYtrBEHEoTd1UWWIKNAwKQAhTbN+5tBjYfHtGeEIGGhze5eyn6094BH9f971BVN1
uRQGOm5ngMnpcsQVsI4qV8AOx6+XPxB+AUuzm1Q2uAgv/GnwK2RiCS28wxLse3Y5xh4N4Tl1BebU
iXnqAUVvZsNq3uWMuU3TZ/kubfDaz5G6hcZxUw+YhJN48rCWpQJzLPV1u3Neekd/gaQksrSB1O7k
R01QPblbscbyOwDNfiQQlzZ5VxM5wnvsnxj7aVwEqER/ZBhBy3pmQNz4zt6Gn+uOlwRPc4XbPHG6
7h3G8ItZlO54pJ33rgDXLzVQovdklqyjj4dhQwT9BzWMvxUIj4GDykFHLQHa4rQGQztDnh85SEyN
flGlHNzhym+z9ABvevpwUTXgaRt7LYk8qrEGl3qvCppaUxYG207wJK+oG2Ro/2wC2ZDApw0NauF8
X6TeoKxnossNMjoUpgkOlE+i05pbsthllhugvXLZnbPIJfl2na7jpdPeIr0/cLawkBmomPuk4YyH
KQTr9dgQzjfdfVotD8EKARhXyEaT+TQGTaUMmWZLmPJXS1/4/79mX5iw4fbtXe7Dz0oABiAH4NxR
Kk/xqXQgj2qf74GNb3uEQzv1VKhNEL/ylkBqV/ahbtRSh+Naw3QvaxA/GApIs8/xYpw9yrc2veL1
7z5MpmCZtpphF3/xDl5Re3f8zVMxdx+FmKZpmZVhF2gx8Wm0NP036s0Iqy6265ag2P/TYunaKwZR
bv2/QrMJyEhLihFP9W5a3bHNUOvzF1CtcE8mGeKOEE7tJFB00OQWp2oB72uHkXV66R9Cf90zGTfb
CInXRxBIr+ppND6XVFBfP/hI+d3++3lJOxC+tO5XN+/RKUZ5TCPoTUKlHjd/f0VQ4bB2NS37Vni8
Phc/ZXQydAtEpNjj7fulfUxmOp8cS+KPRClxazt3gW4jms8HDPa9je8TiGrbhP4r+ti73QuEKzDR
ZyKH++jWU0M4Fe/4jJHHdhXk0QSr6qaZdSqJ0AQTHGKsbmFJCr7DCe6fFB490AWsD6DrBJafbYpv
hA8zx43hl150XtxTA1eemBMg72J0jVlUskZ5DbejiZNt99UtYtYkapBPzaSwIpjneiRh1tyQ28mw
L5O/UQGB/LGcCxLKCkbLboGDOsuBdOqZiL7TZAq8491KmTbVZ23lxy11dFj/M4y2vJhemx3OpX10
ulcd3OmzLeXAnBd3cfRLnsuW7l/yh53+idwZ11NXX4AXSJEsQIjQZSQKjrd6mXg+eX+E1NAkyXpa
nuJu2QTbplpru9513YgQWMlHX1h0TJdKKY8SG0XGSrTHqQqigSBKIzgmbilLujtCfKZ5zsA9YdQG
OEhRZQLVqIY6wCDJdD2lQFhldMo4mSHSn2dgn6VCO7uV2jYeROt7BvCtKB51tQ/adr7jTv3HC8j1
4BnQumarZOCKmXZXKlqvr0hhZI4LZ14R4sDShbZC8V67w8h9P4hXrwIPu+F4VihnhH3BKu2xfq7y
mfzkXpq8UB3UMQqiRmNU/AHSXIK4INnQTAr5pwXffIfL6/TiN91C9tudQHldMpUlmgZnqWY5n0u0
wZs6tNXudkwy+xK8Wo8rNIrnO9rbe8D71Bub82ABVopdxd9o5UdF/LydA2prkSjuHVhBGU6f8QJJ
o8utOLANKQiCpeBwSh+3Yq8/rNt2t/n/LQS0C7WCneHRJERqvIOB/D8AsPFJM/iHv7AAUe9Sejth
0gG9kyqJZGYaIzoV+hrcfZFR9Iu9xtrEAxMsnN+8CciFTjsjppho6FgTt5/e+hnrhuI/1f6GNjp2
Kpz3tA9F+FJG8/pUhrF+tPiPPx0KXYuxWJXJEXcGyJoTo19k96qvcjaRW4aPDpejAagoZ+NdSTeT
JEcpS7TKKqs/YET2OsHDZimBxvBExvR/oUQ9qc7SdlrrU3bnOvsrtV+110BKAqRosbTh3vOgPHOT
z7n2UIHJniVzG5k8jD2100LLFwn6F7ZDcu2Ghs3l33xOpkioQdSTnhAyDxXhNlofqVkPbpYHQpsf
LEEIwI5/vzsP0p3NA+Z2/lE6p5Ps2D5sGsJVQMncHqFhX/93Ra+rqPNhXKDJZCAe74qCYcbdOAeX
uwcFtFrLTp8+69bnOdfpcINKcRMxK16kcGvN9hSjx929VYhSKC+5luU/yqJLFfHEn9SR88YjPwZo
PtBn742/KAAI1HIbQGc74toJH9DM9OBqlccOR76EwnfJpk7QcgCANItKY32kQFP0t/ztzcxXoDNE
i6UDv1lDDGvAzMefAMG1l4z3U0F0MOIG28VW6hMFq6ifuF0QurnsxNUIgDS8w0dtD8H7ItQ+kg0H
vtWBQrIFGkKfy3mfCbE35pxyjAfK/KrGY2+yLvGNr0Dwme5sJGQ3xZ5O5ugj8jYVy+lX17RIDvE8
+95mcoWjYD2BAy94xwYDrL3LcbcJi+dUDJ10ir1d5vgef8iBgrAkUb0JpW7/vZeDYJDpz8uKkd1Y
gkNIhAqM/zPQJVknccdwwyfAcDiTsDx2yBwcK81pP9Cc6UCr4IsGtRPSup2snK7hYPthopf1yONx
ElPF3ZcJoKi4svs9wu+i4LssxY7ek06GbVFXoJfQpiSRBOGerb63O3Boiy7gkvipbrtlWvgYBgdF
RC2GF2l6zrlPILNe8SuXjKYucq4Ej2wvWzXkoQB4yTs/dHeboTSC8gMjJpvTkr2WhHoMAxgeYq/U
q3oZy9F1duFYxB/dysbN5I21kkX5RVphBVXfzbMXJ+T4QUE3xsd+Q1Sr/WQa71jqG39dKdbs2aXe
h88E6qGp2QXpnO8W8zesk1CXf98erHGQ44HOmpVzTnFvHXEBjshqJAy78sYy7od0i9gQdaPY/enM
o5UzOdQlSUiono1DDlmznkAG590zcuWYpiFaRe03MgXI0yZ5gJhyulklzMtBZcGTSCo5Sfr91gUI
oI/KuJ3EyJRnIVvAkHFGoGlo4VS2MmcPHrJmlKjfRXlN9/QaNH+WUEjNMOG5fyIRr7wVoIgvYWX/
PC9FBAQ7g+HmUYinT6IgzQG4av78RFOBbLRDB5LI6tF+f53FrSWlbBxvdGvGtE+zGJd3mPhDQBsC
hOhH9hj+JdpVjHnlUjpQY9G1IW6+UHBhL18Wozpblg1ACux44uvnYgW7+XnkfSG/8JNgRD+0clUD
cdBJN+T8DNZaBmz4hfJHUhGnNrEXGMItm5lw55t84bNxQHsra6wpXMCwASxvVYhPCmYSfWrbQFrU
PJW/4qSffkrPjgsd+uZ588S81RjBvgLnEnrXZ8tCGHVbEIDK03xMmc9P1x3vsM1NFUyZLJ38NrR3
DRIagMqVehMi+2pvl5useIXMsxucIEAITu2VBsdDKcTP5r3CmUbc9ndz2JA78UxnTePysbGi+/Iq
ektkoEUhRBvUJXNk3u3LuxWeuCWg/LqUJZ5b36PAXxs2fcTIrwIduU2VP0Ec8jTqjNOCQzFcqRc5
fXIIp+RmctNZnnqU6YEjWi2H1UNh3b6mH01AkSmkZUaP37BcLeo6TCli/G1ZuDxQ9ID9I9VTjnYf
HPR4/crQkYLYKpiAVr8kjhULGZfhozQMCEkYrIRrLI54HjOiRqsYc9kFh/izaI2GQoSrx5a+EJIi
ftjpQBbfkGn4ybl32k342kP1i7krxbwe1jVL1eu6Rk5jiS2Cr1Wj1q8uXO1B74yi01ofOW2jSWFX
izK2iDnQU3I1HJXQzkqOhI/N5SSIk3xbMoiayW6tiKbgaTy1u0IjGwRfm7u16Hw/eCyvXw3cgpbq
85++JoZc+uqP0fCr6uqNd8qmPzIZm/h+XAOLU7V6LQjsJZqTJcXrdtLm+/d2fwSuimiCElBVeCDj
LkQHVp1SoZ3AUusZO2JVRwi9W/W37m7hLVde63NqaasdBUjuW2S+6bmk2ZynuRmOQt6jdvBFLVPC
IM/zKGKGL7duvSqvIA6vPkRckHzCYPnATHDyocdO3KvJ1RlOHHaznKITH/IakJW7yiJ2JiSEx7L1
s6X9n46M0GjgyMFOBusJwB2HKb7njLvZy8ztvn5vfIDvVftw1tP2ypcl4KVscHca4zUqAQZG5EXd
IJvaJ1/tPinlvEEit9O2HggY1g9M2UMPmyleDS3PJwsB2HJ8Tt/nu27dD01XsNY1T+IitTbhRden
Aqg+1MFzIRc3XdehTgEBnhhsrEF9uGhYtgKkoEhvM2L+vA9+zcHpHc4I1FcyXq6RapAR1ByTNyZq
IoutgPssrzMqyzn63kaIXp9Ii6K+VDtYygiD/htiaUerwFYO4qoRA5ntlBz+NEIv26PWsg8WZTGN
OBy8dlZIRPaHze7pc+z6ZULpxbj2PKHkYsbvso7SH2SwpGjDXneXju2azXzFrkAaWOJckmrDdiHh
9DZORAfaZWWs8eiSjmLy607lh8QybIjgnjOgs4vtHuRq1I4KMsjqFIYV7fDd2bSG4YA7CohbK1K2
63K7b7ERmZuRuNdbO8/2xypxYxlZejJxUz9T5mWkYofxSEX4EnDxU7+nJR6/NtsjVi767oBZcSiJ
LHgTemkCmXsmtt478ul2rHW4YlYr//UTx8V7g3XZHdTaZAAY6CieEOMuJXnOPJeZQctd5R8/Xjk+
nlc3D4/mdiUR6jnozARJEzjNYszeQ2yXcSXjGT030uRa5JIArjA2dOSF3ErnB5Td8OjzaMEIZrbF
qxSSTuDfKsH+4erVNOcyM99RIxpl4aiPI8Ag24AGnAgAhM1qLzcDwzNrUlaxJ89wkHy10bIBQHFm
cUUWjssrWJss7l7x9WjGWj0RjZ6jafdDHBUH5dtoACkhmgIV7g2flpBugprE6DkcQQnxJB1Uirup
X7DDKnibcWS22BzgRmGBuMLqztD71qduXE0sJy+W/BlIh1KAiAnudVAQ1xAoNTF5ZY1K5dbA53EI
dUWGJ5mi6RcBrFxRimiRyN4fQJj/qUSGZqpNZgQ72ZGtcL6ABouDu1IppKgb4jSzk4Nku8wA3gBX
Da2ADL/5lF7V1wL+mdRvjQps5evrMcDwVdO04tN1lswlM0n09NXXpg62CV7zvUJwBxN1yM1XVSS3
RE9t1cvbhtbg60y3MEUaU+hZj/LzoQLDTuOa8vNan6JkBDzuRgI77zJvfxqMWKwj7xFlA77OxWt9
pCeg/ISj2jzkOrKaup8Qehl04ZdpuXXTta7aVO8Szk1rixrtyKoB9hFQ4TcjHaO7JF1jGa0vwVWl
I6jjWL8wvj9hBpvQOp8bUwaB35j+2f6xR3m7796oEKNVggCLkjZM4Px1B06zaGx//X2bGd7sv5Hx
blMCHrIoBde4js3XBOMaPlnw4nc3P5t7iaVE34m3ra2TVp7I3F+RVOKI5SN8JYZhOzoxzE8NG/43
+KzF2zxkox96kICEtTw3BLHeY4KTDWKsfptcUcmHbsWjilDeEMnjsfV3btX7GiCx0DjhIGhFGrQc
NaCa38GsYwOT2JNY4Q+3hwgZDJrsEgwc4jT+WTgHVUroC2fHmHX4Sxb5sznwcwGF7ersjSQ87SX9
PpSTka26e09ruhNVWyTlhHTGNlwC0yJ9Ot+63xui9z2II3a7nFUkfHqQUj+RJLlBP745ZvK8/r0H
6A77DzWbOAUcqIifIQOwidQZUJ2SWmxnfPKADejNap15Z9oWbK+q99JPPPBxvCQhxPcn/RrxMDAr
ANdMk4x1sbEKmnHc6zOCy686oxccQtrwdXeb9Qk1tqeySGLW7Td+j1wbUyWLmSyrOV3+IWHcaLif
RcxVJ5Ao5m5Q22YnG6wc/TexQndYoSiBaGATMVLXIfJz9DOoELy2CFpJOm74cGhUrN50LMuFFGrF
Oj5WrKTwlaBQ4odOFV9T30aN7MLTkZL7b1GZObx5Cw+TEpjD0mT6QJ/o9f+JE25ct1YukJHHBEbG
PFUSCmirFUTRfKDgIY2+i73nuHFyl+/Vkd6npMFZIuUO7SLaTsZpJskf1w3hAJa1BARgpm7nARZM
QPjf37NkcSDmVwH+oPRq3VDgMu7xyeceszqwcr2z5YvFiHSTgFwjsGkWWvaNALBrw1OyldJLwWLV
ijkBIDXtS9j3HXnxz+THntFL51XFPzrRG5ygI8oJwxxAYjYnSGQsn+2waYCn8902AsxjPQFrCxww
08N0oOUs6HzgcFYGAg2QtqMID935zMMSGX1HaQGx8kHHFZ+QbdLHWIDdLbWUKJyAcwrD9QPoV9JR
8nGWH6ZykocIEN6hRdNeYui8k7JpuNMnu+1h3nl3d22TrHN7SHhcxIQ3qt2+qKb+zvh3/zA2tvVU
rOhOoBoGE4NmlVl6zereXuCCE9+PMmzoxES7zt05Ww/fnS89TDeTVwIQZhTfn9n33UgvtoY87N70
aSAxlJamaEnGyc9A05F8dCZRkVJv7w4W9043JDmA/EfBdpMlzSL+3qMxfSNExLerWjxrmDTdKcaj
reiD52PeU6zVLKb/ARuetoVzJcA6smxz4BMeXgZjMK4S71cqotbKRYb7kYOhUhl8yP9yPrkVrGTl
4eiCz3UQMFmdmF/ubqlpBzBFqujKY5AQQPKvhH8wmxMEhj5lAR6Nnfnrl4MpKz17sAOhF8DerfQf
dqn89L1lNyDEhgqUllwzoBlP8Tr5b9dmIJjADb1RybAckUVzT4uc4tAfbgTR/t0vhvlJKiMSciMc
0aFPJ9H1hMYBjrvsIhtrJryT7GbrOOAMGyTfIuMIwe1+nPaejMSGQKAeO0ToBYWJ5PIHX2waIQFo
Z9aak90wXEkbe3jnTX61kgDax+AclUUl5xpLAdd+3VaXXHDFzuaGOQwRivvsbuUG0k0eveq71Rxr
qVevRry84fVnD8W64G+jytYfGg4cOJwgniSRaAK1ERxyw/cWC8UEFSOSiqRz7uwJy1SwwvvseT3p
n9X5qF4dBsRdw5h52TX5IK527nWIGalV4uXbrYIy4+luj7FdeTUWv0VkGl/B4wgSmUNZFqBMWoiG
Zi0mMQjB6aBuOIIq3sXBA7e8cgwgHjhlSzOVAnmKFKqLiXb6LyerYjEou9TUBty23lB7s0uR0uAv
s10tK8x8cPg+MWTe5tPHYcea3+qD2R26AY4Tk/9BZN32hjz8kmA2WpUGS4gxcRhTvyt3YR0F7jso
KBoZvpW0dCg9N/mz0oyaZW97lcKZ61s8P7mRLxvxyeUhCMszk6u71Ii/L20XenzrSdKvKMAuFtEA
DX+ioyjSTvcGOLyYAJunuP9pb7kLhQLRlLNCoH70F0ps+Q3+xFoxlJyEQ0kMrxm+5Y4+gVHOvwcf
30mfBgOMGXSTzaMGYKywerC2afbbm6OmxsuznJKwRtP9ms728DC2NgecyR1X1yLGQSA/pNhoqd67
g34SlyaLRLCI+4WFBjIobvI0l8BnEygfj/T15XfGyxGj2H5qIgt9GLnl0EEJR32J/uiw0Yi+8Kq4
LsliI4azIQh9mSL4ZJYoW+dQSAkJs8kqzdq/KqSJfXpJcSzZLfINYQvR/+RRqBxyGOvkxhx7JeUD
XQ3dwbs4pDU/OJAFOdE1SjsJL8t4GtFAaoPPoUf45mGfcjLjijbHBUt2daKNntdtZ/obdomvhU1l
+qfbKyoUfSD5ZDFHR7Ag16N6cfM2Qbel4ji3Kye4ARR92Z8Ouosm11Yf0Iqy/GNbMyrRxS2kzCK2
KobM3QC5xevhNa9r19eklU/YsiD3MuKQ4mUVp6Nx4age9iakwUwxFkIqw3SuinLYo495FxyIWBqW
myafk6ZXufplRMwS7DzpbXutTUJXCARuSQCN1afvlvoYdM4zXfcQQ9GWYRk3RDm3bq1Mm3lOZCMR
JJWkP6Ir6Eo7MbhP92xSuN/7S9P1CSjtM6WsIDQoK65EdNH4ZCuhZAWVkTZLNa9OREPF64KrT1KJ
KRDIZ6JmZQx/L8Q1Sx/1oETEdlxfI67xCYp/3ZGtcb6mvrOL1BI0doqP1w/HZimL/u46Zh//2TEh
pUuBqePToPZZhjHqn27NFsg66b98Cz9+ldh1biKvego1b6kcuQsbOB1pOA8P87PHTR4wRGBVAqs9
3Qyq6kYYd/WHZUbsTT7hIYYERv0heEsVdSutOZyEe8M7rkltur/7x74m/sMk+hySQsoWIGjTLkrJ
wa8aUfjS+8WsMdPbWHQE95aQ9Bfx+4jShR9qrJja1sijQGh3MRFnfCfM3aQUI99mbTmuYAHdwd0O
Bv4k1WvEHERivjt9Xgnc8ZVxGoOjDbUnaFC9VOBc+EIgGILRyzV53c3nz448MbfAYGqlocxCjVZ8
j29Ep86OXrFMGPaids8yaPUYqQLTivPcopChQMYtlJwn1PFftdgh6GSGmx2mMzcL1jkWg6az4kt9
vBG04uFpKHs/tQkQRAl4GMcoPYOKfL1d/lbjGssIOZQEPkF49ORwV4+KChrxEucvgm9n30ro7PrV
ehXZMTdhcSovDsH+HgWNibv8wbZqLWIcBX4cpYGAtQKGyphBqvgkUfwdFRbvxPVfGRrn9I0wRaKj
bTCnGv2KtrSxr9HjS4mMPQYSJMs7XM0JmfbuS5zs9auDZfU+3PVNySzvnW9OIIHVXSRcFH7GXnj6
KMVv2niq2ggmYD/gvgk4jyrAG3XZ3IbNmX34aJEsT1WMg8sFbsDay5RekHZoVF1/Unq6bCkFJXbz
nV6y1k/yKb/lJtVz4LhTkvW0qKnp6171uHjMRnG8QCOMEC965x359X/7wBehreojAB4mq5KFxujk
4SWkAxWBv8aMdHIdY6Xg9qwXNnkbSpsAqddSmdGSDxBZacNKRIE9z4C534qAoWg0hvDgaQ7CIKt+
et7LGo8hO4i9vMTCXKum4sx0XDWeak0tuBYoH+2108t9ucPXojhQP3aB9LfpFjqmC9he571SStIp
Fo8ZOgmxmRbfnqAPl9vItX7LBmtoftvsUzUpTgscEQQUpY6LV6HssjGmsJmTDVmPvnC6lCCYgP+1
6yr7WxBW7N4Sovx9OEzSAS3KRowqv8irewEclD3fUwFixOebNwAhiwqeLZ6+mxQ01Xh9+IilfgrJ
UB6GXEQkiDL6rIho2WjMdScyG0wywPRX6cOcGASus2A7R1m2Fmq9niiJgXIc07vMe+jeDYgUpeW4
RP6q/UISm25LbYUpQmy8Jfx6r+iYd/ffLIwSQ0IoIg0vZQs7uddI1vfkafplqJTOoybm51v3wNHO
6j35SpGlhmYaqvguvlOvMxf1DXFex4FVe+tZxahvHffSCfjN8kFDlwSy9JFZSnUYtap85rfFE6gA
BNCnl5Xi0IYHsv6MgLzdmsPX/Q+eiLbvQMDDzHqPJGIMkQTWvyaik05IW/YAnriFITXXOdfMViQU
eEgZH31zM54dOPdcN/LbjCMMd2DzRKwX6txO0Pzjld0/oayrRH6R3qeOZ45I/NigmfJuJjtQUYwL
IAfaVkdO/83E0S9Hi5mt1rdY1Pka1UTNCuGG9gl5c4TFKUxfTtVzlpDa5uEzAX+zDyPNnOTeW3CV
tzjJ4dt0vNhDp3cbPpIUA2i0TBLsRGz2S31GGECw1rAGQ8J0AF4CquVZSWSST8zoHZqsRylDUOrm
rc+Oi1fqa5HziyRfRwDiR8W/sZthCs4oCbcbCUWFgzpf9izcgB0NxDtnIzmaPEE299I63xGeSX/5
onSE70zZw67tv2ctwWYCAOfi7mUvF93womw+0VDUpS5ATjItiKrQD8TFVf+jgxDPFg7enbhK4Lp1
eoJkLgiBBryAyvrDAhTwqPDQv1PPcU1sVrnWO4iSR343xVPSJ8x8ij9UgOn2dDX2O/NH945ZkGDj
PhpSd84c390VGiNNtcMM5wHVJDoKXWGInVFX0l/7RC2F5qkWPGMM46iMLEOJ6yi53VNcStstGBz5
8arfItX3h/ms/NBhdw1O6E5HaLR91+d0ijIPoc7wEwbmyU91OYt4bvMMZKoXCHSi59VKCV8vL01G
0T79s7rE2X0uHB4vlOj7hkl75fP30Lv3M5hr3WBV41jq5U1bCYM/+LzNzIojIJtr7WXnblCCysIH
4u19AYqgnYuQpZWF4nmpUmSu8HoIOxfhwqGJdW0uuBSA6jxJUFrXe/YKXvOyDj52+NWjttlp2MPt
zNF5xRYO7Rs6PvF3VpKHupYB2EXBSjFpJswKRXypSDT84lbHDlz1CQuAQtUHt2+LKtp/Wn+sonW3
xpT+O6GcCao2ybXn6/x6n55mCOFoiR3YKFaUdeKhC6LqlvdGivn4PEKpeSCDx+W5pbOejbyLDuWi
HOg8A6KIplj6o9PiswxXJ8mwhNGjOQzO+4AXwr0mhgiWHZ/oN85WVpDE1g5ADSV7+7+gwr1qrHFk
RI+w3XEDZt7BYZ8eblO+fBFBqV1VDIgym5NhrP7p53Nkrmh/UsGxPSHB9YT3vuS7aGOVqbaWXP64
ATKCogTfx//qhLC3IdnSiQfh1a+jMxKPhaWZHgENu5CVv15VIct0RYdmknq+XB7GRTowGDAvMReP
5YMF1Nkd4eAaaSn9o8zBc1sqj7jL14T4bIfqFsDERc066slMDQkcDki6P4x5zgvHjREICufpXwS7
A5XlIiRuN/NepVuokOlEI2WYPI++eq70pY7MP5CW/jnS6zZbIMb3v+Q/KG1fV1oovhwlAqIUpJk9
f4myfq1qmZ/LpZmUSxevf0P46VorfUUDazt/A1Cuj45UhdRo64Wd/tRg5di2YVPcdXKTeZ8DDwum
pVoUfS4QAnNfe56F7XTPD29P4GVu9bzszWnrncaFY3GtQ+Ju0+6aK5M/AD6nqkPEuWqRn1r5804S
AMtXR6ChFfaOh6zpF1GPgLRjjBG2nqC7UaMjEdj5s8vnz+ijtVbIBg3gScetLUR+ScI7w2QnZ4KR
mrXndxqgSOdrKRHpfMed6uDVbYeNimF9R7zKszL10cinUvwxTiHtbeujP+fQULOXPWRwRgMkZLY3
H1VDUyggN7C1gaF+DpTMMgSkSB0bdEe6miqYHv+McuT3t2zB9rZyU3neVB9yZRTAyecJTkRYAdSy
Jg4VldLCrLblN+Oj/bNuLo5+wCJfuQLENQIQ0D1JgV8IDWZ6Wp0RPESCIPJdWFHMgHsuXP1DKZis
z1mA34cL3ySD6JLWFrnlgYrbq2pr0QFgrdj1XvHXCVheVdUveWTejWyksSFEyncgqUsSZ3h2nOHG
2rfMerYrSJHvXq6UF5iyVcEoVrA/gxEO/YrNE2FYpVThRpqbo/LH1HLd/FzOd58V/P45t9EvPp86
1ZDTcOYmUqztyXqMqgRG//0aTUu+m4zKEV2LAiPJsvHqwHR5RkMfzlGoOn6xNivqAStmrAQvR784
RuZKY2YQ+qbsHyOF9Cfv5gbmHpOdaMo6gyfEvQGgcDWgvZxCymCfIht4bqMbF3ZsXZcvUqpmgSBC
eTZF5ToZH6HavYPwt7sV4sz0E/hsgJpJDRXzxKXbR9Qu/QNMe6NNQSxACGS+UuAnIxEqfQ1yeakJ
6wvS+DP3gSFtOAzPbjlEaQ0CgyQm05Fu0C38VG7OiN5xwVb6K5KdbY4Y6kRWjKSx72iUBOsZjHGX
NFZMiadg4XmqOOfIdgC2wxNRIYcEbX9YkuRdcEl6uctuvnATK2yf/C8qS6aMWrk/mU9wW5pyt86p
Rm1RxzDf37F8i3GRCFuQB7YdHfJicByELS4W+DFvMVhZrOQOapC7n3lwOCXBfudkW9I7w/07vOhX
b7DRK9vBSu2DrEL6dh87ZpVW2w8r8SH9L6cQnz7/V64saOrETmmLzl1S1VopTQLRLD4m/hJE5pWD
4IKOryrIJCP3UNiPUDCagK4SyPGzAGjH7XIaewrQA0pxM857tQGNMPZS1Pes/NFcXijKgK6W8DN8
lWY8DfXf3lFsYX+RFfofFUCQmsjT8l9Lv6QoMhdau8iAZuOUBltzXroMmqegFP/RfUYudHle3FdC
nycygKcJal+L8InyFmirARm12S0J07XiIKYLMH6QEQ1FTmSavW6uMFRjfMmC236xLFmUBL3SiXQV
HwJ1Poxv0d5tJpSkGhWow0qQY3A63fJjzoW2p4LEIVemxdjCDxk/JMt4xroUrtCqHC3+evS/xBCi
8bIg7gEIcBnfoDVAir721KrbGH6bR5WzXoa7a8JIKouEVCLxpGpuJnQ9N7sFgZIFnNgT6qywp31m
TEL9OJaBMiBST+RJALUcH/pFruTLd7lm67hEw3qt+2TER/P4OavvmXosE1SpY3K67QUpAm6W1O7N
HNlVtoJ2LMZu/EtXPgEqaCK2Qhmg/Iua89ngekqj+i+M4NtNIb9muDJb7UnNKwZFsRw1rm+A0g1G
LI+10GE+c73v4T/pb/rqdycnR5EU1zodvM2btk13ozuWVpHl/BCxk863K3NduqTsxX3EHq3tkr8I
lkKuOsQ7ooXB8QRi35rPdESaA82F7t71wMlfjEJD3bhT9BUW/0365TAbM2+8rdBA8t4eYIb1Pr7d
WEUWjL5c0BKCqLDm6jSTatn0K/2IvIEtrwu0+C4YBfHt+I3IDPz18jC0vsg1zadUCI/DZv1xwFGp
gtC2zBOxMyr2vPF98nF32MceRxeKvSFwr8amOzSl4xOK33dfcJImZ8BcAUrfDcU7FmupcjWYm95e
5zZTg4nbzKL7iCNTbVJs6sqqUs532qBxVJXBaZ58B+loDg740ovMbSuECu1c6d65gdbr28oSEcvZ
CPN1TVq59DefTnTqxK2EUfbz4NdyuoYDRpyPNgWpnwMa5HSEbHTfFCcH8gQybrqT76dtBTE2HiBU
WRZENDmnGv60JqZt+4ZIV3aThsy6/tRzH90nFWl6Gr7sAMijdr0ex1yWZK9qNDLA5o3UNS5E5Qo+
f0qefl4JIP43rZuPvZeE9oMdaDsYmPwMBxx7xNUvBClVfbVMfqFBQ0AfnAdVn3IuyQgk9OnQTAWO
VN+vIgCS7zppzNA0NVoiuSvuKvDSoTQR6/9Z45GcDSyFmH2cEczadt9lKqF+yM7jSS+apBN+7Ial
t5Y9rdhpXX5eGwTIA4Hnqaj6KFIx4oXaXLx+j/IM2ADnVwRdKlYfNMC9NtQ4yEReJ3rJ92rrDrII
NWHGnw/fapfOl/nO/lOlMH3z7QFfbQvGpRn9zB8xNblmIvmHHjRmuHyi5IyPK0aKx4QhWorgFZpn
2KC43e5fPK3a4zlVAQfzeK15XP+ExJYFqifI+pZeVaFUJS7NArs3YVQwivDe7933JlbVjLeattYW
Mr1rkB2YH33foF4bMx96pHnI6JFoui/YMENNRI//KC9PrAxhuizn+sCWl1oKPoLNbdebPdCBP0qe
Z8HABnJ5f7EdnThmsweFOSvJXxELIUyRZzETFGXIre2+P/xrcbdTYX3E9aXj1PoiCDv+yUBsNEp5
VTbQzE0gg1Z1id2nmj4iCZub+H8GgjQrZdG4jw3GSOvOmpL7wjJPYPwI3cnsSKx6qNLrN0Wdazbt
RIiF3aecfsJdWb+WyKOA8h8dHjy1JnraAzL/8PgzOLKlb860kCY3N0vRC7gbOLCLPqd8IA77DJ28
P6GdBDd/uPq5Myn4EcrhuPXR2JnSdvydI6ebUZRk5KQWs7TUFvlJRCP4dFG2rL6Wf3VNctwxC01h
3tDQCFw2vNNfTzcosRMfebBTt/bRU9ClDcVTJEImB7wuJtEHWNmehPlAk/q0AhJf18w423RyiHzr
f5Hzpzc8ydyhHeDmG5LO6S+rPlf/y5CfsdZNiGtNt4bfpGHkNhlfxZdiMyGhdQfN4BX+Lvo7BxR3
45ukXg+Keo0AVgUnhENN245pcIB6nsQGJDhuEavci2tJ1m9WdBM+tpgDs/0sMue3IzBq8rBtQNL4
d3AdAIuWHiPvcJL2aydVkoYxmnAcHEyzlmjbSs1feRVHI6ZANsXPcAdIrxfGpMV2l8tvAYi26HEX
QviiLyGZlv5ncqO3KlKoG9cRECiqmNXCvPfO0doaYWb7NbLBvWBXRzA/Yhihr49TqvYXlv0dM5hL
n287tvSMy40jq1RmauDi69DS4+KrQyYgujoyR2mQi3caiXA+Hg2DersH7hkgLbBQNYngGQ/EPK2k
/WOb1tQ9akVNiSktnWJWSJc4vyXDC6BPYuAIRXUSU81xj2FvfEVW1ljPq3UO79OgjhlHdjeQ8LLP
JHIabBK8J45znmh71GrMWWwe2fxRz5DBQcai6cNkXwc3NwOYzNZqwYnYUvbAUAHIrRnpjt+tS13w
Dj3+DpROoqnlVxRGE7NGYVVWtSidNbptnS8Owv8pYTI5PkZ+UzER4gpGARCOnXNsX90lnB+QWzto
G0aMi+s5H/npkqUl5gsLRR//pO4xkOr9xWFgs6qJqZUUlFj27t7AzfKLo68pC4LB9vIHkwPaMmsS
oamxD80Seno2nS/SQBE67CjAVG53ufVYom8WS+Qy0qr+u/Bj54KCBMoDeSarciLFRmkZHJf2lsE1
9G0bIqk4DbqNNws7QPTXfQiETfTefkVEi1sSRFbfsUUjvXgwPRay4PmATp2IRdhziklgj3g4/B4Z
sowXkehAt9Zi0VfpkwgCHo9H/zomtn09mdcL7XQ+CGc/F+iD/22s9nrBnglGAo/FAu7aq0HPm5P9
kLspHZofrMw9YVvEdnDiUPsH9LFHLQjUI1Krj+8veFAMnW4iuqwlECSaZznHLELTU3yxYSGjBrIq
JXR2VsQaPIRGIkNygcZgdESunAMWgvl5az57N+0iSVLfuWa51hnGOR+iu+9aKfanZjYCfbJzW2hm
Y91sIaCH52SuPbIrNJiqW5cfgKlVlr7Xaa9p+zNeES9Mcjbnfyp87dS+eqsvXjYs1S6iaZudnQuu
o5+skx1n8V1fBgpi2Pblnlv/oD+0+WAEbj6Raxov68JYwVhcYBP8xtnECII28IQAc+NH8pBkxJN+
SxulfrD19oyf943ObOuCJztiT/Ku2p34c8nrnu30tajoFWr33qN9H/ZLcUPWtVtU6+VLo5X5wPIN
a+oPHv/2IMJDxjrEUaZlYh64fRjRPvkaNlSa0xQeV/HbsznNIZN6RQRnU3tSdAJoItdosKo/fRFH
xZaY+5T4qaXMG9Tx5dw+JA+NPFVyxoRiS0f/DegITaJDrEdU1XucQukUi42fs3y91U/208YDkFCS
wI5TVJYj5DALN3Gye8ocpSCPZjhxWgGmWFYpaX7d6NjsiA5LbKuzM4meZ7aTJAysOR7f+Vlsl6wI
RdTOo6TpoxL2vQRsQOsj3DSL7Ka4012DtOXWuOmY3DsJBw9Hf7htdeKo5Ol1gIEPDmvV1DPso4Bu
/GObiQpPqVLouYIVNSzthfr9yUFatBDvwHC9MIQQZo1EyBPrlHY/WxqGjKTZtyng7VNjzGSAoYW6
kABGETDUgiqzMf4dkLfOD9p88o0COXitvp5W/P+h0kaw+1L/VNLhkVMOegVZjUMhPnUbQXfd1MC4
YtZawzas83cxg9w9ahljrlshEBYrHjMi7xIg6Essgxm/I7fq+uhzsUYfiKrkG66O1P+WVjMl43u+
oZdHR9Be9q5Wf0oLvw1AY9zgdjr8U/q7M/u+bFEWZQmD/OIZNF7OIxw5aTf01QlCeB3B4Y5q3jIA
qJvWd8xpCMwnUq/u1xRynNJBnmEOd7dURLF5ZN7GkDm4q32pJWrszqPTbbchjaec6sZJHwkOa0RL
/cChZvLWrZWZEWFpLWeWMW2FHlPFuPva9po9sgjHbJjQeDP5CmZCO4Ou3mnA1eOnJZfKLcicUTe9
UGFuaZoCIj/QZ/zRMiF1nnBnj/xh95/VbZGTuTJskBwFdVAQ7JdVE8w06TTmR6D0wYYd1KPm17b1
q9MtpjYB72nRKsVlig2xPSAfA0F3/BaA7QLmcuSJxm/VK0QBmr0z1D6F+9RiHhHv7iDNkuz+OGcu
aRlEG6v3vdhlwYJH9YQuvCrpQ67PLPiDm3fixU+XLQA1LX2OPgJe8WH2qhvj5YBo7f9ehvri7/s7
FH7om8MDp66p9eNCL9fms0JCLmMfQRB64VMcpqeEIPdhi2qhLKQ/y2+tjvhJwzjRPOfC/OtYPk2l
XMq1QSmsSq8Rz3W6IM0JOpgOqX/Y5vS2YVmA4MNxb9+ZbrcZ+H5H2cFjtekGtMxXLAEAiub25O9G
MJ7E+/PPitDIyVN0Nw2aLsZdX9N1ZJ5aijc1/jnBKMLKQR3q7ulPkltmpy872mnV8BIBh92M57CF
V2yAV4Lb8qB3q1qh0fuidTwL/4EEVn6uPk4tCaT1e/6kyIZyOphiX9+I1gt73TD7Asb+W68gqQ8I
JXxtYCFgfI+CwCS6URlhHcwARoDtfSWgCV/WX5OpA1L1ziYeEifZOZqe9GT75PkVdi9R4wALilV7
5FN7FmN2anGeoo/vviOvOcrejzzYE/emw2KkhP20/zM4urFOPhDZC6bPy1wciAMLeChVN4HdxnSd
jG9oosL2NU1UI5jccP0D+N7LzOYrcPCf8EWebr+DlRf1vueKfHTMGcM1oHqCS/2aYCCBxXe4FcE8
7J6+Xjmx4e+rQbh5+Zimo0ABtV8AnVQRdYGtaNXdpcsCkLxgmA9bZN6oiiVrlRhss2htiUk/FZkJ
h9y8do16+JGliVgWmB62skp/7huA7MEzWZ9R+elSh6N3oeTtw/Pbg1t/x0BWb9GrhkmwZCSkh8Bv
0FbrqJpaxsFv5zIZuryoi9trvVPGiCo7kZ06NOvRqC0d7CH22MxfPPUA9GU+2NlnKQKoARf/o8Vh
f+1TF2SiNDXDg04VVn3Hk3aWXQlcjLtHTtkFENSOBIfobWrfn1ARY8COh9VswsispNF2URnZkatV
n4lmsi8gOfkj/P6x3mPee8uCRHhPfSdj1F+n5BwxTDoIPgXDt5lDI43pmr+/FFa6mhIW0wTtB/Qn
brWlwdGyFLf1trdHexF+oZO7aECRvG9+YPM7Nq8bfl6g1aYKOXA6RtJuYJdbhpcUxhHWISu59Rh9
sYHC70kIWCGqn0pxI319yYz82bZNApc2NG0GVXLhR4TwFGK0wSDm4/pcIgEnDY1D6aTgTxvQiO/D
fpnnZxEfp/AXouGRW6lWYDXskuwXz9epNnmKit1TvwRMfj6yMbyXZ+kP5LFf8KIAKnSN9k31j40y
Li+aZhgu8aOF7CrDIDKSnQ1tUX77PEbx5t4X4e9u1xXm1O98YYHx/g9TD+M9uALwbaiTDv21S1eg
Zwj/oadGk4OBj7K5ap8Enyo9CUbjsZibdScqTcjkYDFFrAyEYjxC56pXBRP8J2l0QCWlPcAE/VSB
Wz+2KnV+pd+upDSM2owK2gxa/s7zCAiZ3xSql/JzXIO4PEw2xDOe/xQvIFcpCFVxAMD2FjF5n2Jf
5Mp9Wl0ivpKi7BffjQeRqkw1QtiQVjYaotEELZoCXFagkC65mTIQa4vcxla6i3B3MaTm/foaAcRO
GQldiwRICp0HyL1icYikkWAZH/At070FEDOconkkT1EOoCpusE2XZZfuN0vdXBgG2EmHcQI0A+G1
pUsQ8JRMvwY7Cj7T2NUV2Cr73pgR5m136ISdERiQKXdVd+NPZdjdRdvv8g/QKnEiWPyCm9HRbm+k
+0WqZlv9gIAsEiFdIT0dPsUqaEB3k1feew29DBzi0iHiqWg31+wEmOM6liwYqwkRw7wQMzUgsEbM
hUBivyYhb/tT+an6ZMh8I5axd7QhaPSzEUE+OaremxSeAtauXl41XZgHvd05OoQlJlEXpX2qYI0R
gmrPaTOrCFbRVkg2iLU8JC90wZWqrfq5Guih25Vuj/8nnnejrDNxbNvMsJgBOXsdceZak0DMZR5f
KGctQ86IXjlav4CVEJ+LUhhR53+1xHaCFr5z1pWaB2/ejCjQM8eoW19pWRN40cYC2h3xmEzWNll7
CyinqfxtqvBNu8J1yBAWPrfhlKAFpVmrvsDmQZ1QAruVVIotpl9JdvV9Pv9pG1MVUXxWMcj4LYMc
gl13dcmG0WbSj2BnqnxQj8l7720BfGVlfQ0fip5DIWC8pvpG/w5RCWD4P2wR7DEbfiLLJzo6aX3k
DDfGwHtLgRNBWdFO+wb44VBYB5i90/ues+011aeYoWenZS8efheSV3FVMzWE2ZNhqXYGr0SjXQW1
trez4K5NJ0fzck2vUR9NmLuovp3+zBgaJ+7QLgsFv5BVbHEUJiLnrKk/5XzaaA1s+51jiCWe8Oyo
+otS8p/C+rLP373pwftcSAod91iX3pU33yIoaPzk+8XkA5/ZGVdrQcNIQRzXl6rWBd9zpjl7/Y+n
bjRUCwIyXpe06j98LJv31jBVvHhV6/uuwsRnmM/+zpzjSWV6Z2pCDk8ODo7T1HVIV8Nk1VnkAnlW
BRZFT7r430UHMfY8ww91OrlPHOYwJhQUgyXtku9n+n2YweNk3NTYed4a7O/Fc00m4e0M8cmsrWCr
Lg4Na+mpNOmrdKG4KHQE1rTN+iO2uhPyNxwZ6pCngXf2aOoiIefEaXdZPGP7+1CyHsKVpoX0a633
tYFUGfRjVcVJfiI+nbvOlGIPLuXWJQRkPGBgsarUBmKTjXL7wgS5OG4N14zD90xMdPmxdet+u4Gf
FFHJqAOCdfqNBi9X6zVqQJUwlMJwzOgQHYLgJgFt+GGvP/tAH0BL4DKOqB9B6OJUtTXkC+lFOObW
VEMvFBY5a1OmWHekj0qE/VEXuxy6HdY9RfDFykXPPXL2gF/SlQ7HsdsYCoo+JLMwKL48i1AY+j5n
XHwKrRE4YUKy/Owv4I7cX6siNSZA47O3bp9bB7GIt5qC0gsbqEp3HzKQGP26nTjOgB/+GogOWOtv
BHAfupzB0JT+zkw0P0g6Kg79lxebkEx0Qygmm/wpE03L+QB2D8S65zM3PDfkIlyk8NgutVK4BUiy
ZU2ARYKL/puFuhlvJtAe1AKVgexSWQ8gzD8Xy5+JQbeLybin5Cj6BQGo16umdoRXohV/VkTqGX9P
Ze2TBcXL9ZrwJYJDbeYrtWEkD+wMgmj/ODuHZgJLsszRg4AOwvD7nXwTFGtIqMIE940P9+PY5kv1
IzSFfHAEjBqbKn5cyQZtiMcjeQ69ZK0JyCPaJV2GcPrEbeomw5x57Za++z4cac+a/mrNqPA1S1zl
0A8l9+osJT8VxJb+m6Hdw2G/H/Ma3N7K8uvgDjXpNYeNUMMau0oHpXNjUH24DodZ/hZRkdHm+F85
5CEGBb7nWC4NdrStcwLI6FcLMYHa9jPa0QL5NvIEimNhjn5e7R3Xqb/4qZ1tcKSLTY/ZWpOozjRG
40K2ZW/8gOn2qJ3r7illLlftxn47WN8YToVCl+hgBaxYrvRkrY8VhUVy2GCQeTVyw4dQy5JQB0Xt
xmq0ALFVcmaDlqt4IIgsoK0uaMiZ2NbBsnlBgqlcG4S8/DuXPR4c67wyu1U1ICqJriIChBocxIjY
iDgAuyGWS+6Aa/6vx01yT2QhI/lth75pvK79CJh7p23i/ljNlgCAHjwoXMs12HbdRIRI7rhAnK8g
+Osmm8zLCLMgUdcaLRiD40sfWdHgjtsUbTLxRklYm3QCRFrtsgk3bpr+PHb2P72SzzgCXWGIf/xp
LfU5tjYkFf6eh2/nmRbzhQQG0X0rZEH1P+aapPsSXugz0s6kSYnYI4PcGH+9oTC2WDYeBGYy0Qub
ZgJLt2cWgU5THy3LjDxI/XzWqED4g9rdrMc5Mus2nSbFOHmMfnO3YDmfaCMRcsbX1414wRvGLE4X
xGV5SazAxjx2+CwgdW9xBqDLgQMEovcJeDK4/bKXPYN45gqT24IiWcQHS5FlZodEdZvR4G91VgLg
aGNxj6pBsOwt9OBfMgOEc6c/3LfXkuYC5oaGCQUAg4CVRVb6j2qHzN+dqGbNEhOlGd6l6IDTZNFU
A4FlFpWvja30If1xBByRX97gvhtVtJnVAJb/LaMhSz8VQxBYSRh/329TVL6gmDp/El4OD8znhpjc
LwV4T6PNSNb4VeJsvXBXa3mPdSjIV6csMjVkvp6aV9VEfFi/u8UXyP2JH4uNGLV76fVY8Y3HCI/l
Sa47zesOSF/rw/IpLKoizgrax7TRg3BqaJnFvA2XMrDHAvdo1kIyycrzrt2LK2X+lilp+ax5MIxs
n/6Dp+AuW1PZcgD3c9ijGRt6OKsmFJoetQT6mT4QeRwgCoX6mYxoUeaP6MeQjomFF6Ch8bVfnCHa
HPWGPCx6rGWRtXnO4vYGNsiprmF5H5wGKy+9vCFL90xD5ht+eNSF0k/33m12/PnngQKv13vmi1/B
eBc3dWTtMx2NDcx+t6/qlDBqH7xlalI0XN8sCZL+My71TDcSJWR9aalRBSUo0uwJDWOS8SZ9CUWx
0gwFBNz+3SCB5O7NL2sY+2z239FyHXe+ZhZKvWaQk3v2Z3Jb1E7xjEuB5sIoltA9R5cfZsc54Xkp
jwjpQf+/JpIgvLE1rwmolfO7vAPggXGRpc0cBQMQQfPmBBPpvfUGxParcALoWLObrx8sgG+V0Zw+
BdoJLAIbKSgVgVurtQ066bQlb/Lzb3Wdjp8FINXIMdMLBsQcpBlLsUU33WyU02LRGX8Iz7FcWGo4
Br33Gys6TgZzkSkBSKNPujRK1Ppbxo/ilvMGhFu+2IXYPOKjlKtiz3oCCK/ZwjoWh3Rbv73EZcOl
z5n8SWKrKtTyw+jF2BWr3TASFU4seNRbwSxmeDQJT0DCovVnkG0ghRBi710N2wMmGaJXl2fe5HNU
FYJAfcKjimlTtR25Q8/GnsdOnP9792SK4bMT514TXu0L0zGgUll6md91ecKI2Nm4Z0++kKCm5DuE
8vb2VTJHqmfwLNWX3qyyegIKiI08QYxXWL1194RIAM7FuYLw90JhCEL/u2MhESFKlvFxXQjZjN9O
P7ebU/nhuv2XBxNuovvhdP0xLRZNbRP++cxakLaRCik0UjCv8lO5ZAHAcM2yTcNWtsjMAJqw9H5B
0VP/Ucx9+6O4TmH/JVCYrhRgqSoovW++tZM5RPWnD5rLIk6z9hISWX7HoeswYQlYWTaMXB70Fhc8
1UPf+fkB2LJEmx9B3UT05HGVmn1ME7zDBZHHvQ6Oxh6euSMjS7wIgBjlmzIMmS/QSQFuIb/bFJmn
zElQEpdcU6x9n7yPnfrqGyfC/lbHu4oCPk3Wb8k4dMjWMDzboL2LAUgzL96zBTJLnefAjSAySe8s
Fc7VhStpKbIOrSBRsAwWMWqRtlZdsgTVQWCBPJqJxzRMOLG7fQwZ9XZrpddWEYpXCyiW8HpkXijl
FXgn+CHl21VmfgCj6ZijfwMjJnXevEVsb+3BbXnv+p8P/Tdtk8he+yBVfKxZK4XkSF4LqT84b4/3
Q+h7Rh2kwqkNrA810MUzyqGapS1hY1Xyc6TvE5BZrYmrw79SeBxKtvi99BzXcHs6HDQu2EId3D6i
VkWpEaH7F9nuBLboqZsfC6GwlHHlI0BKCVep0qiiB7/6f/bgzI6N4DrE1t/Dc0/1ppSVfe1ehLzX
vbNNIAEz11pb/o2j8OEiQOFmlOdCu4TFuySNGnDqVLpYlJEvpj1N/2Y/IntezmkqXzbW+L1ehRDL
rVAQqICxeIUnG26NxMf2a+8+EA7idkQhaMy53yT1BTIP7Gv6Bcmk9HaAD56+qAUwVLloDsP25cws
OSdzz7BpB9TTK1x9OWptu8P7FMxzKTWhdfV+wjhsdYAPQU70P9hn1N9hQtM6kpFHCIVtoIabtsHK
t3xgilBD2A7bl3xkr2tr5Zk/CnZyzRzQkMXr9dB7GqP/H2/nHHw2nxBuHG/XZxV8f3TdPtXT64/c
Q6fhew8Hgnja+SUy/tAGoZ5JN6dLaKJcIiWuBfLUhhxzo3dF4DpmJk1fc7FDFAzZidxi0RIVAUZp
9QCDw3xALoUGOydraF9hLmkKVGmF8iUBgssxivqBPsY0KHe8qbB26RLbZnKhf9wqk0QzBUIiTbCk
koLqrotKatjfbGaB1a2iCyHK9DpM8IIYG8Qff/Nfiqky3ErnnRlC43gatmHlywIW3rnToU0fRL9h
rIj9mOqv/jLpk5KYvayx9rLO1WINy+fFNL3bq+FijYeBD2k6+IlGo+6qquXr5Mo3B+FOV0UbGHlB
PmLIIL0j0WML34+dC4HdsNTKj7AYF6mmzJTg2RFmRxBxzcj/6H2fCBNQuEN4loSVnCoTlAdeBoRT
pm9O9Jj+F9Dh8BAod2uKIiz/1ECFQEMJ6I8hhgajrQe0w+/cECbKKGNftSBdF0k03keNYj4twhxa
Ao7UkgVfa2YYPlO1x5/oD9IQrbUr99UuNfxVqYtfp6RIjBZFElY5bblE/zQbmtciVNKKC55K49us
6Bsf/Wi9FFQY4FK2XY4IAcfS0q0pfhjytcO/WCmEQsM3CJtZYY04fFEsN8Es1yra9PqBCm2BvPP2
OFNQCvxFvfxLCCX3Nj1jCRxBemRwpfkhMHe5jTJT+gRr5KHHtoBvIZwKeb+wglJNsni/5MHBC6aV
7/yXycZ6wfUYjbEQhamtfujLoNGwrGhCp9C83kFi5pO1UmCaZ9ZAkTzF+QwS6EFmUceM6DfC5FuH
UcK2jQzYRX7cwN1+r11sNo0n4YyMJ9EqIJrqG3fvN/cDMeDrMhJtKahTYfN6dsJC83VP4Urah8jK
Y7tNrqoQOctb8S3odFWkdSPOwtfg67yuuOHdN1LkK5ed18BmM2L/rZRjuHzTdyOU923Vf6Yaa0N1
m1Dpbu3PasZo5YMIHd8K4V9J6BOnX+QGDm8rZxcdRT7GxkIr9HDJH0ad6UmwrB72yBEP+MjcX3ih
8vk0/RPR1WQ+Jz0Pr4H1v576TK8i0WJuxkqjMn1mmxj+9d9jmm3KL4tgELc6I/UVv17RIZI7xLMb
1kMeYkILDSo7GFWvJYEXjp3q17qQnoSn+DHbCqVvhOdH+ApwK3gbgPJ7jUJgmmuZUqkAw1PjIiZT
nwx4jivTsUAmBwpGOwvDhO9yctDIA9ZYBlKYSixFMWmUXizH4MIJw8YhFeGXkGcCGqMeGNTYTKEw
ZE5cpV2dAmUn7RiHqym7mh5vuE2hbq07ISzaZEVqEFawufYZn3EW8rNVTzsEvrTKIP9OQuAcTXxH
+KRDI4R2zQVRtmQBCKRseG1jC7r8PSTwou3tKYFzoo58TIO7qi3VSVhm7pVCHQ83+zQbUmZf6ZEP
yGLgU0+OwtMpA6Xl6rYyQok30LnsgV0DGT/N11Xyn6+ZEmmfZm3ZEIDbLSHpAk9YzeU6XTFu9Z8T
0KKKr+aNLRxp4FSFZh1u1EZdDMBpRMvtR4WSXSzpBHelp5edguY98TLY9ASHbvCjQLHQIqGRRptJ
V0pe8bImIndK0+TFPh1lTs8Lvt7Ma32ufTxNheIllQaNkuHnCCg7P95EJnHSOsQdnVrz9IgFlZBe
z1or7ywUbTYP+LqiA5tlW7YnMfg39tdN0P/KK1/+PIPrfjBsVzkmyeYjiKYzVk+AfgTHZi8JceAr
FVpFi4uGlYHAqaBvOeSDoOyk5z3Cl5y2GhoORMfQ4FUgxx7OIU+hid/tUJT+5xy7hkmvcdFSVdzA
iv3ZluBZpoQj3ZaeIYJpIt6OwTOgeVwSyuz9jL96AZY7tMIR+0Mt3vBoFIBHCpXkJhfxvqC4M615
a4wWdoqwZzQO7cO/yXpwZ7gm0gZhxHhXgi0PUla2ixDG+i108/OhvNcST51R+BUgkrf7og8pXQjs
glbfyQsq4rL1CwpB8EGU5ngnH/XxHGilCmL/GHgQJIxeezEVWqnmENpJ9+kfs8RIAPyhFDqgGK6t
WAzlr64HI2sURP8nL1euGhCF1kLu3uJGj5pJIGjhHCAlVVNY392fVwGYUmldwpVTumjxkcy/7fIv
+PRMrjg5jLN545APDF1xElBsMo0wjGduO4ayEdT3skVRUybrhbbJqaf3fT2ZC3NFd0UNj4OH4bUe
h6OlZpSEv2EqIX4QpB2/Xy1VL8WDPIPcoWwnad8uYzVNXnr+Djaiko/ga3iiCpuHuhOMmHXDKbyu
6zZdHW+GrZs4mXPN3OYP1Kj3T6748A7+LuJLj5RUwnnYCwCE2YC5MBH2DsAnx8FlwXWEOzDgfx6p
SLtxIjlNHVXxp3GH+VU47heipS0qCChv5ewvb/6hL3MC/d09dGQoURiCs8ZpAHJw5BQRszk87ZS3
AfKdU4FfPcSY4zse6ZIP99U2FnD2vGquZWUm9bpI92cY44kfYpm6lLAShrf1Rbx71x/jngDa4m/I
mhnxzR19ycPUb/DYoNeWrvqtUAJUvILct33AxAEN00mzMJ3c8c3F321G4hGRGnEKRElbu6zgPoyj
e6FX/OEh4psEjJqBZVIcRwnFw4hyosSFAEc7gMhOKmZlyVd9a32xSIE0NYJVntPJbU8J1xZJl943
Ve1yyfBS/5LS1R2P+QYyyf98+81C1Ksrt1XyskOFAZw54XZo+9a5NytKzO5hn71xjZ4QwfjZjC9Q
TVitgNPahWGL8eyltoQ+gHMQZtxJ4ceL55PYKYNV6Or1WIJv/du7/ICjxuPLYCBKNRthhhmFHzG1
dmpO8OnFAwhtqEltg4YBdjUJ2qYTHfsdpxZLBKsQ2iuVfdKzjbOCypbnAtN0RIvDbnZffruZWHgF
LhDAJErFhyxFABUCcl1Gpwi84NcpwMmHvDHcsmi+btqa6baBf9sw4IGcRrIZQyg0ZBAV5GSrIs9G
6ymb8n4WPgBz7eVn79Ri3ErKaMQQZJW0AQz1R1yNanol/W9vdhOMDtRiM4ej8InJnRTftHauBAbH
Cc2zUpSUd58/CvWo00i0QfftTR7ItAKvBiOPC65iSWufsANBo6/kXiCNtpo1NEtnAkMgLI3US/tI
/e/3jpgWtNWw36PJx/cn3REwnL9SPoko41/HObcU/vXOP/8FYUwuKW5gPTRbVDTUEj1FH9mYM1Sw
aQH0M24SB/hZOFadPhv7n+nBn34Zjqfc4TEj1kMAPUUOLNuUIfc59Sq1Prmowey3qDjcjOtLNEyD
lGOOgOMCaUFIh1T4wyDBHExs5SjI8ThebcDvuGwtyKxnKqA0O0RKLKUi8jcSYEiBSX9bKT36A5n5
bqUlgryT7t2CSVOIJ2jLeS49PC0KpUmyERDJV1a3YrfQQVQSl/S5IiwsJVnSeRO7I+Xv8dRVI4GI
4QhZsanrMitjpgZKqVxchLvJ8MJoWykigvhT3744p5ZnOFezCGNsRZyczqMw2+2JNR+czTLfJLt1
F2xq4SshtLcMFn2TFyDKedpaK2BfB8nM9bIhl7/WkUedvpc52VrkV95Ovavcb66h+VUXIyWEF39x
DGL7t+h6zF9GM/uoHMAUMLh3yGLVVXn84Dir4E/D9CFIMsxvPm90k8TfsKWYwOOWBio7fLWE1q3f
M3TZYtlRzWAi1L8K6xSmV2q/YUlkEORbHMx+Px5z79/3zBd+lzbPc46IiJI3pvFGZFNTq/SzDWxa
7rPj185ujGfi78BDJVYmg3YUcKxyQ/yq101PV0Oe218BTTAo8AYtYA+XDWBYXFAaTR3mEDWm01af
wUj6TPGfsed+zHUGuEhTDnBPpke3Vr01lN6JtmnhI99vzMfN8HiKIKXpm9co2HguABzZ+/lAOdhy
aCDZLfSl08ZHv/b2CRnOdChViPimgV7gNt/VnjFFs4A/mRurHSbwnaIYJ3yExVqSFvvinTD5Nr6x
5nyA3CkObhLNwvBBfRL+ZaexzYXucfWSeZoqxZgeWYRxcB3aIJQVJxH0bTU6u/7sdbP7Y/X6BLIJ
fZpRKIUQAc8CX16aupEnKxQQsOPliXovitPGhFixhTjdrLyTKLFrZzb2LEx9v83lGAVQRUg7DHv7
xGpHLLTu4pMF/r3wXLpuaeGpKMkb3K1UoNHYNlfMZLIOuHAWzIJExsJMS3s6AjgjNskqVgekGaB0
YVhfx/ocmgyvfwzud+2beM6resp/K0R/jEeX8jvelczVRl385Zvw1IzGHQOEGFNn3vVdMMUBwDwI
BidD0B54rfLyAxeU4c4m26lesVCL/GL8Y9H4at/J6oCi5vhpVB5BgmUcvCmn+Mt/H8svY69lAzpZ
il4M5F0z85EfAKfnEm/I0R6NrMzLpFwsd6fVroYE832LPqbycxE7iRtFEYQiDCB1KajhM8kMJ96e
ohp/bp69+EzB1aHyQei4CDSIqY4fPp3a224INuSFChUgEKzJDq5a/Uf3+QvFsirneEOLNUL/Cn8S
A94IdgXJ2/buI61rNf6RPJFgI0stWJjOH4XziNA4tiPMo/dN/kb6TrP9LaHqR76f9fqDMMApk0vQ
VenVOEMIqfiRTSdgqDHagj2EU5mCuzlFob29HjNR4alA7kSkr18TcJ8qLw9xr64YCGLXAUL47nQ0
GOg5s5oaF5Dl4m+o4gXOQT+LlCKGapev103xBafM/aJwNsAc61ZvDR8yIWbecw+cdzg3OszUIIxe
5wJVE5k66Ta5s+wdliwOUnCtSOSR/4co7LKQCZKR943pV5dHx287Sh3JYTn7ddQJKRd8JLIOK/3E
YF0mJfoPgjr8zFTD/ui5p5Ovt8u/Dy6XyY/QkP1redLw+tRCUrEv+AncFsv0IjVQon86PxH63EXz
tDEevXcWEL7SnucbLS7X1PBLjS7+m428uQaBHHXDTmStrHClau89MT8/46evgqwa6wK8jRFqyBlx
mvpkqdTAL5mMPdMJWSAFBJ0tRNNJG9pvIoMOf2/kRpowy2l/Dalx8Fh3Mth53Rz7UdJ4UOrUJeus
EHpJmyIymCD7nJp9If4up6yskY9n9N2Z5Z4OyZ6KS75jaMAyNpFwj/HOAG097ua1DKxy0A5tuz4X
6xdyQdQWLA7nZMDUtfGMWlGmWxibzmxcuocGloymYJJNnNXvphlfncpDLeoiftWjgzT30LAHIi3f
0u1jQ8c4ujEAIqSzPSvK69EKgHUwrSR0PQ2UBxaOMzioh05VPekmuXmhHKt/o75eXMJbn8k35In7
nRVgmb50z1UgtO/Gqb7TP/rHXD19oyCPgXbEO02Z8dD/Hh4vpS9q+/vpqy9RcwBcxDRwio1Q4iAj
LFFf28qee0k/gBycTlE/1hdGKE59SFV4XmTh44wslKwtfCuu9HRuML1ko112bS5M5iqpTUUm1E8f
mcDVpxowoHguqHis18ZhBA/edagypcneD9BtDo+damNgALTC5/VPkIUJj+Xu1ERXyx3maPhUq5wE
nMrV+rIEtdcwql5Lfn/Dwdm6PuSHcT7m4AeBPHe2XeMGJ6ieKGqaXf1BjWgYcIhd2j8fehCd4nOV
j3fpVRr07wI87LrCvrBa2/gbbYWhRfMakc8bV7zLgkSotg8mVG4AFD8anB+l2oHwU9xji8do5vB1
jcSQJxNaAdYQ+SDdLfR17LX/Q4iHtePfZ1p8gbCefyboitU9Cm/yWQ49r9M0kI84/hEdmd27ogPI
qHffOHihBJ0ElQ/8rmeb7b6B23xOWh+z8D161NpE4xmRyARe29MtNru+Ug39ylhwyJYiCa/1DjUR
yFk/D1sCTidSonVznFy7i+sxeb1SH1ThEEVdvJaIxYa7YnorxpN9uD0korfxFRz3smcMfjeKLBe8
lXpqRJQmgEtW5Rv/ipT+Aqydm6b0Mv9S/FD5ND0Zun9G9+sG1TyiS66qONquYCzmciZy0BcmOOGo
BfCJJXd7lIjApPwessRSJ9HxY6eGA6YvPBHW/w0EqAJAfK7FagaDRW7IPN0a/cvlrSFRtKOBij2r
KgXkRsrYnfRUP+yr2GtmKPl7/DHnWgB3izY8m9W8jDNgWSpLTjb6QOj4Jkx+bV0jKJdfZVTw47Fn
vV7u6AYYKsx1CixtIy3NNwQqsz6hXBdtI5qKvClDKWfALyG2uKswveXzKqImosn5PuhuWnqob1Qz
qggOrlB1LkYiXiuhl+l7st+u0dh+vOzdS78yppbE7zOFES2m40w2Mv3mV0VsG91uIeFJ/0wDdXVJ
xmbmlt2c8cqda8l+8jTGVTTJME4/bLicpb1lvOFUSrnljkCNl0XAm1m6aVnmK4xycs0DFfifze/q
zde2Q76pNmkFidpglymTqhPEpaPq4G3dQZpYLf8r8mbHJ+xiAj2iwvNX8LDtH0TaOX4pcXFmNpVM
0vFBSq+kLKP1kN9aAWrQhzX0j5c3hZ4O7RR4l2Hfd4oSUAGuMuB3FIaqYyotmZhu54oQk53XjA27
gSy1ii17amiimINxM+1869fwqc8IquWg0NCopI63FRsnFzcL9lqZCCRiB4qNBbk4Kd3OILp/E8UH
ZSV+kuSMWezqnZqnNwZQkYkaUsL20L7/SbIID8sT9RdZeON2dDjMqfCayOQym44qsIM6Z1+MCH8Y
ikDQJ8yGnQX+bDCSEOHDmr+GKfvBD5eKMiz/i8/QTJfqEiZvVQOLF97I0MhEJzRXBOc4oNYNdE2T
hLSg97Y/d9LAhxRiKxr3PPfxq09pTYOoQlsOvJ76Hzb+YBb1GgTIrIutiTK+pch8eGoQ64g0HNs0
HOx0VmX2cAJddxBYCgD3/jlZJJDFC/LSl7a4qC4ruX91wjrKXADSo3RbdFCHMVUbj4MMrfTfALAl
UShm3xVJSbOhxdp7gOTw5qzKNPKvuVrerCWtvKLE/v2ib72vWQvmVeRLgimpj7m8Ay+XHAEejvZ9
TDinEjlz7syiTrDFnKAzAN8HHH7AEcwChwDzFejhTcmmjpJK6paTRIaOjpD4sfuNCURGT/+QlSz2
ZAv2O1IelP8xV5dIAlkbi90kBTh8Id9rA8PeitKY+GLdA7THABA+05xOG3Q4vECyru3/BF95Nm+U
l1wd1/l3UxT3v5NYOS5FiQypx9X6wZg31Y8L6EqQari3krciWAiE6BN3nH7gEpR+OiQpihvA2kgE
X2Ifujvx9f3dnn5KhunWTyFyusWp+ZHj3URGmEvbvm8lxwDxPsDIjJhCiw1jeN07Px4Fq4kL/Z3s
e/PbvACKlpqfNyHvXwqpPasPcckrUiSTlYlf/I4ylE27tH48vJHCpZ7YTE5XM/ja41G/pDT2oD0J
4+KNRgnBw/xYcddM3Eobq/7KEsIeL4fUplY6pYuV90n7qyJ7TF3z9mlSSL2WbCXrnLcfw/vPQ70H
09yumiUy4ohMGZH9qOiOjoMcwGxcnlJwqN/MZie5YkPYcRsE/pKMVc+iw6BD9RYCReOtadnj/BsJ
jlLTqa2CKKi3y9I7Aan3l/AK+qHBmGrx/+SEAoRFLwJO8t22zJ3CM1a01+HM1MUm4cnpdxflduMJ
CwWHxD2TDTP1BBr4FUP01RcLUSVuAxgvmmmalUvJgUIZ1JfpYUyVt+ACIFV+MK/DniGDf1+s7Kle
Sv3pOWCjZaeECpOibhnXPDUeU57fPy20WH2d3GihlabWDAcR6rXJvRjjJyc8Q2+eMD1xvdS3g5ZM
I0DrewcZofOkO3n2SdcZxhnYO+9mMp5m9AOxtgUgkChQ5IXy9UnAHmTkFi/AypyGEqgtNZTl+iyd
EpIkAHAtPrjkJxA5eZ4OR8dmiq/CcGuib636y0j9Y/PiIGpyeXEoMwxbpcfGoTXpq0aIcOdUwjkI
9ibSFgn6maAXvrwWNqXeBWSxXfKovo2XHmhBwmo5O5na4VtoVBu4ZIMx1r++NeHq2KXoYNTKSpzx
mm84X6kf5r5hV1sBNAAR/7Y7spTpyRV0SZ8xanV4qXCBxWIS92rA+zgJxXHbGxYm2cKm3inPJ2o9
eAkvu43zmHkCEEWQx7YjhdedC+Zw9VbdVzVy7F4hi9om+7eU0ZaseBPoGWNFj4mVL6Dznfm5NKQw
mzdDc42FNDi4L/VaQdfSxoHHyKtAQcC6NbrgjPgTQKsqgyTW0TkddxronCN+HMoBob+qogf0PCpR
Lzoe7+pD0IQ4uOTP1YX80U5it/a5IzrfZK6ejXc7n3kTz4VgY/+gzomnP8poScUWXFXTAcEt5piU
Bf8WYkKDlRQmA4BcJ6By7HhgZl59rYofFcPmjHRvDqxsxgdZGST6msfM9tS0xmPbx3tLeNlI47UI
dxx+9p0H2S08tTkr6ioH3olWKFMaAUDEBdchB9JdHW1WPFfJhUaZoAcZ141bDx+lWQSeYVLoPlXf
ExJcO6j81/5BlJ3XVuBdtxFl95FLF2eNbCtb621Nk9ybZjTVFvuE67e4Nb7rrSfrqglDsosF8jsr
eJenhzFaYNoCSrP4o62ZjKF0K8C7iTl0SKiKiHWJyCkgitevWS1Xf+y70xeYJO9KV7gUlvcQtV3r
MFpqEh/bKdcvE8lFTzoHchKnhCavUBRik5mSrJ/BSWaZYkBhMZTiOtJLzs4+GDFfZSRaXyyJbu3s
lEXMwTRDXZhGQjDeDBA2cI495/Q/4C8HCiNnJXgzGn93HtGO+s9UFRtvpPX/LF12t8LMEsG5Wvb3
9Qt/QCgu9oUvTHGgf2pYl+3WLvzmN2jKMhrtgH1FWLyjg0cS0DrzKl2/gXuGfA3pdGYnwSd6L+/X
uLTA+lM0DbB1GWEnMXKiqocNgBsTaH3zRd1ocSR06iGODaJLqCewTEZqOL/mQgA5/H8hp9wFurd+
ZCpCG16ZBSHDSOVID+8TUL7z9iH9CCYyIXknIHSe2IQLvnyYDfqUDHLLhvXX5L3+MsABAB6qHniy
IfoS5p/wu/2ZDSBfqrVVrzTeQGyzVlwIqlxL3CwqQZRsr3l4uDrHNZ9jC7fIKyxQUMZx0D8Dh2YQ
J40fEk/H+qWJRsou5ghhakKNuGNP8FGztEKQmZpsoLQWr4KkhgK6vJ5o4TGcYzWQePF5TLq6MKqr
H+CDsAPVh8+bR+ecmfeTPdYSo3xZ05Qh0mlo31pADkWIY1092MLljMB9EGDfjJtztti65j5X7X2a
S0TktXE0ouNK98YQ/7wkIoLRfO8NFR7fmrejXseNauzepWCRSlQHmcNVaRTGRV271vLOOyB6D69g
68LurnmUxMH/lxBTxq+FzXZ915fbwn7iNrEz/3nphRw9xKoWfaR8KfhsM7x3w5SBdv5eTnAaf5o3
ybsNpf3NXNLftCKf/fi1RkLFHH66XUb3m4gEIPBvBa70C5+RZLYv8L8KNyZL/Kmw8TY1XvkXHuGB
no6uezFv5h35DWdUclG7WRfR0LEXmo4RH4mpjekr0Inh62UQNgOzFcT7IGK+Y770gaIATfY6c0Gm
iFnTBkoZxFTBFEYX6vWEhGp5DhvfNxSIlz1daCLrgEKo7knvmMUYp/wvjtSdbI3+i56A3Fp5182f
e7Va5RNgftTyNAlPPFjVZs2ZozfwJgsWGtS33nLVmOX+h+Hg54gu53YsqJ/A7auem04c9Ttz3wq8
uK45fnGYb0bN/y4xCU0vOPj3XS1UDQZm52mWR1IpCXuQ9Y8P4drjl0MdqYBBZwBwnLc0rb8I2CjS
Z1Hm1vPpHUdimR5rZRkliSwmfS649gm7DSRRvIqDCN9NvHhmZ3wNgWBSYIefdsYWHQ4+hRzTby3G
r0XCF3n7blJPXSVzWmpT+UmVHZfLuUIod/N+w4ArQZMZDw9ez+xH+Wzw9dIqt8MrijW5HDZFWqOl
0tbFzUQvulr+lKMu2E5a5ure+GGyTxN5oc4We42Vxw8E1M+ZgWzSBqes69YVh0OLSc0VRSNWCShW
NdIExCamWTNMwSt3nLZ0Z5P4ZIZByNDc7s+XS+ugl4cqPDAc3lhmhfg3OCrGfE4CzBtuj8+Zv7J9
gQjegB1be22g3L1VXOpkecmBM5O+/qRprENmyY7MGWjN0pmMx75bCLbsC8D4Z/8tqkY21eV6WPGs
61TyZtnT0qcebwqKW9F1mU1zvz7t90nAG6xbNQ24SKcRXvEv05GLJsuQj1rUsaZgCWuPmsQYqYx8
/GwOlq2tXBmlNgpCGhl1OdBIvmNAOUOhiVESr2hMNR01aRPw+74umZxVlgPqJgwxWeG2IuAU1Uw5
wbvUwhVJVTy6yxndRG9utT9QhcdGwvV2sg+yAbNXwa3y/w6dueKgOwZ1wx+sWrymCvO0VQgONzAX
UhTQKxUYeYDKyEtoqk7RxnGk2Pz4My3fosUyxyTRgsB+BwSbOiiJVn3Sy7KX0QJYYW/pnwnEfB1g
Cna7UoBEMmuTwF2U50yUcJf/jQ2BmQqGhRlU8/R28ilbg7rEEh0z0macaIHDTNfzA7urK/pYnZ2u
RVUvUcwXXxvqcuDu0LRohx8ibBYPw17L4nzZ/TkTCLupBRRbFsvu3L5TUGTztEINLIDa5slwyZqM
HgDu3r6P7HsBhrHy9J717w+wMT48fptFOeUDi4OwEYvuuBPqhk3aC7+V6ksgQsaUkv+YkO2DZG7R
mxwyaAVP10tBEMZE+RUDc+QFGIX5O1TzhvU9ftk86mWk2/IzoJx/NlT025RP/W+kYaK5HP9iVoDG
uUalCjpcfZZ6SyFACmAAJKH3FAYcCivP86aryfRiDAPxPsmxBFHsKyY3ZIS7K77Lwyl93LrLQPgz
B270F5SS8Xa7ZpsWRa/jwFSzP0PrjzQM4uxxovAZ57lhWb03M4xuegr58mTio4pIkqvG00DFp/0C
JDLlyYCCBaUFlT8vV0nsyVc+jmxp36KqPUpO+uFeOaXpSaIAGXKHfbo/Lux1S+d0GBmefQr94G6c
wpq6LKuq7gSBB5KvuKLRxQxQBc2cGSuR55WD3pp0/SDoY49vOjq+R2Q6Bknyb0PHhILApwecRfjn
icgbbEt9fYht8NFa00MQdivy681ush51ah2Xl0uK51q1zTuP0+4YYAyQJmeV/JcwdeJJd2t1DrPw
NLBXBQXe6Nznmp9CeoOsJjOpnzcDz1rNg3E23XQtEyaa4DAlvtxyq+kB6+xebjEbtzDWzQ8MtCiU
sJu3DLW3Ksx4lE4uFnTAY6VXInWEpwMA/YiPNtBxXM2rfDzBO/q471q5Jga8zMhIl89eoCmCS74Z
pwGPMBu/2NLZNsv2sGdn2z4hX3ABZaMnF4wLhR7HWFk+vwBsDyHPWbxIZalAueZwXM3ldUW1mSQH
itEOWxgAMtDXHyZah+irRxOleBjmEqTaTFri4Q8+lwmwlwlrZC44bj7xzNlHRM0rMBiQtp5AxweQ
yg72TqbI1mknEJfT/VjXwCXJyY7q7kQlyjg3qaSMeszAi5Os3Dj9/vE/wV5yM35jfz4Q+uI+zADs
UzCzS5tUbHHmkOjSjhZ8KY9RhSsiJD4+7Zwp0jZ2LvNgB9JiNIgqqBa7ibm1rgS4EoDV1qXzJPfC
OXPWY6HNH2zZ0i+jTForH6QKZyUM0pL8kzIlujd2sEG/jG5ZiJsiv6f8G/tH80r9k94KB24+CEQj
Cp8tnXCGWkXf3FDrTVmBsXk9aaBZrQeFLOj/I8fmWO5tKuwwUzH2RyPxYou0A9u8WD1Qh4qvtbE/
0MDbOWEb8pBguL3Of7K6QuNkPrv0FqC69EK9qDu5sJ589Db22W5WEr66mpesw//Gb80rZT29cEH9
+19Y/GxKIyl3WuiKv1MPa+jfTfKFWEJ4N+R+XYFnRkplo6RN/BdzoQmTvCt4YNU5BVzv008h8ys1
9+thRsmVZ0MQ/f8olToNgQhSWQefkcj08z2hdm+laBUNn37Bk+ZiHFMONm2VuGbKkAFTcmT7EK0+
NytXNANe1X6BWosC2SnSjvCg1CnMveThVBtKQszjDnsJs2x7yVAu562qHS2yyOoXhbCEuFwscdHT
H2XVdVd4espe9DOEEGSMKMYReDm7GvXedIgcI6ckzHnJS4AqHt4wtvPRREYKbujFln+voZxkuNLx
xzUluORk3+eK+qNRvHGsnNjeyJXHQEwBzbo/HvyCnb8oD5oLN/jNjGgVT5hZ5RcFWNlAGUZwFkU7
YCLU5D9VA3GxfSUOiGUHPAUeG2D0h6xq1vubYAD86flLBkho/mvoZDETXEB19JQ6akhgVeonjSxM
9bhdPAzbcMlrwI8LuZYkqB0n5Fvddd/Jg1zHTQiO+dn1kr7zjVj3c9MGz7iuldHHOHzhEumFFWs+
OVzbr1pT8NDyxiO6Z6X3g40nMyD/oDhONoB7sbk/bAp1vNfjS0sNyQqeAbUXDCQt3BM7uLrd/9Zd
t+tw0BdIsAFW5q0kIk0ib++LVvBFeCV5nrhq9I7fkjiByLmDsTAb4gZP8yj2gTBfU3EgJpBp6kr9
UNAxU7rGDzW7RdQcA9JWFhtWy9D2JdhJvkDWaogaJtMF9Y0wjV75l5E0lKEkSH6X2qpU1S1DUN7J
OJYZKy5RCOY9O6CP9LdlpX++AMr4c+Xk2ugDwFYCbdHLdSG53h8lg0sFDNU819z2yYLUBvFMN4kY
HXfBaFbSVhj1TADe77YH2/vG0Nf1WdLDRj9F5ph4u1JyNl/LkCTGrmB7MXYuKDJLS5Z1Ogbuws5B
Q5P0iEH6ZA8tvqBiNKXKgwwsezLO493Roi6ceNZfHMi+LGf/8GB4I5QY2HHX3Q1/kJOYHSanJu0q
2f9KbFlHoh05tLycbr4gKEXOsYeGdaRMNOe4aXPIBQwv+GJ6+L4P16ZXzuE0auV5V/E3saYq1CG5
H6D6nToU/84d8tfcYrjrL//at0FvN2/42bpLQiwjO994Oz0pAgPHxNCz4GgWBEtA1riuLZTdgkPK
g4L4IAcN7yUadCopW7ZgLlZwt/8GILrab8xSaZB5rVjJdaAfGt3k++RKpU+rYaPUfOJlrnV5kl4P
8MqphCZqRHNmD2ba9ebh+RK+YXCpYtOKBdUA+hL9fWZHztsUmx7ZURcg0HrZt1zlpdkvku2KYOt3
8JN3xc/LabsHXnIes0dQsIO4RwhaY+eo9z7YScsfrIenTEq58W30Wob++Cm12OUhi8PJTeNfS2U1
fOzunZwHqwv8TVgpP2pu+H1dC229xpbYanKi6kG8HB4JetR4J6UBOVb/GcF06gZ7vpR3vP1xCMHV
ibUGf4i/pJLzuyhhYxdj0H6REzPf0lwqFtjfUwLK7mXE+UlL6K85/XolGPKmMzo2KsoiaGCSDoBS
aEuR6TJfSRfvVI96zdvV9YZaqe+dZr9XnUYAYyd41f5ldwUbRp0kAqh0iAGdU1X3g+KejxnmnPIu
KnlHmIcJ53EbJZvuto2Go3rPe1wueZr03Asaes4NUnzhPDfhlMr62UzUJBrV9Iug0AzGE3zuyXC3
j0pebBJprnKfiRMxUuy1QBbWWvlEaRWwUH8V7bzpMPPNk5nFaXJxPjLB8bbvgsbaF8qRlpgXym4A
sZcZ0Q6IvPUWvIRNXvByQMDKovsrmjzA5Hu5gW1kz8gTWIfPBkzNo0wDCMOgXYTaXsQOPbtCt+zj
s2bJu/DDwZkCJTshEwXCHu6O+I9p7+OnF0bXUQ0jLR8MhmzrR7177tUJwS4nBjHMD0WNoj4UCi9j
6Yu/lsentV9D5O8lqpRy87e9FsrOknE2K3fma8niXZA5jUsolNQdIL1UIsWJkhjZ9rk6UtWVw0NR
2cqM9Glr4ozBp86dI+/5+RQCckHDt2/JSO7EPXmdx7n3ee3LcYNi8sfTl4HluuSNY71euI0udghL
ikfNC5Bpp5WbD/+3XQpC+8qAL/uy20pvH7Vb81S1jyI9xnEMdidVTC3+FG24P48GjckrQKsyldnm
FsCgYnylfG6j0e15diVVgFmfVizgivnNqTPtT0xRA+zB99D9piLwJJohyZKLjEiE0c8ZVRu0ucMI
fV2vFffCKWjyhq3rOOC+NXaaKsZpSQs5R25mxME696A/aS9Pj68YuDIXav9ZeW3NM5qQ6Vg6dVKi
oAnfE7IwnNpMaAfX3MhaWEjOLbX9lvyheBxSJu0gzjRXSaT04bZBjrh19I942pvtSyDzl5kXTgnA
anpaOh1iOusTIOJaolGz8dfocxEgBL4+mP130rcdBH0WxMV+crS7xGf3ZHcLFuxs/FUcsPr7qQ0z
tVDPpKyXw9H3I3f9ZOsl4HkaRPhFTWpTBXYLIXdA+AM2Dq9cJqYdQD1lapETh3mUeX7VJ09yFxdL
bs3/CD9n3Pa1R+MiKjExwb0pzquqHOBdV5D3TNpuUQsVD7I6o0XEMAwZowNgZ9VTlxrcb4hgRjvL
HFs7ntzLwbIb8WGZ1kJ+jDWXKVGa0Kxk3IfcoJzF4FEuGwfXZDp4hHI0FcNJjzpINmR8+v7bpzgM
ANkHZiDm5Zz2RsBoPozUkMbRrqJ0Wu1v5R6PzD1TlU/clz9CLR50lLh4F3d2ozoB07yg//WbRME1
L7mv27opOx9PG8V5K13bYI736tk2QRViQAHLZkaIV4akeROytstmdSH2AHp34ejSDK01pIUIv+it
EWJRxROkGAuzEXp9tdX5zcCFnpOsz54cgAtuPjNYHdSOhCh1L41bR+o5h9hvb537uropLn0LDoJW
TsLY1dJ0sXz+0JcDnxVoOrTRbCpVaXWZp6cfFj+Re09IK1Q8MUWhrKdRgYRyfzP3To+rNwMWXbAg
LnIE0ivDp/Z072UiZT29zNxCc2KDEnRiXg3tD56KGT6yau7OtCCWMYar7TdIASRSbLnU5NUGMTd4
1OS4cqF6S+hugM1nEELtP6flHVC//WVgLqxN0f8O5SYpJaKnYti4OmlSw98hSrR9vpP+TbMFfOHc
uf4QdYizk/7c7n/g+uEnAzhfjnblOBYS15Ie5dobgJ9EhuNlw35GL3J2xlfX6UBhjR3muvci30ic
3KFMbOUyIcSPRAdpGSJ3iZhuAJ2HdxyLg5faoQr1/uV/4GDWcGjYit+Or2Guoe5KnI2xYK57R6jg
qm3mfpqc0cyReCt09Vx2tI9Ifk6f1n9rof/5N6GrS163N/XbAIf3PIJznz8rlk0YCNvjzPYshnMT
W/rsjIFCaMuY0oBzygFSOMXDwyBOMhjSqMFlTdkCHoJ7o8oqKMcP/kqOdkHio2e126BalVaNy/Eq
NqcRcaFK0QrzEXAsZMl4EwlshxBoDk47/qnxBvdkpyR8yMW7I0Z6tM0hSrn+ZmzfQNURs1GDbUqq
fwR2k1ElwkI7UyJ5Mryqm6tnsdbd7RHAvNOLyBErh/McEGjPHSWexmqfNjnbihzGuruxGXnQcYoC
YgDP4mmhK/24NccciLbSJoAHg7MCTydbJKcEqiuyYAUG9x6Q4mnKnKk725Cfg371jNaFAxIh5HaX
gUKE168r/rapoA/YAJ3h9TJOURNhjkh4TruuAQaDvDHmkTpJqHeqydf6xraprqnaElzZu1fRpYJ0
YVSin9lvjjtITIaX37NVs+wc1REgyDmIwiDhIVkOpa4S08BBuzV/xMhEpvLtcJF9JseUuJqDa29z
wgx53vuaYiWD0PcsrKNiw2T4vghVMLbov4wOOrvx/2jQczHn6lx/cRFQImpTwxpqO75MTDIX250Q
0e5LxhcI1SZR95iRqvFxYhQ+uS4rd8FTRTOsElAI2YrBrApac67J0zHgSIH0a9YS8AYq96JxUH4K
pzFL7w4TwLNIVEWowelb8FPzTmvNUBTYmmasQPpWgm5sG8cRl0Fs1FeU3FidbUdPpXqsQvZnpSky
XUgFyAj9jnaOQh2OemVSwayHWPlAZXbcXZXcmmDe9Kqf6m7fYmHFBllZe5+NHypSXbLivWBhBC63
G4ApiCk5eB/cogjGFXx98S6HB5PVtc0Sd7Qumn3Dqat/UqOgQm0wod62MZaRftMfNp/Qkb1yX7wp
Po/w8uMZznvd0bSGFHpKCOPApSi7ytpYl/9ck1CZbMMNNNuwWzB9SgSYHmBXKCShwIUFMYnijQlW
2ophsRdKhYlqbs5KgAGuh5Qsvfoce0Gl4/Gh6GO+gaBJ1L/q4SJjHzahKgsnOL/z1LqkR/kvb1aq
GNRE3qzGZhPwNcBaBdUMlN0OWbbmdOJ73j9lcxb04TYbj9Rod7HDcPn3Lthreg4qNXGETkjOhxy7
PdF/I7Qpp39z+ms/YD767ZFuxyFHh3eiB1WnK99tA2Em5dRg5RMAaiNdYx2goC94nzj/Ul+g3lRO
LBPnFEL6eb4xVTpEWFfatrVu2zHPGLmuOm4qlbECRjVfyJX05EqggMqLd55M2Chb7hwWNRdIg4E7
AsGPZ4WpG3sEkctU6Tsr931VCGYzZzBt41OmPrlbY1MX3u+gDkuU736QxsHi6DdDbXlvIfG2W/X/
758v58PJbo1ZmK8AAZuEdu4wfmXacYLAGhoOSPFKE5D8XebAOCt9HK1EhzzDwIwY524a5Jr2mUv4
gjzAayPB4spMum9pl36L2zYwiyJStvW7WJRZomKranvApMzVXP7v/ecLwYWF4RtPQvns/i33ZDXT
BjvZxVYVwVOl75eL6aCA5XJ7U8rCpFydechFjChwsWHPcJIvcyvz0D5dHCGX56WSFIXyAElpJtgh
i/HiDucbnqt/mGf3wkeia9B5NFAoG6DEA/7KMg6O7GxF6fVKyJCNnzko0eTCutobSf9r/xZwADxw
YyAdB6QzWIOGXEH/Wyr93wK7D5AvySNdT9XwC9s2Zw37Ap67PUlJTYyMffXsrebbJPtUdcCxhE9O
WLlCvaphLlkukUTqLXA7axTHkX9wZUyWMysp2RMOHXMKnU+SAzT8bGqd9RVmnQPxsZKDqkO4n7/9
J44bOu3VJOkCappdd+j3cKwf0ZdLk1LzM+EfOJvL3GuOsxpd5j2Bk6y5WQNsSIDoattatzNqLY0Y
/ksFMwv7jkmWqSXvvXbNQ/nZmqg8LYpYQNNC3IXmqSmmgYZ8GS6R2ToE5xC90CYN6Lkd346Ye96z
DOYh3yh1QfOWuWYtU8rDPm7jKpS6JldEx+FlsPyU2xqOeLiUNXPN+g+xmHIFZjuSvceppDn2/U32
G/CMKJKhLQobSmzxnOxJDyRlgR2VeBKrUHC3wjhlG20+1F/VzKB6FY8BGoDEypGGZidaxyktG+v0
mJVYQpHTRh6b7BpB+YC4Ez8vISF7OrmngECTYP1ySD2qmM8o/52eGPUa983S+WdmLEcID1xE3rZi
oA4HTdso0GBy1SwfPsAdaHYij2WIvH18/oE0zP8incUFpCFBmKXcvBQWEi7jq59mZ4oHYVnY3Zbo
ulx5090MiqHRAdXKgMB2hLv0YcwAtLfV5jrubknsmim+hym+a6yjrKEhyaDktuvDW6z47IamMcuL
JGguBL/NXIS7d6r8w7Fx/dLkjze50GRKe+M7p4SjloWAaIgaql8LXZ6klhx8CVUIq039DH/Nr736
unJQ/uwIs0VAGiCgBmk5TkJXlqbgXO8gRK7qRofmhoIJdJQu12paFX/HZeWGZNFZUpCk+fM4gYJi
X1o/xg+aZjDQN/Izbq+Lg0vOyQOEaCyNTqLobDr6K6hw5Gy7Yd7saq8U0+GHdliFz54TObejXE9v
5qKLKWHuGaDOibNoyIlUDtSNJPXMEzipQP5G6myDAMtX1G3wbDYwi5La/syFNxBodw+vNbCD433f
Vuedj0Dxaaum6rAbYF0MIZxe+HbcJbMBksBPVnAj7J0kXTdRFLVKZz1FnkdPWtV6wGEffaMOJsDs
W1HaakDfAVE5got+Xw7LOLIm+Aa9bs3lb9nyav86rjdQjpWsn02Bz12szQzrtlmM/eM8GFukVPHI
yKvNE0PCAgUhGPK3IrAEwk9eNOOSVplrh9LUcQRHx396UJnXVSGu/zWSD/qcr6b3dPzX9+rNgHOq
hUXW/pf+CSb9AwVKKEFOqhzcn+g1uSNaE4n+bhS+tA6SUUozEuZm0SGrZlxStu2FEZOVycPAboEC
pIExcktGPIduJG1XDyggIcQcHH5VddxddfmSa1c+WztsZXGBCssXvfj2DeRxGlXAsgWaPJHDLa3j
K3EzdGcc+OoT8V8F0npcwkKkmnnA8LeN3fDLuU7KLDwwEUjMXf+DOacerjPSJmXSJVyFEdxkWzEL
8L7GsQRFN0/eJiAVTYSB/I7FG2v1NOTR5DD6lr5/aDRd5krRCVwCIkBpRILZevVQhspnBcOmqdc4
KnaH/rBr5YMd8OnK3wJ2wdLGsYDe2j2r1/JYEV7fjQvgKiWZcFCkOKGt+8tdl6E2r9qG5fQ5A+qo
ZF0WLv/tgBJ9HvyUJxHhCXvCwyNl1BqBqLKkIWDOVjrglEdD2pdYjroCpX6xhS+xXYDDo4H+dO+r
APFs8eG/UwFaGKlEaFe0mLRFxEBV8jZiRQH+2raftvocWIJUDrDwkXUp+zNqaTtDaibNC++h6A9S
+kuHcgN3ffxtUBybIncxmPtCT6OHV2cpj5RBOUYUcc/fFibJQRXsenkH3yDB2bAPHSV6wzGPsEZw
2+IXxy8MvcAE5iTdZ3JpWmCoO3v9lp41PAKm2+ZAY4LqtGEYMwcdEW9ujKmiRP3ZeaNL7bsFAy5+
+dOjOcidwF1hW5jfV9XLqA9AS6157ye/za5kS/EVUaTCpKkXW1UlFZaOrQfQuJbFe19+rQSaA+T0
VVzv5xNDuYfEFMMXo6GGkb8liBdEOnJ01UVEhg4XMg55QAKUKUtqwdlV3CWCSjazgd6MYPEM93BB
3nm/92wQwIgokHXphFvXL33LsmZEpVai/4V9n046xwtNCmKPabzqT73aFyzWU9fPGcVr/Vn9Ucwa
KfBo6V9KnQiyJlv/cibSE6KkHkGyTdCXL859cBTNJUiUKKDl5XIQKy1CRf9dBHUtoFHjLEEmQRow
OWCVfWk6ZteLSoYvhL5S5pDahOhDEiPq2/XCO2pEmKKEkwEzJOM2lhVrl41Zjd5Sf9t0CVdhMESb
+b3DDFr7OapdsCOLBdMuOtkODiqMpb2ceDWMrylJ+YADgFTwvkFlAaBuWgudwwuf29TSmGAFkEFk
oVEBQwu4/P1KNgXJxX+bchnY85hW0HAv89Sbj/camaEonN78poYfG2ZZAADvSLcjzvFRyUCzye+0
Epz3MaEMjZ3GDgIfP7+fqMGdj97D6ooXGeMj8SG6Mip90ubIz5VEhACRQ0t6rcjEFa29DncfVfja
RShsjXerCGIfDKRMalpEryVUnobJqYl8SQYlEejBuJ4ejrB9xITmIepuyBFKCiEwv33t8DEd5TO2
do8m1id8FUyTtu4ULvt2Lyq8HPzQYQL0esz/A3NNIob6MUJgEdW24f6PZ8LUYkdP0jY9XKo+tiDa
vUKBGGXOavUIdhZ1v8wCght9lKjttGyLo9JIWTwEbQz5mhxKhB6cE2ySduO6IzAhGh5Ko7HlpvuF
6dvbSPA0ahZWg9WmWSQeqGsN3JobYkn5zbjL3k6gAr0bWs3YdWQE0zKQ39aZqSqSWjvNFYbMfhNj
vy0azIfzl88xOsKqlC8xgCKgEh3I1qUznE2zcTCJoqgUq6gKzHVHQj4DCqdsAEyGYP5kf2+fi+Xl
LRD0C6QnSmr3Id4/B1a2TsQTLZBQ5Y7Lerf2+Fz0YZtzf8jYJE040cjdOu7lYelqFzE/k/gWShli
32udnbZiP1Ez7XACNKWv+6/cJCUyZhHD4sG2ICLuLe3E8VVLA+YEqZpan3wS7y+bACxFXVOrzrLu
IaRllxjWsmcJugWAC2lcUZJcuHD2TtaL+mFlex59+RUdNEXky+5H6mOHsVE1vMuWSUa/yufwzvhc
PiZqZd15Xc0t/HMFmvcmV95NtY6f2RZESq/bUDHt6Ii2q0ERIRK1eyctN46B+xq3rjTah/nS9sDX
8eu9MgEWQY0ShiUOX88lSlju4uJZSTYsBQIOeE/B5pZ1X9ah76PMuTgv6SDIUNaRzks5ISpoJUVl
uu+HXs1LVC2Y5cBxJXfCpY9WCQhlQjdc5rcXfzBZC9v10h7FjTorutWY4wpbaDMjFQI/0PRNhn2w
gIs5kBhLtqaiiMk0705svbHsUbp6msxvvcWIWKbZERGZUR2U5VRoMh/Naq6wuDmFZLWyx6EHgmlD
8OZ8k9qXHpQWDrtKjXySLPCl4FRhe4FRgO0Ytq6T5Yw3jhwm6ylZDjpzmKa0Es0N0hiMdW17HTyD
od09njXqoEbcXbHgffDEtFoEkxWJ7NSCoyi7rfKT3031jg7vC1jn0fr7RcETsgsb3XPR0HbMznkn
UDXePTYHhMr2kctJ/bci2TSa04Yb3Rk0Bbdn5KeJae/6w9Ji39LhBAZ8Ko9/WQWEZ0pGeTw+BKfV
to18AUvRgtaFd7zxSA/po1F4k1UM63UkxZ3Oulkeuks2mHV7ETkz1nJvNIGWYuNXSOJaGhOLSIu+
/cjqTcbJfGBgB8nmwQzlQxiV98pqeiXB0PBv/2Bpm+/djRih68OcUFZQWP3sgkldhGGeEDQuLv81
GZXfOjYoVaJBBk3j/vXyFtr3qEmuxuk4aK6kjrPtmjH99WFP4GXmLGt7XAhtYdI2Y0/IzV3RrOdW
uwyr/wVVfEejIO41C716z5Iiu6UM4PzbBlrSqBh+N5CtmDNbM4asgpVcZOUohCEvlD/WqxVE1xlT
RQqUvJH6TkuHoo1gF0wyihGWSH29KFPz7+DRZYCLqjJq4OwU0N/vEpkmxiQhYF38NpdFZbGV4mS2
r818fYqkda3IGehtnPpqS2n0lVsC2R/8z1pfpJug+bUR9gZJZx+w0LpNpclOtGS020gJrZPT4UVu
aJ5KhnXRI5ZDc5qGFoE/5WR/xjbD+I0Gep9ZC5Vu6qxiGm2LEjBILXqpCuze19DnoVLTupVfaWVX
+m6gtCV5uCAwJly/xvuYmEfR8flH/6Mm2KppUSjcxSVNB2OgsKXgy6zKoeqoW/eZughX78Jy7NSM
RVVl8kVjKtfITuWz59zE+ZgrHfPTe/R5LCQ+6YwOHFJUXy8/aWyQzTRnuM99dSuJqhVZV90KzZtb
f1eQsI8vRH2kWRLMJSbCh+G9Sn+Ah0S0t/xyMuXXhf2m5oIe99jWbqY1WBb0VLxN301B9PKnu9AE
1qdBRlFd8C29qqYF00RJo7Tf0KGuo4SD3gIW4F3BxUpnf7/NzbxV5jJezLAS1deFyzi66vcq3VdY
zuJkfiyeyBmVZUn/Q3hk7LtY6tvFyF2wZJIzet7DEZD4i1E/6Qyq++eqhXCWLdC/qJKd1kb52FeS
2siI9aS6+7rL9058PLFIcePp0zbD3keOqAHEDRvDP+ok7XdjEwAuHhvprRwV+I9dm25OD/zBshAu
2+vhlO4iyWTFaL7OqC9jkJuBzv7cIRdqOuan5KglTBxWfFT211Epawl/Rvh5L50G/hI/RVeVNwvW
ZEVEdbY7B+dBQH120ljTboXDXxIajJjJN+2ltFVdz8/ciQohoPzvt4zsiZ6gf4CI5gBuTWEZUVsx
K0ylxVmXcBvrMziVO5UDd33nLN6x76c4NYOT34h2zGP/L05bjCXdILg1hdGmI9wBy18fXCzqkx/S
p1ay8iIqqV33+jmujV4D0Jj5NrarwcHr6ePg0wcMWgzOHwyA0hVhZF5xMACVr4jfyPogxsvLNo09
IOLtBVBvjTgu71TSrrorFqCpwUXTiDR/Xg4wDa4u2pf5fPBUN4/RdpijbIdIEHn/XaNifd6QDpuq
XsvaGHDLoeo4zwWhoTya36K+WoZCzwqhMeZwcDe9eeqi+9jd87vh/22qvcaqcVG3uoSLSdOw71BC
02bvZV5X4IAHR5xmE7SzKBfE98+y5/G5pZCzZLOlNGTRhU1xwk2tTlo0HLaQu6Xzlxh/bFKdcGEX
xmOumZSJ/UdJpxvJms9lMAsdmtyhqea51Vp091viNyBXpwN/e/COqU54wkVjXZGyUXYVNj3l48um
dT3Ooybv+K4BlFx+E+fLI92PHEYpLH0M9Wli26o5Q+5WD9ddDSKPybns+bXJQBhRRgb39i02PV8l
qnSsJrIQZEm7FkcVCOQS6MmXdJt33tgRkxK8ftOUXFY6gkWGosFwjDQKwaZCdkiyIx7L94i8AK9w
7R+6kT802Cx9PWj/2WOY1P4/in1vhYmmF2bZ2XgGL4N+vsg8ozEc+4PHyvtrA1YbS5p9zIJiuF3d
TPwWfam1nGDL9Oq/DwinJpheGH0Cywz/whdsz28ih54GMuHjvNHsZaa42ULsaeluJNlz/A6pPz2A
9EdBt04o1179RC7Mwa+U5YJNcwVNB/1WKgbGZAmWM1TmUG7CqyyOYFjwJkACxcPPoG3STGbjbPRk
MNDVac2y0CBroPNwOtIplSSqhRXhSEj5BG5o2tkDYWmyPM5aOrnMA5CLEXOZMO0zHl93mAjq3Qq/
2Yi/i0CVTn8ZNl3uQxl4IhH900TdTAadmmqWaNx41bMH1A694dMKhRudWdHdS9ct6jWLlOftmf1O
rj8/MeTToBEXxbsSkp2MM3m3Mh3KLx/xTOEDUZE5AyNY+6rBuYgrJCYqa8UuFcGnnFB4u70CexDA
RqhpdCaZfKoBlnVQYbqw2KTz2Re/z0bCVUOHiiMvoLMRz2Ve8le/DaVFbqpSbqztvCtrJ23ZIOnu
V3bCeWIUGEUUQRzZQNIBmDfVCkWm71lR1XHsbPffmgtAi/LpdQDCeidhyG47FTLLJNetIC6tezsM
osSxhph5Jr7gdjheTqsCIxXjfY9zfxMOI4SX12g55g+slae6QYYTn+WtnFeDbRtSjVp9r9pBuGAd
mPy6d6TCdmMUvfs180M/QPWkMWioZ4x8G3dS2Lm1E2DUWLCBUm3MP+O6c6eilxbhAGUcpw1ZUdia
iHeqNnGcyYZ3yVw3kjdgoKCs1Zdx1OaAIalQJwekt3LiIoVPXv94heEtiXQkoBde5VYgbksqCNjt
nwDBvKiqnoO+y+mcepwVz3wuZ4hrjRTzoFOmEuV7jCs5YKoxfjZ0z1kyB8kird02KyPYfCILT3NN
3bW3JXbYnai4cr/PVfqwPajgXjYzbr4UaxItdBmV2Dyu5RIeQwV+lEWP5oni+r9+anpE0IahQMYy
WnxCm7SceaBplsPqAO5lTJje8LeMLc07klrYQYr1yEtKTKma8PYZ6ms2jti/4M7BWAdMgTudcnot
jIkPtgLACcNzzJFIglBkSpS+i09GEhQ56rlQGN6s9xlMdECXIU2CotgV2OLpqUuVkn1oOejXuLfA
YC4MEg7DHwucMYKkv34+zkRoohzbKFzwPP2KCs3Jt5mEe2S1hKrMDfQd0KtoiWWHlipO7sAmgw5N
zbT9UDN9e2bLuu/YTmasczjSY3Cnfvyxb6WZ7rMyQy2akP+A5ex4toFtrVe1UvGng/ngJgvyjb7l
r0EM1K8BHJkzIDYP+wrQv7PsR9noIvI5IcJfKSk2WwzJXy79PRUjCcKiw8IlGEYQkpXb2qpEm3Nk
YnuZZ350s+X76+dkXSMk1Ab0520y/t0MQuydJaBffglsAH2rUuKJFfwYp2zpbm21YwTFqZvJHY8a
bxAKni5ELSR6zpy32ktwRCio7D6UkHYAdRvc/3hWsM62AxH7jRTAVtyJioZmr3q8dELNQcFJCCVH
5BJrQVshqnMDsKzgkDXTMP3p6tnw74POx7+qsYG/5qI76j0knZkp0HwaYzCK64xVnTD24vE8AZIs
/irKiOe5wf9ZJFMZF1uKtu+vE+y9nLXGr9XUNd3xsdG4iLJBIVgDxOSvxippd4gIdv0eezT6sqE+
/ELa7IlLU4i8RGgHBlG3ludvg6/eI0sGZ2M4VlTPw4kfeeoy6ByjhqrM8DOEUalu4uE8M5iMpo3R
XdBqVZZc5Uf/LMYT0q8rsVNEw2gWpO0WPIEPAtAFiF1Q/augEB0EWwrZBv42eCpBi5nScCNC4Ub2
o+AVgfVkXDUMNm4nOqdSGEjIZmr4MO+DJ8RKephB81YLMqmdqhgH/5c1ngKKDCuNc35G7KpUKJyw
BOasQ1zGtFfjOiZWo97klejSO/1433FWKih1Zj+wiyLW+yumip2mx36KGuN31nq4CBpJPfnmTveh
f9dlcNHFPF86kpLxPRsBegIQRdA3QwGOLKptJsH1zZIkOYAT3pi1xi1Zs1XxmemMnm9FITSaWUDL
OxJ1rGGY9E+tJo9PCSNms9WJikJBpdtFtbfk9UZIqoLRYTDkGkFDN7VeSn6KwZ02EmLin5j/MxzG
OPe8GPMMDgI06m5tNrRnFKcVm4JVXU93ZY/teMMb2+T/iic/SPErWPxe1e/KFgcaVkkmzT58+BPt
1Ny/ePdewXP5jwYRy96eRk+LlGzFkY7vyBUqiMMDwGC+5tfroadtmK36Pdt6Rx4Oek8sV02BoncN
HvJorHaqG2AXd4EgORUo7zjf5DMzyZN9zCMdpFp2WXAyfEErU7VQ+wnPB6QTjNh8qyYRduZ3ZvA3
be6T62ZOPwXJXJCDSPIInSbul+PGnzWKFugWbl4tIli/JWA3V+c9cTTjL/CQ5rkg39sRRclZm136
Y/1yaLozhpFxHQB0FNccQ7bv4HP+3xzMfif8EuKdWdQrYd4GuRaGKQm7azwwfy2MAQKiji8BaXwM
trsT+DOnsZ1mHmirMS8T1Vzu2roIEl2qHaSG1ImqfHykdJcKLiygZylrgFIVDf9gfzqUwEAudqma
2c6QRIPGLUzD/tYkrZ/CIQvz8ihW2G075zNHQrXFNww3HOhwPNq70Cu7K8hOgFexSaWpeDQetggv
4IgAGpN5+HGoYHsqBSIy2J2fdr7VgyiK4TWUYaf/FEFSALuJ2nimxaL5oln6KTMHp9PJtOlyRasD
F0v/8gR4pOYF2ckh+5g700AJKsdY4L87WCb/iXaooFG6sCxEqZ6wT7hqN8mf0vcXc21ZM3oN5jQe
CgGlrgrcJt0YjFxJ1TezEFArBJL8FT6o2yzFd5tFzukQSy6UyUr8n3Wkr1J8tHYIaGeBDP3naD1t
DtSg2WJ0bIbpVsl9HOUu4C2N8/kfkRqf+VHZtz5mWBKyTOu5Qnq7PDYcGTuf/hgmE0oHhJQP3C6U
wwk37npEY3RZeZWncijZetAzRAHUrJXRRt7fK50C1t0agQVplaGqLvPv4LG8J8lhlYLZFCdmE6ed
FBhdIfhS11wEEdjZJjw1cf6/lW+gwGi9iEzfxb2zzFWijsd3hsAgZcYUfsyiWrWhOPLvQfBWEeFJ
hZt4TeHh2xv3YqGk20a1v0iLjwubIT1B2sWCDKq17HQxUXF0rLytcnxzOGee4lx/W2lcRrXVnrBS
rECl6VYtqi2fJf/AfRSC1C3zu2nNME8GPa6kL+s9ync99WXW+41fn7BEWARkIuOO8JK6EyQz/Kzf
gUEOIqrUYxw+fwWjZdwvm8hd7P8aOb8GbgLD4kJJNMKerM4n4svkk7/mUPc+gAVR0scqQ5dEMdgt
E+xpTQZwGS/5K0X5+8ZIPznzHKEF2JvrMutTL32O+Qxy48JDNSaaIjg+KbM0dozA38Y+g8IT7K96
8P89Hw5xJaMzXUpQtGFltQodvjJdxSrQKFZUQFXgFCClFnMLdGI/L6JzC1ikziX0/XfrSjEcHKD1
j6djYaMFzdXLpPour+H1XySYR7CGKbw9xe107bn0V2/KfNxUFcIpD/gUXgVtvrdykUGGZ2cGFNIQ
WtX8l9ZqwQ/+dILWz2UYPiRMsi9mguaddBgYAMWM9hSR7l3k/BQBeOA4lkAK29JbT/ChvJHrpn70
W1lqm7v0o/WCBNu0c6KoyB0EEPSBiX/Hft+Iv1x6el7fIe506IPDthElSxEelNpVpwnRWXncZhYW
ATpCnoBLr1k49nPvxnEp8hLA8/9FMIKUB5FDVkMZbCH5hvDPTsInvK+AFEqNJnHHkOIxXv5XGwNO
arEMLIbEDZZZT/lwQCIq6T2ZO2K+SWN2CLqEjdJCqOSBoww1PAPPoa46tqO0G72NEyFP6I9U/dFN
bdjCJGtUBJxEdcwyeMR0x+GnP/154I+iSvvH9o1M/tkdqqt7QeiaaDtibNIPq56rnBzvAowyUQHy
wfP22lNNSVQeTTHv83oPul6mq2hBWErWQ2g9eQzu2l2QYu/++h1l3bZczOBGwbd6IvzSxGrmWfqw
j1TOQiqSg2PqH0mL6/MRf7LRLsZoXRmk+9dISy9QpLSNkS4OECop4hq6/4qe0/RSbHrBDhkIp2Pb
ILn8I+aQqnGhGkk19ReEKqASRf7GGIbzTyFz6x3XrL0cGID/WwCBNlXlw9SBUsFr3aG63JNOCrLy
GEIe853YuFEeYlMjAFM1gX8ynm6SOhGHuDiephuN005wkjx95P9Ge6sA1+OqM48QfgUGWxhCVB5q
Ru7lMLKT1jURMV00ZrxiCV3+SNJWhzy0oHMG06FJVsHBhNX6NT8K/gul2EJzZIhzFM3XIbkrlosS
A/Mb4YZENLlDr3hVFLfOnTMNLyYPv4+psuV/lubdydwxPnFazfvYrA6E7UjJraUKw405uHRq3fJh
EvSvQOuIU6481ENEXdcSrgVrbNgA039Z6Zd8+6V1p6/OKNPkRjEH218/XjW1UanpvlZQ+XKXwMRn
QnSbIFsYYbICPzQAS0gPEVuU7t6xDZaaWbzGV+fNQKkCq5NlBIUpEFQkZZEwbSwNDC7maYehaYGl
ZKQkIGDb5GGpIpVr8e/HfH4YIEnezLodbY/LNvcK9ST4WYokrTtQzjbIUabgVNx6x4CNFpr2okiY
UrEn9ctzh9Ffz52RjYjXwGdaduNra5Hlm61gUzeRJwpHcqy199Ac4hYj3X8yPrC9JHscW8HAqvGL
QfaaaxqSYV0zC6fcg+K8ve+al9eLBVBabDGzH8FAw1W3PHHRYmD1xe0B2TO5cc2rewSFkl3FEYw9
vTMqwpl2FpKKc+MzjjO/5cBmri6Ml8jowmPQ1ccjBxomT5Z4JG9n23nnjPG3i3UxI591dE91EiWu
PU64J/52In0Hc/u/YU8rgE2K/wIHqP1hYOApdXCm1XqP0S021ELizE1Yyv48AbAiFZ/6eT2k4i+Q
AaU3OMr7Wx1fk7KkZorWDIRXba6PyUvJdtaupGu4bn3u3VuCeWJ3eC9kL3I6q1n/ox5ABB6YBRle
Peah9nhz36roq7hwdehV0XD+kobu2Ji/oU0GrvFJrTtW19CU1vVig6F43PtfCc7VfbHkxVFWhxa/
zs6WSjgdnLVAEJhtexWY4Ku2wPtGvXqnr61XQS9HM86unu/we/16v8vTsSh/FHxhqx4Q7gw4KrfF
vDKRZqmgXhieK3yn4thjQybDWiVRFWaJasyy68Pcl9BVA5svFrebYGtG9qufJgIW7xYG+IzLyXWr
9Qlz4xGJ+SnCVfMeR1fjyNttFaJSVBu/s+ZVQi02TUbCFuZZniTVrBHg5HdiUTKBsQBYIRkDRYD+
bWa/7zDqNqkdBdN+epAJyR2MZNC4hkRBUQvPFP/j/8+W1jdrY9pYshhdCLe2+ItlcMwTokzmaXzx
7pho8t9ngwpBjMsalJTDGwEeAldIeD53CVMfCce4AFNfDCMMK8yCd8WtUFMtS9w9psIza3/dIyRN
JPUUSHPn4amqnbhIrBq3bIdeJfhyAuzDetnHO1e8Fb4GM2nJ977FhMIR21QAEx7XFSrgGUMYik1K
UK3evpYqrXU2cupVmV5hw0OEmNvo0XjeU9Bw/9H6ouKZ7Ay5bSeP9RfuNQROJsvP7VvBRSfeh8c9
A4zqk6fPbkEFGn41XFbVOFSJNcloN9mnIdfr9iYQjNuQtCVAm7j1Ad+xPMuIm0T71aoqFNEWojYb
C9YVqiaej9HHU0e/8QQ3Z2h6+xt49n6A8XSNOxztgznk5TTIyJBla0JtSOIz5wibSZ/0PLTH2iQ0
Ugkze+HzNKsFw8HDI+13EeB24HEc09+b0g+owawwa04kHudwoeyqPt/uSPF2eDI9nnT/zVqldEsG
a/x7XpV9uAp4sPy3duo6AmSdAuMsf9zI7pR/yfQ/uzSR7GMmTe6RBQjA7B/wHR7kzPcILxicQ57B
XtgTUbZruh6H7zPYOb2ZCT5+z89NPCf0yXycW/g4EiNh3zI99rkP6D9ljgnnw88Wpozc9VNxqEjW
VzD3CE7l1PSqAos3rlZzc61iCqh9G0AzenflzbNtkyn95U1RiaUmU9khC38PKYpSsnovNsEFOH26
03JVdFmM4Jn8bB6dr2L0FsuCPrX44O+YraJlEmwn2Tq5nMu29bg3c3SW+WsNzTKOq46ytCAuyEyr
kds9qF4893j38LaE6phwXsh2IUzZ5hPKY4IcfuimqAE9SRotQP1RjNpurEbgCLlet/QcYksQaOAj
9oOQ4/t/NKe82blK2ArXdtt4b8UXfhhGJZyxOM84N04oUti9VV4YQBpG8oqtlM6AVOIqTklaqNdm
20I71ZanzlebchAUuQKrevmcwOHHkxqsu++Swo+iISu+Zx4Yj7x06XyBTAADZJ8jqV9vgTkZ9bC/
U3jsX7JTm6dgmHrUR6UC2j2iCjZfIFOKmkWfXQvF43WS7C+gE7sFesXPA550SvrspzZ5swvEHuGD
0erjHj/hfpud9hQsXjcNeFRYAv+PAmpaZTxkJLXlVNf/f+GF2G32LusZLN3T1vZ01h8iBzi8LZsF
eViCk91Kma3XNvZYT5kXSYXh8qttNjyWyAemrQXGW43yNPPUi/1U9eDSMpXE5f+RXCRwOXKfJfpN
DV9MwIjgzn/NYeU4De2AVjL1CKDLY1XA4QtFUYkLI9tX58Sr+GNtAwzpiL7Up89sVZ4cFXIplPBM
CX6EGaDh5KvwGiEYBnNbTIYHaMZBHVBOze0lX2GOFNqDKS5/Nr0QlGPDztPJcMXQfhSFZ0L2yEaT
LiIzSEgYI9VKVlDBKK/TEyK+wBFf5KS25sIaxBvaHPhSjoCneAzDXPhK7w4k2v78LYRRqDUfX57M
YVZlhKxhdg52v5Uew8MPmdYs8+TGjRI2NLaTw+80O6p1UVvB71A2zcgKC08JxyfVaQxM08ge0Bk7
AedgrpK3OnrrfM3KX2iM7S0vuC4THMK0kkjFEBODEHDCzOWBTvwD917o4r6ALH6ZrKbuz3PCCu3A
RFIpvRvey4qwIhdf1hmcBOcz1hzHYQPyPYMsXUImPAqLKBJEtI9MLkNT9ge5oGbaOcjjtj9CKOhg
AJzOBYGmHXpX8L783PMJN+8VkEM00VvFf87LuMiFzUHaTsOSiWBtyGONep60biv7t4Mq71PsNiUa
eAFZu0wirrBhKoTGPRilcuv9f2bO+SFtclAO1MFksolAbXmVMz1f83QZmHfyzab8oJ2y0KjQmfm6
2QQTWdQToar/to25W3mz5sViV1eK/dDTPGoQX73m1g4uF3DasjYfbLibD/WJexl7rANF7A4hZsV8
WbrqF2OGxm7fyoRj52PuNFUc/Sf0FOvqBwJdcYw53JNuRzacVZAZft8qeuNwUfeDDwg/8QXczbvQ
gXz332RwlcQ91tVdoAKMfvyyhfFeEjkY4Gng1sHVuM7lsmnHvLsWja3dZLJ6PIq2M/HthXvNAtNH
0/bF3Bs7h0jWtGpkaosKJqlk4mo82/2wicC7fiKaa6NtkwxbIw7IfQtZSlWlmbPjNSP6La6q0eDm
5euhYcuNwOHVBWqHlf3wgy8Z8UmPeT1Cn3siXYp+Ie6hHyoIkujZJAmz2y1Fc4AJBW+U678Mpy/F
qqcIOJmKw1vk868NdNf3q2F9D2u6ujLATlholNz8LC8kHj+iZ/Uwj4EF8exJRARcxCmzgOCLquVS
RkVsthCgO1YnWv8C4aLGgB7IQm5w3vhWVC0cFt11XvtYSSdFqbmpH3xvUNtNzHM0b1Udrpz3xtuj
5ayFsZPAzNKRBxIFZyOoiDLd3CMpJhcX/LMUeAO+PFp0VIJVgTtXD4aiYvS57z0Nl8bKbhZhJ55A
Tl0YZzT6FOTMwq6h3K4uAAwDm+zb+RWnXGBAimxxVtB2jd6SZOxpVXhuv4Lxetki1acNEKDbQLgR
BspkiLKdlItZluLyQIq6uaexwUYs76kWpqZxV0n8nxW5texEkt4QWsJNsD9SPzmcZepQMhlHjxxd
pwE9VtuALGTE2vf2+XGq3qghNdPiXzNQw6bnhBjEaBd6txczTGwrcnPTPXtzGpbcpvD/7YXVP90Z
EQi7DJdoDxc3ABs2XpciyGqwaNayKSYM6RtXm02/KBado5K/Mpj9Ps5TkIDj/EFQyY8KBNPZKCJa
1aOHBiJrWBT7WjO/U2jBBVsWaZRkudJU6WU+J1vQtCVBcDouQk0GmwAwAEit3QKdApdRxIF4tXh4
9WmpRVWHtdnxG7bo6goNqyYbpn8frNGuulfzi5aNbcHHUCPLDcmwaJGhuZ22BleHM+hQbjmMW/n1
41bq0LtZ/lWvvWdtwhgdoY1WAqCU+nyCKvoQCv90vAZBUav5B2rYEylLe8tMInBS5KYF+C1Y4L/d
P0vLXhu6r3+FacCeFregnPJBbUx/q/rvqaeR4+olTI7vdOYkZ7pcTulPq3R20pwAqIsFi7uAtM8F
wwMgCLIcASZzRQE3tb7pWG6sUQqdzFJB99V/WyqChyP7Bxla1RAGOALVpe/2XjdwLAcQFOijfzoB
j3oBcIH4Ruh0CUbE+TRfHRm2vj6H7FIzFJRJnsYziyRaR8W0UX/yiUm4WyrjMqsu+AA4LyPS8rCx
fiq0rv3ran+bGrC9AsOr2g52GcVOpjEFhpv8W3n6Kvu4VEYod3xFtnXw8UTjZowiCEpv6tXkQi1o
pWzpQCU9VtPHmSDHKCnk7BJWp1oSKPyscVH3NnG+uQCyb0uSh9aGk5H6H7Oohzw140KERK/SpYnY
6FciMONjo5PvwB+q8XhotejNfQpARn+dUMsHp5Kmbbcmr8CsE20SQ3W7q7l5lKyfFYYQtky2+B+H
MTOq5Ar86fMi/PnuREWKXyK98U1wz4r3WvpjzwZJ2B2em9NmcqkKxlDNH8UOrw==
`protect end_protected
