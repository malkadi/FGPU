../../../../../RTL/CU_mem_cntrl.vhd