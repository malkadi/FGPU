`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
gD7l84kB+WAh1ATog3H36h0/cMgn9QL5jGe9p9PjvP7N+FJAVvGVlrxcgBw6dZaWDNZqNANQuRFv
ZSE8fsSCFg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
YQUcxim/tlzHeVlJ7otHN7u41KO3Yg5DFb1yF4GCsbXGLtUvWNlkFjY+UPIlgYImR4Zo4dTHJQ+j
3BaUNSUOqAVzT9CfyUelv2YD2ZTfAtzIe1Mboyb3+StKnuzxnZmIhVPiZlowdW5lQ1r7BjDPOsge
ztxOfUTbvYcTUE1ABIE=

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
eu4MFD/NMz3pssr62VCh1XDd9mthYydX9VaOq3lWUwHi5/7e5dl2SAWHtYwTnBgGPY+jCcMycJhy
WSlkhQxVj5BsMm2aAItwXFvH2mSbjlPggtI0/+DNGQ4x8LQSFLTDYnnQbBrHlJymsS+/asMkXACD
SJ2tF8LF5tMhAlMPZZ0=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
rNAzbNlIFUMjdhvgzZ2FokzvR4AuFtV+1AHGDKa9QgeBsZ1e0Fom48uKbJ9iakvqUoUcKKAvRzeY
OBkbx9P7Imx0gvIgzFsgiVw23cBYWOhbhSqVb7mef9aKx8yeF8T48n7gKldUkwBHIPeqaayRI9/Q
HCZO+k2+HCjRZE6L/Gzd+IOdEVUFOg3NtWFPk2JFkfZkxs8X7Vg/xxtvH7uvp+/EbVyiMbnwDT/p
NSqOyA+rJwBJYD3xRIPTFDI83XJLCF+1i4E8hyu7Y0F9MtjKugqEHwAG+JK3jde00nzNNaeLVUQ1
OfFMZJpkk0Cg66d2cvJY/G11oPkmvTq/JZ4+5g==

`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
apuTRT8aJu0TR7Ciy6ONiGK4AT7TUEiokS4gFf1g+kDg6PdKk9VRun4HKszIadRtahjPQo0of9uS
yvu3GS4EQo+Y+T116wnAIXnZSa8EQaEsDkziOI+rCvXv8IgaPYN8Cq0aRlASFL7IHOWNI49V0c0A
FIG/+5U7ZyNQFCVwuE4gCgK/pA6apm5kY4FGJft/EdZ5YAbR/nCTzK4P53+XsKHrtGfw+/MthFWz
tI0OtloKqc7laKZWKOVFqWq8Qmq7UL6utFODtxEQqzczH+q+Gw4rkUyOosIY+cbB67hX+GlmXXEF
jMwvUcen9t6c+wiH6rmBDcUIiuUHHz6q+jCwJQ==

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
dfDj35aI8y6zqcW/IHFxmCDw2mpyex25qQAUnsL+tIRxivv/85PqpCOrf3b7NWnwUKMrsxtw+JBY
mtlPsVxQKR1gn6VkaHwbEgwxXXxFe71Z+1nWQhfF8Nt55jGvq1joWKMrurSV7Mo+HkvHMSszXj3v
8ElD0S6sN91oml0nObejOhxzHf0ybK+sGag+CFA7aBr4k4rYglf7AzOYrPl3nNoCkyrFDQFa46/w
SXJm/os7zUHbsDI5GGUH3BU+NktHZV6GK3iyhtHTwrMgDtpGk6vKHMKULM1Gjv9g1/jp9Ao4cUhr
bCVOXM1v2e8A3564rmh3if78zTzCKamPRAB5Ig==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 962560)
`protect data_block
KwL5t2oQy0aWVwqsJj4aeSEHXCHCxaOJbX2Nlria18v+Fx4J5prLcyZ/NTVPBRMWjm5nwRxaQLXQ
EWZrT/j3YoJKTPrxwqdSHHHxB73e6B6F5JRoSEhoC0FY+Zdwavi/MerTcS2UyZfouWMjy+wdQdAU
z4cTNW0GySoV0dKvkY5t/e8rBiNEmjfxCnjosV2X3a4FmAiPBPJaLFVMPn2vHR9UvHrLQ3yFNizS
MTKxCgBzAHtIZaewd+F9/xPl3vAEY7HxEAZgF2oZS5U1I+01LCUVWHI9eD08MToIjDRIjKU8G4qp
elFF9gtlET/K0nLBP2nAkouMk8r0RQLnc1xLoKCheXXoIgvvvY/2s5GhnfE6ym8CH2N77JaJ4Vej
6Jhmgv9Bom7xd2/McOgBL7ul3Eykg5/4R/NWyDgXhsv8cjFZISczc7htB+h6uwoFTOK3neVF3+Y+
k5F9jcV55STabuyyHse6CJQPrbsrkrzzYB1tiY89HvYhU5jjJP9BrcChvqewLde8yYqWbDI62IyO
liMz4dETZP1rrG2+xqj3eBmtOpG1PVK6Yj+GJMha+rb3/WkmMsWtAisZPJt9v8uIo1KhsoWHRLsU
VZTBo3mYdKZxj3oQSDRFX3haPnT6s1CVW5sW+xg4n7eg1XzBXORyZq27lCDJM8t0KjPxHIN4V4yt
4mmekNEkUf5eNSVxqdRuz2YKS+ctGXAbuAimXLFSjQ3CLo2iwP/zlvINZgxCEams6toD4X3Omv7T
HKpo5aOepiqRxhbtLOhhDdGWaF6BQXHjalqp1O7I4zrGYmxFXuaXFwuLHVMwV3cKck/OZ6zA7Z23
JYNshpzCMhI0NANUM01/fl2nsZXN48wJq2ov36qv/sA8ksZlYBCxU0IZ3PO67OM+Ecvq7cMQt6NT
mJZPI6LD82b6+Cf5aIOlhgqKcDCfEmXkuYiTKJD/NaZtAnSYdHyNW5nj5mngP0KrptLkMXEKwPYm
E51MMkJkgOI69A4we4vCQ1IQNCTgif7A3aprNLzKNQHZ42CuxdPk/5HpOY1l85tX4QPfksCSuWCB
8J+X7O3NYucCvd1uGk6fYpjFIJm4vakgd20xKyqILSTxcHugiJ0bji+cXDSJnzN6SbbkQUxydei9
CeYYCzqKyg6soSwgHJ7AS5cYIc0W9mTrIyoXLnhEtmwjNGLIzhAusIayVbZebuhq4CRrOnM/ES8D
UuiUYEMXpupw5UsCycaVoIfX893air53z8k+86UZjGLAsCtRxTPSA78c+FXtF47R1sQ/bXiDmxKT
3SrloX5tnN4bfZXkAWgdL/336tMW5n+6gbmrbPCCcaVjIXJoIL+YNFEs9RbdXLM2PNzu0Inralaa
4ZMzVnE4wK0jh/chMeZNvOFq32sQFs/+Q4QuUdI1d2K5m/MNVn2amtTsJDO/n3pjh0ILt+LVC0jK
A/UTZg+VrIfj99R/YyO5azqY0lVQvjOBQcpmJQOxqCGvN7cCHO9F2wwO6U/kru9Yh6e6SX97PV7H
8isQAJsjTF3NbY9h5Nbn7nFxfjcPWFJvKjACqVdK1MAe1vZAumzfoxNuyQr6rxG5Xyusgx07KijK
1j32hxE2ZTzPR25EVW+n3rUzkO0EOiCjhy8myFTMn6ZS7Gu/hCm5zFgn1HiyCDSI69bMhK9+r3Qk
i1yydyjbU6o3C68ieH+N/UH/QKJFu15DTnDJM9FfcegYpcGc/0Ax0VV69HP9Mt8BONVEQjw/okwG
5mHDdEEwvgURYIHojogOjCBLbmo99SZD6EbHo1y4b1zKYK2JtJHqLRHGRX76OpKk57/Zo2x7PCf5
GPA+sFkdAtP4PRt+CsV+0G6qWMqWWbp3P3P+aU93pU9odEhOksEWU/Ez00q1m415sQ1ejiOZmDUp
5NXGGhYZ0QdGfWjIQhowtALrEAyPe/ry7bWL0VZpK/T05oJunDDfOYiHwMfwCfOAdKUEiHDrAf2y
I/qdCVSR8TfcRJHbrUyFnLxmlxbDUIYh83MYzGv51y59RDprgAN4xCSTRjU2JGEjVb2gGoWnEbyf
Vpqm1q6r59vZ4GoE04A3J218KHkvPvGutQg65nKR08exoEg4rsOzKK5QKe8CRFh6dWt+zRE7+CgC
DB/kbbNnWoSvJ58fMUwujutDrLlBHOQ9D/orDe89mNR76+8mk17f70oI6UImmcb0/vzCrA1cz9Ez
J80HatMxizrQdaRAgPIpcIJ4FuLctDONWUUyBnaZhCXFrvoUdc9yXq8sstFb5s5etBz3rCHkYcVa
O4Dn3I9cNrt1HWdEMyt6cSytbwkgjEX6jE63QRGfgJDDpggOvy/lt1NoMK6JG5VE4tlptbxFm0mw
jgWNyKGBnu4DiEn4abQfo6ucPCwgok8HSAAFJlGSJ1ZXxw++bK64dVg9PTMFI0tUZqmK2IvGxdSM
9I0TqNM18oPgXYUavDdorVubiDSLe7vI1FC2RrhJ7W904PXPtmCHVOcxvT3rcIRULzKKOQUMgq4A
N3RKFEhhr6Nx4CDSDsRrAP7dwRSexz3LZBSvCZWD6M1didHcuDxgEOgyncGPJDGYGE9lCnpfEv3s
QCz112/RNf2eJi/iE9Yrsea8uuzjL2bX++Q139voLVnMn+0s7QvR8Siu+OBalmiepbhtTdPLvSJS
VBxJme9NpUpa/V6kGCi6kFwqFmGvtLOm7wm5hZj1ZBuidRAJ1+y6JPc16yBEtTeDJ7vSIiz4+kai
/kc3CLvqMoYZZvSS1Mqhl//8v6cwGkmA6Kb24MyomQSocSX+BXC3E9/ax3N4h83eGjpXWnaTQpgP
KjFGPm/1PgnvOZhbS+hscsqr2gukGmLaI+75SwdhJKoZUJLQvaCd9SOXWoAP/lDCTegGu/ZpwjOL
rAwPuJN8i79UGDCQI+AKoIatvH1FzGQSN+5SuKfWu8qOC6zgc5xaGUd6+VUbW3Z3uKqUcZARHOq8
tWSsk3OC9D/iyN2EXljGP45B0vDZHJ/eYrWiAeSSLtGl7d0v8hYgQWhDHAM1MrZhXSfWf5oVTGJW
3xEbrOVB9nn8458lCzQtKVEaRZh5xtEP/X8VUa3AhrcDKr+1CF4rFgvj+wVy8GvyK2ze1UBLg59V
ebqjnsbF8NibaLza5f5NsS5eF6TdZPY9tfiwuhsCmjA7cifTQveGoT/NNvzhtmUzVzqbcdgviRDx
hVSI90z3PlN+IVdPU9TrU+d5SWlmOc/1JTfdZpldvp18EdD1ZBwHdnwEra8HY+Pnhkd3t4dF/jYL
3Wwlr96VAKe79Lm2WZd3C3FWK0mw8vs4E6BhavyOfr5r9UdF42l99q0YunxD8crm28c5m7jdjkRG
28QwJkU2DnCkKdxjH/W2kojEy58Wny+WdSyHnKksl/MmNFI7oi7KfC5SSiwajuSq4TiurAl1VuMp
itPvv3rGpoCNCGQB/hByaHYOaInMUvZhgZ2zsakpTbr1MOcJ/DCHX9kJLK8xEzEfcl3hiDmICBhC
P5pgGnWEYvbj1gjCGGv2qb2m1Kc6m5d6ede0ly3Q/aSvh9ptrGFjsz8ujUtFrlBNfQy4Zp1azeZP
2rIwzxQoDfjGQBpAAfYAvQew1OH557h2GtSHXChbsU0IHNNJbG4nG37EqPU6hOeFtyOTL61yPEgq
O4ZSulebXIAFlSljdNNCRpRH1rKmeqUnGQEnLwzPqfzplfkQVDD5Ghd1IgvszAqB56lvX+1KzNWK
0ymuPYL74nnEjqrQMrFkgewT34vkryo5I4Q97a/0iiYTjjYO8t0xUpyYng4hKxaNd+Nr5MNKCPuo
xoRJlKEnaZENgcxEMkpKENdzPNdZo9pkYvghu8p6EvP31nO/NaNiyqweuJvJsYj9g0bzAE8WXzuG
C15OJhK/b0NTi1euyp+mtp+alJGeYUlhImk7eLgNkz1TH2ekEgxTCVcca5wgl4OBQh4uKxFX+Ys8
xUbGks82SZXtMahzK2mDnJJMgl7xrvDtcmgaRY3vLdFxm/XVqdSRzGqjoxY3xadxNKRQxcGAMyZ3
skSkSit3NxLLOcUVID7CfFkJ0KfcFa6y0k79vezwldFmzloxz3e5MDlzdDWpVVEMAaCBomxbOS/X
vJGuBBnSzBzhjbaYgaSQQr2S6or9uVB24oVp2XrNLczL6wiuFoI+LD4T71Z0JGMBCWqOr3L3zNi1
RXYgQhOooTux340lw4ymPkJ96LF+0MdDkqqvW2U17R3tvT31ZFCxNYEnFskYSaaYoNY0wgTJ4YxD
K9hPSdLIVgkeTAyM2YyNaAeV0AxqAdpw2FTlO03ss77IRe5PX+1UFgqK7NJJ2lSqNy+ttQUbEYSm
Qzq7vlURhSa7GTm0jodqA0OvALO2bdQZ/LQ8cFGqHQv6ngGx7qY5VYtpDasXqtbyO7o3NXP1jTTW
5eQrDN5YPhQEx27+5JfKGq82bC63psg88KprTVUSp5Xf9SCfLTg8wMXjO1a2O3ny4Q/km8QUa7bT
4NRjttgRzK7lbxwKr7si5deOZB6mRAh8rKFQPqm+NhR8iJnBDTKL4iL5EOGE/1+RTyedPDF/VALc
n31etqCVQsoAcJhFXAzI7x0FWeDeV5csCPD5LgBnIzi4yOGmVWPwlN5QVK9CgRGecEpqtOT4Wh8I
PO9aWhXolxgfrhtSiRgJDo+1UyEZGYbYINOdWhyg5NhCMvz7qO7M0Qdb0vZ1CZdNdnRRk/WniLWo
PH3DR0fuvviZcF3ro+tQPKL9Y/hanNKqyvbqEgbf2wa4AoSPrmjDa9kXLb1E2k0QJLYHxYrKY80l
AhJyPW0yGBhyzW2dEVOK+eAYMOvlXLH/fFpSEoezzvfQDYEmmH5eyCGA3Kwqno6MxPgCwIS2Bvxv
fvpD93Iqdl+wjAlFsJfMUhiHrg5/sm+WLlmkVhn72y3N8Qct2uQj3upPA4oxtFaHUArqMFWNJbf5
hGqoaIcL6dyr2TGgma0GxCxJ3TOB6puyErl4qAgatn1ONr/YCnIUV4Cdu5yH8286iVxfSTvbdLcM
ShRczmUOb3/Pl7EcNcMdgWiyhxePSWKlNb0QOSggWW2gNtaDCpCQBzRVh4WIv96WTQjnfOD/WZHW
CcEpdZFNky5Q7h/KBJ7/0/gUpWXHAwTrjdHGhU/vKmNmoPFHxfarnPiVOe+6gjlKkTtG4Q8bF4B3
nj8HhoI6I5w6RSsD/89vLY592X819HiZS2skWqcxoFZAv6GIUre8NLcMNDHd8Ce2O7UNjMRGOot/
7LE/dBC5VM6c5toPbbFpF5NfmeAQjf+8EM2l2wGGBd57HHAeAg5dFG8XqBeryOYk1yHALvZbLGI7
G3BjeJGoewcXIMmFG3OlidIF+2CkqJuUOAhyqEro1FFlf9lo0daZkJzJ75sW9M1yW2Tit0jpKjPi
+HAVhYZKMllwQ1mAiGj1dqfcIMuXSGTHipnJBUOd95fbwuI3GhSfFXWZ6kFDmmMcxsGjBVsRGd97
Wn4bbqXvQGzOd3k2Y2iiuhtXvjvMiacJysOcwZ6K8CMegjFE5/jQaKLCUrDnSZsYnxQzAaRH5zPD
trC8i26JKVpj3/KmtDWaCeAMQQEywD8+I8YfdIC6XaTKFe5q+3lJcy3X09Rnqtj7FyR+7Eredk2g
8jzKMC/jsiu0lJ5szUnOzVvjWsuSVpbHcZUELHZPlA+hWB2M1lNxgVK1L5Y0bmQLk3IQrwJLnAE/
yRVwaWscqBNRcEndyBmX4iHf/jSz+lUFZeZ0DK8gJQJET4zqF3/bXckWjBaQQh+aFTnCRVhCStUS
P5MYU/Gw90scAeSFa3VsQJC/cUWqBbDCKHdYoo2cjlvYfnpCymzvLAEFhjDQ973XAO6EsMQL/hAv
YqbugJidTc/0UUcuGv1Fv1Q7tg5s3n027556JP+Opg+BuzugFUWF+vOWC5fcpik7pELmcQPQsAuw
rTWyuXrK4itTLTT5e0PyYYbYHAlFPd91DLJQlWZY3znp1uIx2Pph5CdLmNw3KOANbtV4+IeBK5sU
TVm/P1XZcpl9CTCqgcy5kwK2fjnIUst9HBx4SaW281BZv2M3tB75X07nBxfNkNpG8VzY/CLDNJrI
OirjRvs3swwdD05i8RiYPVBW/gBbX/fTkAY4HZH7dYFNMm9s0y69rBmoscntrmWvi7+MUUvTWUCb
jT6cMY8XBpQUrROJsXqyzbz4xzeGvngZsIhbOBtkuBn0X59WBJ6/xVJLolqWL/ozM3GhwKIe6zFs
4AHpK0QhrhwcEjKEm0Uy//Wgdm8LdwTQlAyNLhZl9oqLkwv6ZUN4h+zCDgU/r0DLrYKjYItieCFf
DsS4meu3pmUY4XOK/hdit8BdY8HU7NFxc7D6e/DEzJaAWCa3TRBNbRZm5H1ycOu8lDvijPLmu43l
/C7baP9Q94OYYEadTe9QdanMpmWGGYCosYJpF0Mi1h8x8+3zFl8MATvYIlErLo/nbaFj9lqcOkLm
tIzFw97iZIT8xgrZ6HD1ESprkNrJg0wUTQnttwRlxGAYyFXvBwkCJuEl/TMwArzHtDHe00ILbsje
1wT8Ai7UUF5BEK9PvHtAx8iHvcgiJicQmc8ABflpNUGICWXWtZ+HgDOyaQnA7Qi598XUD5VEkiCV
wSgkMIfuW9zTAa3l+ggPG+u4MvFAb5805iSUYcWREufS2CF7Ztuq+6f92TxXu9NDrdbnxj4XhR3E
s4fUgA7STXuwShWkUgiYCMOXyChEk8Uz7q/B5QtWXhKQmC5FjEHLmgte69TxZ3myFJw4oyED8oeb
d5njyO+QDeKGsG7dT4mDTLb1UpvOjuBJC8+JgqB7n0rIOzUM3Z6wLqZAdRfb9tsdCIkIek/DrwC/
Cn7eHgny7H1uI1OgFTBnggRXkwb0T8GrA1+KO38b9N32JXkpLp6Qi0rxrknQkVFnfeRqehFhwagN
igWPazDNcIzEgHy0e3uO8V9p6geqvJ+4GpdYBwcabKsmiLp0OuibEa6+PcyDcHk4oIT6aLVLJq33
oTsTEIgVz3RWyJlHRFq7jKvuP68EE8l8m9MSW4HHDN4DkgO7EstYDRZOBqWP7SQsTY0dCFgpBolR
hTZ4duDB2tRDSY8QKhB07zTuc4hdk+ssGgdHsGrKHLd0JeCZtlT6Zs2KSQ/m94wFcaHGaPjrz0W/
/ex1wSmlN/nviA8HfvfnaDKV6Hp+6pSMmogi7JysYwd/Tv31Wlp+Uj6eJSPdJ3aoognzifBhFC5D
AQ7ZuiEjXzNZAx0tx2HTriMOqMtRz3Kl4NIFDsK89KjGypO25rhumnHCRoulg0THr9dn5kD2/lCL
S5lM8TpZMNyBTO71uUnUbercFO2BB2tjDoI/ff42zgcWFV2qkd8IhqDHfGOxj1khVOiUYcm1LsO6
tbBLUO70lekhwAOZCbu2oHP/Zmh87ydNwjLuLev70Aj++xUkFalorG83DaVnpbGhn3Zj8Vbgk1XX
iWH4a+yWw+EpuL30RxSNI3aS5hAnNxDe5EBYJmpBap5otxOSLCj1RFNjPCLTggBj60UbD754yToi
UOoXAP2WRYN38lLLR253q97XH9xkr0149Wf+KPpWG2dfsgxGLR+BqG39nYHvPIuQ13kkA0BqU9dg
yFPelrC/QV6PN7bE2Egz1mlg7Swt1Aag3VxjxzNhsj2y5RD+DJTjEGJKEcQLGWIpE5u5KRqoCnCo
YomjNC9MCsZX1u+1GQme4vOwE+kXekLKXwIYx9GYCZNxL7DrNXhis7azK+iy5Vc4BK3EPwXxLcts
i1ZiHvBX25w7kul8pvF5RyFgeh9OklRrdqEpD62XptY6Xk4IEUcAqRacx7g0BMhaG8mw4YHggA31
xGFVKKj5zrO4k5qT0PtMs9sUgRnD6v3UdGbNK7DFg+rdQy6c7N5lr7wUzrLivLtxcx5KQMhqBgAM
gzUcNAKGMfQ0VDQ1OAbwd9hDNfuzgHFo/SZ1cGcYkBGtf2cMpoAutSgFaoaxx0SQ8DgQjn5xBkaZ
UTB0t3DJ/AGzWk6EdXHCFTv2MbggGUQdPYEDAsUwZIeQc0uGLWCzIMUoYVablstgQEmcrRnoSlWk
OgZRlpEv0b+FrgWsVMWFZPcu2dTUt9D4pFLgeUrSU03x83lxD+nC0nwfFekKPGG9eNEAlYOnnvqX
AfhFObuRtMyYjKDIupxsRTnycqvYYlXefWx+CzY8IVyeyEJjmzNQFLc+5berfLXffHtGJKBsr6be
eKsjmN1XgF8uAy7aaIdZ0h9fazSD7Q0FxTm8d/osZ2Yt5znJERfUG//OLo9pjNwk+JcFnsRxDGzs
jXY9b86XmbwlxAuVKQqnrokBvqP1TnQfLeFt2yRgHzsTlt7GJnAKdg8mZOjOEiPb1EfvbIxaKOJB
vbztrGsu2q80+6rkzi/Ik5LXECoC6/J3r7iqUwJKgWOtLIyArBf7X1NOrUVCoCkcC+/og9qjKK2r
AlKMbejNiLcN1ohY3OZ1ORJdqNoXzJIKSridbnkgWnfCsWOletb/Bexeq0CQUNSwhObgOMEhtoZ9
kAu9Jh2ZoNtDF2rsoLbOKY+28FkR+NfTyizPkrM9OEAYBSqHJyG4EFW1qKHwT/Q0bnfR++BIw7pC
sKZDTK8P5eEbGJ1nISqJ78AjlkGmHQM15e+7RjOofseA2vIdC2ODG1PjzeDujnXmJ0sxldUzyH4E
0K4vrsesTFt9dxJankjY0bvOacAw880SnjuGVrEkF0NfpcKUuZwm+hqdRCljTNlkNwjHvdUcDryX
Oq/UsrnlLzJhfyBrDoSg8lmrcfYn0jozQrr82MztwtQY6A6Z48m3LMlE0nYSxELG2743g1NedxXJ
7FnPB0MqC7+BmPTMv+3Pk1BUY4+yjFItLyf9ElZQlFbMShI3ejqDqhWTqeAqO2o5psJbGLilyTKV
r8GUbAvtA+FHXiggfxPyEzhSWdjCgkNsDmF+EV5KNzkclTXWv/X5YZCy7jKGvwAzD/dMQ51+G5dr
omz7YHZw8O5tLIkC2fpa8ZAkUZFvriyUPGMws8zRpGHzZTK0MKI5D7/3poas63IRmm8VpDLlmIWl
M189+tJ5IuPXVJe7MQKAbY2/trdRX1mggjSRFCsqwqxJpDdHWz+O8qXoqMU243jeqFtc1CVyKn0y
iksr1IRhjAQ+P9pXE22ymuoiJv1Lag7gpmJTFAE7cr9Vx/cVAr+0Yfpy3/iVwG2sGs4CC1m2YGMV
Ib4A0LQUa395EkcQoW1joDoRz5BR96zzHiO2P8f5ftUN6sLBKgf7YVXBivBA5tBFYuf8OUY91Pbp
sUZyRzAjnB+lcgvps/P9P60AU9MYb45QcYuO4cFIJm441irG6lMnaJUgUIWJFik3PrcsanTH28Bj
28sqfBCdHsAUKo7GGGyTJDTflT3bdydxa+NM3qW6CEuq1dH4Pd6N7cwBVvgFIpL0TMwf00+nWrdP
FcEVxzY4hOcnLUL5GTxToraA/U9Pzz3gntw7o2wD2PqEscDxoT32djWq4jhpPsu15kHBfkIKljhY
WoeQK5+pllFkBgmQnBivDgZiqDiNJ7jWVezJxUrrKeyB5Kzc/4qjU0QU8fl6whA2ySofPh4VyE2z
Tk/znkFdZSrDTltTOvwd0rTSLpJBrSGW1/ZDFNDo9tDICnm6u2JXCj4fREYwU28ntkx5swWTipb4
N0qTj8aMDEn+9fgC3vskdU0dZBjmuxehyuhsnbk6c0Q7J2+fzXkeM+ei0hxYyNQKIcyAC+KqnJTe
vc8+8oASnm9j/IiNcHQtGooeg27ZhkWm3o4rimsQLz9sfr5Am2qSBoXXtx3L0l8pPYiwfy4NtGiK
2ogS1dePwmUyIGdt8tqpXpWI3GYUIV2ala7A5EhZKcM00stR/1IwYaSZBqf0s0+BFyE1enLgh3Vn
elxzDCs6zwb0INDal3xybLsruo+XFBZ1IW5UZP9SvQ7b4FF14Ks64eIuH26SVzKclwu6/FFVy1Zc
77NxxX8dcvKt/wpxbbyQVYVlUfgbq32if3uuH42E9aKA35p76M8a9JkiVIjD5DBsLmGy4bBuDmY6
v45c6PfB26JS1RmnutR4ohJQcbN4NDHTeF0oBp0p+DOm7ZIL0N/oTTpbClyUYWzv3vZrHu5l3t1x
l3nG/Hco//byzMmwWPo+TB9XVSKrn76fM+E4IAGWaffJHAIjsItw7264q8/MU1AQs8tlCT2LqeZ8
jEb+EIi+CEZ1ieznyot7eSkprn/wQkwqAA2eUhdINFhMnUnFgHMmw+DI8Y07J8XAyI3EmmwiP+BD
UfBBWhaEyyOyQZFV/MKc8mE3mm4/tRYG8u6TMkqHWyqeyUYM+8qUFf9e8g6gkzyoEe2zJeQIp+kP
Onp9YwO6KQLS8G/LrG8EM/aQwqUBrQ8+9XTHsVA5RAYxlHYz30m+FZ5D3pr+RAKk+h1r8jn/yL07
oZ9JHfvjh+w0x2CGRlUm2kbc+Qd+16Ie3r3H5p2mg3Pl/gLIXPFiR/KJh5kNGAZpr6lUlLhwhGw9
ZKe4p/T2gCQBQ4MTP4PXCh0ZWzFdTEV8fu/BIVkDB/z/tT+Uka1wdCj1VGhfIIYKdhZTyMCNHvPM
Va/f0LFu0zMkF9RG5ATQc/pb0aKrK9m2MnvbrOfCg1TaAymYRW63rPU1oL3vGLgk6lLqmBoR8I38
Ku+6fJb/GKaFozfVoNN7GU9fW8dPvy2RcuxIN/7cP5+CMUiTX/nJukRcXxG1C/XcRYtJg3mrgh4g
EqV/3sfqPZHnyVoItIwylVgZoZhtVQG1kfIbd2eP1E2Z/DHM8HKR8MGDLNxcWOCGeo0ANaBwA01B
g5OqOJNmtht1Hz8cy8m9FjqIxDlrR8ftpInUNoi1RfYHakCaZfDxn9oy07BPKkSwJW890V3Q/ZL5
G773Ez5gSJQB6FQpEHtyEKGY4zpGCF7/JRI0NdDNeDD8TczQAlRIPc//sZbsZijTDo1A+Ti10RX5
PAMwX4wuo33Wp2uc/QMLZW/RSzEATUNRLvLWdkoO+wClMPXuWj4N7kK5eBltowovqaqsWEGX+nMc
XwVTo5qJUxOPLyDATQr/i4iZwg8Od3OIsADwW2qPfICMoPUvnMick26y22nJGC2ULHo0GUbkl9HC
0zZ5pTK4t/oK2I2mW6X7Npb9b2mPtTD4fM7woJNjVno/cgH1LI8ch2BSEmwiAoak4DJiWd04A3V3
TfkHo3xWCejxouWV4tYKigsMkgjUsKgO9OxLBGb97z7zaL0xK3IAUYL9+VZtbH7/9tBih+fwhUen
BMCaidye4kmvvFg/FXl23mIfaG17BsV6g2o0zyd5poCHthWU1I5aUqy/Id3oKt7smybNuQTE7nf/
Elr2UMItCmm72Z65kyP1aZ3qeIT7cOqdb7xdMyEiRYd0uuCTrTJ1QsxM2TPA4PI8EwPItlPay3x2
rXvXupogLv8DX3wdzYXn9DUvz3UJbwpVM99+ubxZKCMai4j7l1G6lxxq7HLq0HykLBuTaERtskyc
5gyejHMCkLzpO7xD6jVCGgISP87Z4GBRgsIH3VQa95UGK1GiGwjQ1l9bAnyXJzIBDS4jE6CsSDQD
K2WTOHsdc7awXI2qqLHQY7Mtu5AuRoZT+IriwHElfByhXQD94/Uwz6z2VA6Lzi/t5kfoOr8P8tiJ
NcD7nIgPHNrxKAzk9gruoDHk4XASBz8RNRdPgH6N/9jZtjk88CT3SyR7U4fgX4clbrv2IbhwzCa2
9x6F9xfzEhxqPSFATML79k6fz1bkN00BtUoJ+mRB+5+qUenrAyfiGO55bpIVvgB6IlQi8SgMaRqL
pkqUFFHG7m71ZvowclgresqVYSqtnYSEhquBLHHJAvm/Sb40aP4NGQ7qZfkKr7dEtIHbYkOL4wBv
NPvXZVUXJI/cfO8KYGx6r0gO4dgE0CqoQcBTBYozu3qKlBzBtOZcs06AlXSeZNniGZcZuc6G0eyv
kd8FweFb0efWDcd6ddxYG/g9JCGNrROX7y3Qs5jZXI11PhpRpfDXAdCzZ4lFe3TPztPnjt5rOAzW
Ed99WdbkXVBN40LqZVWl0JhVTQUfQBZoiHgB4a+dqHzK5/VAj+1Kg6IY5EhqdeNGfqs3bO99Wohk
4g/zbzP6VI6hukr6gI6g6Sm5zC0nGh6rDI+QluExA2a41eMlYmZRkJwJ5HEdSEqoi77LBLLFgzXS
fOtuTFRB6YpePEvE2d/ECLQRNVsNKV2r85eg3bYoljyw3TMIsZRYSckQjt2nv4nlCUsakKbhaiXc
sD0IXuq7KWB2N+3LZ0SsbjnT4Ln/jmXhsvo+8gN3hg542khLmZaJpAuAgM0n6GlxPcvNw30tVlyG
yEkedYxxTWX4P2WW4sXjHNWPOxfLNT1LuWSEbfCyMr7qMxpT1is2Edu+2okfxQ4VimnyMLCljfcJ
r7hVCy7Oprg8JSbMKokAjl84l60Ow6b32V1ZitM256VE3y042o+xRBQVWdTaXjqg1+JDUmaGMKwR
JlLGodf6zJNtvP4LtN6fK19xHP4/WsKfNzfqLpIs/Rz/E/ZFvFnzOoVPX+osYVDN6avfcCmU3ZpN
V0Mrt2MJ14Cjh5z8em/368iCtbdv397Nh7ux/t+B4Syx21o50lRuhH4GIm9904cmzAfhUueFbkP+
rKYqf7lKFB9E+auL7kcFlA4Ge5RY+XLjPSeu6xM0bvzzjilI3MC5N2O7isEvy/ceTRTabzRv0g5W
yIj94RJyOXmCIBZhJBGkrMDoug2nnrzrnVVqICE0Xh4iBjC1rVH/snuRitP2vzEvr6kd3ESCe1nA
v8UF3K9cX4YM1LS+sZrm0nFAwQ8z63XEj1du//OOzqvZ4SPwm3gUhISE5p4YtJaShve9JdVjkQ43
x5CYAQNHo88riWhBGAJdesODJre3GRfqPnlW05wWgbGL9mvxyS6nA8u/Y+DbANxcAltj2i6J24OC
9T4SJoo0UkfDGd+H/J41Pll48zG723Yyb1wxcMUlGxMWRg2TKTkSKxVWf8Gn4SZK8a0uaDpT+6pS
W7urWbgYBT+LBH7v0q/VVwplBYM/HwQlJmwZmTIGhNl9vY7uPLsico7AzZJdvhkP9VsSb67OtxBJ
oKXV7Y7CSjNzPLUgCAxoldj5iJ+F17Kils5tazbtsyknn0oK8ThJXsEDwTfuoIMoIkPpmddnyB1I
UI/sp4hJ8xrdkcFLnraXaC2Q+BwXj7Z+s1p9UAQMU3yrlJ7mfxOQceP8r6SgSOPecLHhciq896/4
NoukOkdbRdhqgU1dUsKH6X5qqsHpDF5F6g5iZ+vVyiQ05egc4m11x1mPVAZ5ry2VMbdMHJfG6Lt8
jcRtB4PyxUEyHSxIrqsCWV/kNr1W9ezeXX8AcdE2BR4x1VxIxh23G2kMTKjaBfgvuZgDeXIX/VGS
wARDW7tDFYV6gc1u2/ueF/QiBfsRvevy6738tKX0W0lQYCSrl474csoSBoS3ytxy5RU8+aGjxhP2
4AQWPjH8vq/1Lb5p1bnNi9dQLXjqLeSochNOKMxs4TiKeL82uSvVJcq6tmnDG7DLEzBAk1/yqFkz
4oSEAwE/0s3cw5MHf61FeQVGhJsBBHrTmDCc5NdeUcnT+e6Y2YGTO7fHLbA4+x8gvA2lyqZjKOQY
ZPCwXUycuAjYWnJTHumRIyhEeqgA8fb77FloU0DPvxM9FI5y8ejzeod9VhjsxDUO3XBd2gULa2zN
h/S8IxCz/qh6GYztV8RjsDzkp90Y6/jSjaE7B5A2uJyZ6s6VC2WNUQ7zZt9fRUrwneK+QzvfnEqm
+D96ny631Ec4Q4Jvt65IWBoC097UxEabkkM9T12av60tpruO6hJbHJyz5uBQDvEOdJuI+VJB0KhG
ESH+jGKoXJJBd/ae1E0NxEh2buCTbRYZ1AIB4gUrMwoCp+BQjKV5kt+s0/VPZvtzDbz/g1O8Eyie
MJyxH+hVg6pUv/6a/saaN2U5AEbEKz9RAKI57z0kFhIZD/JjIUf+KPDBNZXo+3epb9RoBXWt+7MQ
NnAG2Axfz+FFCMJu8CZXnyH1EaVefpmd7o8yO8msMu5gxJ+YSORjqlfkbukPj+W2QSXBx74/ffql
NQQ+cr/9pMZHDBAsHQRvVpsSLSdzqWi4+55GHUsZcvhQnj0GR8h2E1GOiSNKWLvjjFwL5Bi2pwgU
+uqWm0yUk5pjgrasYic6eRNGm+g5PrbgKNMMZ7w18jaErPEuIpHSs9e3LuzZ89t4DqU/y/fsSCdC
ztZlgqexUvDalGS+wE0JTs1cZgcIHm4sU5p55OcG2D/w6TzSL0Q9gQBqDk97IK+/CirMUgZXzINv
eWUhGwiWqQ41dzEA2yK2IVEGX3ExkyBxj4PgQjTJrc2r+CuBZ/zI2d0xBWC4x12gI/NW+pOlk3N1
GvBUOWKev6YfNISDs2gObC9bTqRUKs79zG4Ed5i0Qbeyu02tbH2ZhFzkZvBZ4UzYPLg924XELNeN
IeIph3G5QXfvpRL1vrUZUhX2CIuyfs3MfNH2upewgn4Hy4IKNdXq74xPrG2W2pwMSDNRWypmUnwx
BTqwtDIeDQpCtCeD3kwXP14A4hXzvDIkMa+gCOgVAOkC/pScuhewvo+ERbGpmCMUnnLeSgW2qRQQ
H0yBVU1q03mi4wvcJX3LacrfUn2uRWCBHgpwEmiC8nTCgiBdpIQBykyl4VhcUol7GuU8+rNVPZ8Z
xbNKP+vj40hT0GDzoihe24wEmLGUsI7I9XyYOIsVECysxtcFXWBSa6B23i1++jtKzgoGPInJR2VU
14BGAhuTcYB8BfIpK3eLci3+HvW4wPbXWeYqQ0uqfffizIgkkNNxEHf2FfUCOkmDkwmKLj+yYJSE
oB1M60VCfAhGj0qdHSZbOpBLh66hm1Br9uqT6oqJz366v1O6UJP56Nb1oFgNYrTpeY3Q+8jsV6p6
4D2FPzbegaski7KVxBihCspB1GxQLTJlPoFUVqxteW2JUhF/UxK0EnwuMigfNYYITJYfDLBkb+x5
Z1gAl9FzuyJXa5QkUTqA7XEpwp9agwr9ZcUxlQPpzAxehhYV0ccekuWr5djfoUoGcel9SpzpVxhv
5v62xMRCvuqi542LZaH6DYCwQSL2tjpRnBOJ3EN9JrFVcbZArpuD94c6GZVQglQYOoNuGOCD9Gjb
k3SYXwmhN4PwQfV3OmxUQdL1UtLcs74eD7iABDqCMbLw+tjw/NsKbKAxcbAR4vfLWJtvcFHvoFdJ
nA9FxltlWFUAMdRCme1S05auXEPkUArM40pBFD8xSyOtv6PtIut6xZeInYJayFbET0THfDSkpAV/
hS4MfhruEReY5PBqil6vOjoYhnRPd4nGFEVTZ0FJquDZJK+qh36/F51aDtqOU1YyIIYlAoeA4/Ii
P9YqQaUP4KTG6nK8/6N6e1vidXVj2wBeNVS7uhfot0KtLFVzrzZTH0DVWCfE7Z0tLJc69AhGzdLL
4QRR958wxECI6fepFLmhvLSTKbasj2eIgdZtqprJsGnwqMDPL8ugcuWojZq6vbgYwT9maogaPJ+9
QfpfUiPlm1ZuRPEVTIGYzx8EgayDEyxjCHZ1Ytblw/v53ZQ9iwqTjkTeVjPp5vlkXMlbQlL2yvnA
M+gvfyI6bOlbE97B/vF8OjTCZOJDE4coxKaSXPnASb13LicsXkTzn9xNgmM0eZxFtbMrC/ZPmWPJ
pdgXM6j9kYneRVx/1tH10xfJa7MPF0UiBwphHUvAvyYIe8hJpyl/Tq3oYwPbBaFclmVGkKtOfR+x
f2OwSrI/FjYJ5PiZmhcflPcMxUjP8i66TmWR4t0sFv/btg+IT7rdRXVV+1Mn8oyVoGQIVRV+ND+l
rfffG0MPNH6RmcJPq3wHC9iBhQTimyPi5Or978YiU0iAQQPIDVDQzCFKvMtep4KkADZQdDfPyzEz
rrzFPO3ByeCaOCQ9PaEpFuAmM2tjGmY02aUiQcKYrjO+GzzXkKVGNT3ZebmHHXEg/CmQyOIP5jx3
jCruUWsjb5qYr41npnqyJBigKjWeVvLjrbIwri7BEtQ6wpgxvzWSSWnCkRtRL/1LRE8k5CQ9yrur
BngP8BF+0iWz5U8fuySymZrQT0x+1fNV5PNDp55uKTuOsA5biy+h1IDP0jZP7l4RYER6hODta4PA
GKaT7ApB+3wWHIVAd63atqAUapL2eXnxTD438I3IDVFS0qCfNAzUGOYZ//zKHUdfyq+ZtoOBvBo/
GvdAoGyDLzi3Hn3dlR5L8W0Ztrky5PhTr4RW72fg3fYK/cY4UVzym7FiOuk3ksAvb75xWfrMn4J/
YwOWsUYmJytWbe4/Klujm1rkBj9IkNizJz+LcoEXAN4KCHjSe+sXh+yDrHf1kSIZh2+EWfl+fVwC
UIIZPJa1sD0PQK3+nD0VLJqSoAWyRdTuf3yzwxr0MOlyKa8qps3hUHeRVWZtAB6zeISeuvA1CAh/
KKqJkQxSswuNehJVIvpTrqJsTjJIwvkAzEwmWmiGbZ6LUnbeh6eu05XWiZWjSSQdWyTClcbzVs8Q
9KLlXIojFfJTlyJl/Vr4vUHi+1Un3zU/qTTc0zYlIdH7D0GXWfCHHvzik7gXlmMaTgzBY5Ii0wYA
RoMC5uNNglPmwObAoguNrETx3RrIrXJBazfVpz93r1UBgnJTbOUSAWOdHGJNIyPNHqHmxN9yKDh/
hbW19Ul5g3X1Ls8iiX0ne9nwZXMq/QiQO2gCbbgR/n+but0txwkpH0Sq0FC/rDfyYk4DYDNKZhnP
/kQioE7lPTe83IsuuCnedrfHL3CGn2v7o0np3aC6Mj6kVMSyUz3l/uRlQH6PgDjIECjWRj5XE2vj
Cp/+M7nGa3o3Ze89ScZVl3Sq9QFQgjDoQj7XyeNxjimSpKUFGhKrs9ymR5qxs9sxSK499vZVcxuI
R7bhzg8sqUo0wUL1rGp1JNuU1Y2BSOpB6ehHU++RJqP+6hTyN9Vycl9TKyLORrXPx3RCMwm+isKZ
MomjxsKj0t+q82UG0aJRaHO1LXT42AmSlrCEz1T9vy6naubjtk809TkLisbZNq1EHpn5cIWM0LY/
2qZiqfaIW2pNZgdLMPdNaPyU7Jq0aTMb+z66kCvZjjenl3kbxkGr4BlaVGfdppcbwBl7xbZarT4W
2UvbgN14ls8HQ7gzSUJNzVLPlJXy45XVWGMuGy5K92s7pUM5HqFwizKfJGW5gHEU5F92FI59QqUJ
VVYBm0pa5+IxOxkUsZs+l0myEQarqfjUihLW6h44h2pyy+R6NtCCwEg5Bp7+Pea6r/JtkdzKAzhe
J30q9obVAElszwfJiEh5yWtEh7tRZctLU5J9wIRa6IavgBK8QPNCPEQsuVsRFfiHTddhPyJaQwZv
Mx8lyjSrR27AGCvGC+Elywqf4wPFtaR2CDK21zGG09Pi8oAaUawEvuoyk5y2Ud1n9rhwAbNni+Vz
IGtsG36hLpn3U2Kh9p0V5JV0fkQ4mGD0vWu72f4Msvirc5gfC/1rLxHc5ej9iEfhCtV0M3MM5McF
4HUTzLoHmfj8LbMSGt64uX+mCbIU8WfX7pCvU3UtwI/xPsMKtpa5pagppvEnQJJC/FwM1zLhcd7B
QHGSEMlA30+yvgcaFyOe8YCbby5NKuzGsnm/FtbbvVupBcOK7Gn+LoWSr5XKyVBh8PAMRoGAtc97
cAAnDWUMHxM3LYm3DysnLbBeijGgJ3YJIlLr7weq1G5qNpBT0u66+7X7rTdnxxfFaWMsESDN75rq
td6Be0efqweGy+FxQdg8COY/JSoeYATydP+d5yNEBYtg0gdNaeG05ylGI6hq7ioPRnxnGDJWCXwP
ccZjGEjqeCuIofPREPKNlLOb1iKyLAgT/BhBZoLNGUnlwgdDcj1SmYjwkf6zFghT5kjEW1ZDWEOg
MPPn3BjyKUzRRlH2Kni7h3TtPNfMxBhFZ+QwbmEFq10/s/O3SJBTePP8CB0qGU99+DpXA4JpNkWA
xaZ7mnnWPBWNhYJie1CmBYYAq0YWaWGAw0uGYxp6WAHXhUwGL+1KN33DQfqsjeIafQJqB2tA8656
s7bGirjna19cP/UJHvmDFgk2Rn3d4iyqkTOFZLPhJiAkL/vUmQ4fY9zxUWMji81xC6RNC4ODJTTa
DSvh/bx7kys6Im8bEsA5i7w3ocMWdRQQNDehntEsmTN2QtQwXlOwCgOUVawS0s+P1wfn1aU1Mcp1
vHk6aYvQbn3d48DBGxukgpJ+hd+EZTYWapMwv71Afk3eFyjQwAm6pYQFAhf2VydmY0jtax3R1ebj
49v1ZRQjdrw6a3jnxrXzSeYFsArGN1Tt5LFuBNVfVIsb0F5wDKx9vo68c3zb0+GY7taHmfEvsz6f
iRPzLq0Q7sxpvAtk/SdvFRhQKqRYI66sF6gdWungWyK8IILR7GiKW8XNOfCWCExzxkiT/2e+qLkX
/5DDR9BpJ04eMbaXb5TNg5Qa7SFN3i3exlwQhviq2zdXZwvHCoVjNOYzUw+smHmfNfpUDkoXvTJ8
UNOOERK3VspDhLYqlN90Ad9uyzyKhJAXk1xWXzrgGIN6UMxXwwPeTpH+iV0W3FN/BG2PCsnHUjmv
9vKsFvdfA1vBGK0x40OHhUa3tCyoQrMw9FPpptceeTYV/mqta/siis3ZQy+X5Ndw/KVeFGygPktn
q5h6BREV3LmixkbSqjCNfETavfADQF2WkvlF53wCV/rYwvXHmNhvH017UJMGbV7z6+W+Ih2vNczL
FrAGHm2M29ppET2yiVnhmDghfGO5jF24dTb8nJQ7RGHTxTJ7vsElrsp5sRAHfheRGnyKNfLBL0Oa
WVj9yeJs2jBCaBsr0CmZ1CyxROUBbKv9YlAYECyzM/HaIgciGzOa62tWy7RBw0pQ9kTYlLCkCT/0
ZD0gi1R6IfIPaS28hlxXeiIOBngEN7LPR28y5oWkKsyeNkn/KYK5xSLCVLWcrNyB2lFt6GkbdSs3
2Y5LFqVgA8zRHie7g/Rj/TbaN+HwcYGaO3jhBqmOXFt9S63LaphIJ5h2UTKo5qxD+kw52IWfA9tl
RCEnVbwcA/w0cU5Z+QEOlc4COp4LjUN40tINQCo0b/Y0/IttGRJfczRIT1K0yfI8sXrXwiCYEV5d
FSFNn3dl4heqCT38PW5KpvRCevu5cqOW+nRGKEJDQnFWU1Vay4akZq6x+6no3mDmO2vZyoEA5BDy
th899UzrX2WWDfum14gmfqIkMBPzsjP/PaPBvkSPb2uOQJ7KhQgwIaaYRhnjnFHY4HAzRUAteB97
Wz9h8nTKK9mhd5E9H4IyREBAzZLMkqe8KRVITJG+iavZq+YEsMxbpxLyRrTIP6LC4fplKr+0iTHw
SeaWKd6kBl0lNeS4B3eqcqSKCt+UTTIPHlpx+zKn5UB0vufoxEHwouYa8oL+YGBQTO4AeGAYk2y2
S9RHVDbNf/VohEwNbKdD5GAy5ONyY02hQNqK7JfyU1gbW2xlwgHRQUxvOPwHs4hZlaBd3Cz+BOct
ALMqdCD6Segi1MKOT2s4jRMklQkduZD81LqFb3OnLOEpyjp5bPg27PgJpqZwbDwUjtlglA4A2RK5
mdSUVJS3UyO4Uwkjvw2yPgcixoLTBb3YofC0EFDi27D9nDohBgRsjoqn0xxvDUp5D49VQ+0BK46s
TLdQWQM+6PbWLgz4RNwgpuzjdfiSlHeHAj5HUAa+RpZmz+v+w/CYf34ulvamDQMC4uCmCs9+YOr1
ysBNfFTATKi2DtM452PmgUJXFRAFuQsIi4WkU6aMqnq3rZoJpXpLdtgEbtKLmhggq8Y7NlaTtBl3
cGqB/xqI60To1yCMfRGVAfJCpLgJD0i0RHkvQazw1HM+LJZpOnOnBrwpFXe3W3eF32c2DNfbhN7Q
Ofu6254wpGlupNl3FBFaq9z0ewhqWzHhsTjCGjYuSCE/7QD3SiNxIcBFpsG/8ao0O0vLXcD51vUe
rUycqb8Fg3vuDg2Ho6E2KZhP3sYjZed65O0uN530W2vFbwrD4dmuqphhrqBWd6UlW4sHpOIvR9CL
87NRdTDP0hDPOf3km3Vgjvy32m8M4hYJhc2ysmGn6V9LxH0rkY9UL8GZJMeh0w+F3NVZ1Qc7NGZ4
ji5mkE+CW+Kz3hHlcNad3eP4Yrn92vr4WLwSG5sBX7+JPtrbwJPskBqEdAGNNGzC6dFDe/QWkQAp
tQh+vD+9iqWJaIAGtO/VBMTnybllNKK17Fva01gpZiV/8DVr/JUTz/e+43mLpiPSiVP0mABPxifv
9ASj3avbsxcQyUM2vujkhtRKNMz2SLyEXWtnrZfwftwipBITqAp/gk/MK/VIU+JcM8lmMPl2pprP
tRt7yEpBtOKj+CkNAQXlzKriAmLBhlLhkT2cIM5y6Zj76m/Cob4i+t4ZKMfBzhv1pv6SaurSGAKW
4U3DdyhD/jB2+8X9BthMtGdIA2tuwGzapk3QwOgrtfu8vLxj07q6xws/uFylDzmYStNJL7RSrYMO
tGp7hzlj91rnZ+ENc9KVVSbAN7YfVHQij6KNg9+WcphGfLnmsvuOHYitA75gvv7deXwCNuf6ULt2
S7ctPlIJXGKUy/X+VE2R91xwuQ3KGQNWLf7pn47pxHpySKXxGr/G601CbzMWpt+NDg5m/eXqFYGl
xsz2IWRSx/WyXl53UF6NyfcQocIhgn03sv6weux5ckjnyjU5hSWBjXhGXpuptsFQMTplDhn3eF/9
4w1fTQSTySBz5xdtvd6XhooV8Fj2f0gR0FdqQIG8QsBnllT3Fk3LXQiJp7+4senWyuQ4VsP/fpfD
JGJ9csB9sNcrVRlx2GW176A2clF1pvU3g9npai5AFYtURDdSOUtXvrAFvsgK0y7bMhTNuYY2Jybf
JNfjqoojlV60acJGu4YsoaMHKQBTU92Zyk3ecj2GbkKFfa723QnDAEp91+pBVgOE+eb8rRekIseb
d7R4ioOoAWiLaAa7/BuOfsalO5eykOw5yiTqNaSqpMD0lGehsexTJojaXbsBvX5Nj/rCIy64OHwI
Bob63zw4Z8z7v7O+OXCBglgHj3E/4iQpEW6T/sSs388igLerNuZoNKEHVkneiiTYg3HkINsjuGDU
jStkLApFJPdWDQP96Zlo59Rv4IGRnNMaUV1X93aQxqwOnKVh/RQA674YY4SxzhZRLUAbLZ6RPy9L
Tn+YzVDLfr8PiwYxQ8JXFnee1Pb1OuBZjgxE+cMBN8GebKI8uI+fmtMWYf7jE6/87jinLuiwhlUq
IqtAy0ClU3qvGFq3qiEIgxjNlnfGN4rzOxnx1231rzQAsYaIL+81qyRnZShxNes0YitvaSIC4Vw+
Jh87ubiWryJtlznx5bKjLX5czzkN6VTkn9SSPgUzD7bfnwEXrqqzBvCY4Odb8vjtW7hKoprVEXHD
j0Rjfn7RgWUzV9EewCeXu49j1NC7BpVgPUnhxr2mRikmJ/JhM+FgbnaNCz4oJZ/XFjPSXcnT2l9r
nfq603Uu7TTJAqRN1ga0qjuHADg6Ku1tI/12oDi7XQcIda7UvwRu2AeRWLnDJwEUTw9zgUygXrwC
TjcVw45r/Hs4jGRE0LsWymipdb0HFDtlGjhRKS1hlj1ZS6JHAeFsdUBoMrv+EXbpRh79QC4YFQ9b
oHjSegIMs7KSZOEvkpFI6rQKsfaQk6sQ9cqfuNsTUelM4zoiWDothRbsMwd382fqKTe9iIbc/79Q
FAhLrifs7pHdzw26mozRghN6R5FFYD/DmNS/fXmTLURzqMSHsN9K2yqSqXpuJT0cvUBPA5aNVRoH
sF7mkdR+OIogSGriB9InzYqpiYMhqZAFM6yVnr6/nIIpfyuBqksoVWB0lyKWplUE0+xURoSqGIJl
knIkpX8miMHnb8O2a2RPiEl8zfFscbAv5I1jsyjM6Ivb+1xFOFDTqjlFYNnKF6HC39hTSZucd/Lp
uB6q7nFLwfRCXXLx8rc9Ztf/4PuIjU212r15JdJCnjidcQA8QJv9TiFyiD3pOzUOSegMyMB1hd50
gOfPblfGuvbZaEztqkmZjf6qHTRuHl6GqrIMU8jZCuWN79ciayXb5IODU+Rm/TiWgZInvcz0FUcg
DOwaGJYgszblyZlW8S1B6MQl74b8bVZ+iC02EDz2/SPZG3l+x8IIbUkuZ+m4uCSDMagbsIcxPj5H
U16CtCNhw5I1Kd6HhwkMkWWsGfaBFldzcKgQp/eqyTSNh48z75CwiwvuOPsBcQeaAUAjV3x9UN28
8BKN3wscFXkA0ZkwgtR5poU8thrrexuBir2er57UK5G43rE1U+L2kExDKFyZvC12qw7OUnr9vVu8
eNutM2pHGQAMGuaFGDLY1TeNUEVi/nNcyTadA/THg88yFJnwr59GdbXcy3RTXMGV9fojHoKiT4CO
l94KIRDV2iuhQRpYLS3nM2fyPA5inI0S7L2N0telEUpwoqyIpzjG+7sbeLOUFJmvtMKCc7VSkAv3
SEgKirrA+z4PZCqOXaTjp1jNob+Wxt+iUhmdAK44iqc8RPTZLDvC2Fd2KhgTd7Q+YQ6ip5sCGw3u
D39dCpl+PuiAZe7kXpUzarmjhZgAyl8c7rHIRmgDDiJNJMXi+ncurcfCx2OGRHHuxN1E/vLNSZHz
1u+UbHubaAB+EAB1kiKToAWPuqftWSOncloow/zZKC+qDxkjuN7Up5TtW7na+abU3BxDcfv4bt01
Dp018kPjTXG0IV4kK30CAcIvVH1Jy/KF8tsMlaWf+xb9aHEHu7WBuMt8KCSf785DHCOvLWbX92VO
xFaft2d7IQvjCPf5xCt/QvozHVH3+7NG/htJCYwZoTdloD2DoRGtwbSDXpEX1qRpcxsaGl9Xz+UT
o9ffQC13ea4tBWM0CPwnQAFSBAvFq7iO6RqPGCTCRQ+F9cJavlEtEqotYW0RNR0ttewHpbib/NhL
M//EpI/0RoxNwujy7cCdStAxD6Nawn9aa2ZMeKhgaK3oEIxwn/ygfpCc411TsRiB/Cz89oGJUKsH
+WowizlhPifstox3lThxwbp54ROQ67T23tkk4ejzS9AXBmG+h9oG1YwVlXIFYOPkcz6vxrasDTVi
TwFFhRXgnnsczIwauXL/qDIt2PT0zl8ONGJI5c0uxAQSqW0fWYVl5uDn6Iae8q325/pkIwONiy0m
8SCCPSXX7VLthMOywuyutO6qXgovbHhh4fsGUI3C4BExNReNKa5Jm5Cz1xzV1h5OLe5hnktP7wmN
3hbCilHH4nHLJC7lMFf7L2tC0JDQqxkE3ua/D2/jgLNtmZyyGnkQHVYqYk3Q9NYsaSXeoM2eij+f
ni836Qm3SFKrbctPiRiU4G7yf6Y5VybtmfpuRCylJtHw4oj+W1VWSxQIdQSsOAk9yTA/iVNXfY2f
7id9z29dwRoyH1oKfofhdDItNAm06zVyG6KoDmdW5FBX4ZgNPMqTSR2fbEngHNAMd0Wl1kzNce6e
0s64JaugbJLBRhAz8iSibHrLklQ5sVeskByfJ8GFaz3+dLqJCAKmITzsvlC/G7bqIZQKo1Rzlpvl
o1CwQdx4Pav7ILdZxQxdVuAijxl+r1oNIxjemo7T+GNiahLu4tyBbj7hpSLzFpDOidwdvV0u5Bq/
rv7a9+AyMWoQVvfONfmPH6bReIK1Y2FIUhEL/95m2l7vzTL/vTYmhs+h3S3JUAXRxQi5ycg6Qsgo
Kyo7CI8Y107Uu0SG7rgqBWcojO1kqRWSJG1ZoIZb0DyMXqqoCOkuOWw23el6bghcs3uuZlcLGP0V
n5IhDyyRYPp7j62y+9VharaZksJKudMgKyKiZED7jiudXeLyBr5J7rPiC+/g2/R9UI/DnrcpqyDF
AjfeQ+1wVCCoD+UArwSkAkQ4ZJbPIVVVI5G9wgwdGlCFo/n6GDHNr8DL1Jqnm9SWoeqriBzWCjxR
cj4Uqpd7LCsFqqcD3VeP4J3TgWuyUvdprxvtJXKNYSiuVfWzFPM9CPTw6qLeFlsAh/0/4ZhojoOt
E3zSdKnZxQxcqtl6fMqoNnmWqTDZdQM8MSxsPBnJkDNJeoUbe9YG+2HZwfT5WF8qgmA9PVjkb19i
0QTWjPMK1YKc9R9c9O1cI9byeydMveMgY+soILHUIf2Uq/BC3+nPqWuZA4rdWtHCl2lznr6gMnvJ
1VM6naIZe5Xrg6TseE7gtFC8RkaskeqPTXFJRIkdOCvTA6PH5zXtKw82unsomnDzrRsI0BP/ohU2
f/7OMqvUN2/IIYKwb9bAvOJMw9tUDrE5ctNOJRltjzFrezYcyTKoZr8V27XKBe7uRsvZ6FxjmJ7/
iVjlCcze654H0CAUKBJNQWbdJPbcl873YVbVbD294Uh5uB/70BSfSXR0fVgjulLvA69KQZ18z18s
eONkjotpAC77i/qQkz6/mBGseFSybi3d5guPXUz9mmzkFgu0CLoinnMeoGLWPGdd37nq+/SUCdhY
hZr2BPHpSO4sBG6G6MHIjjJphboFEYHC2iwm+69bzdiPbA++zraNqT6r7YSj6AzsBtCYg3C6QmgQ
CLak8qimHMPguR7mM3HBNlkyAsjr/kdks+81LfytEz51mf/1SmCLOIeoMrFq8N2FZD4ipAKBBRCh
4e+YJbG7z5fD12Ptm0UDQ+L/ov5Hdr9TKgpGEpQYqcqcnvRlyCuwiPGCDleSgwtPYkDAK51TUAU0
+++RSAMDdxclFrk8tzBgcp6cBi7Zz0dR0X9sGNyZBmsxYW3UGEsOuHlNJxJyyWvBeBlvq+92UOEF
YXVdpKR8Y9RelKygNSQR6CXEUV2Vv01+Y5NvUTNtgibZpn9Ws3slPVWTMeJTpM/D3A6MuWI9BHLN
az8Wr+OoQnyxikPvkj8b/Prm/2mm5tbXd0foK8HfoLRi3HaNXkJjy5sMn2DMqczaz/HTNfgKDqI/
QiXsnxbQPKR8C4r3D2Ot6PjQsFBIxW4JdYXsU7+nEq8mX08cxtLkRkBn9u6eWiBZLep2mthc2bxc
FUj1tTWRLzAe+90T6QX8w2ZgGINbTdsRQHUX69QssdRoMHGBIkidvKiAWAvcZiKVkjQx3ZivCKLp
9uH0dyXUGuBG3XjxDy44GxTQ60EtulUooul9RgqNY26NhxwmqV6KUznATWUnbr1wCr4ViDFvH7ag
f4qWiXnajGZmWYNR5NqPUrj/7l7cThPO37IvT0dOeqfPKA0o4ud6D57d9Jm3U0LKdQVU/RVAACTg
HGoeFhAobit0pgjbWD2QWwgzEwVW+w2FGca7L4bcslRNEgpps3ZFn8CyJFMhQfEiUuEq7WBgYTdZ
TOrNeAkSzGIk3xfXlTAPeC1/DyQIYNlbTYNGtFONXXET78SOWlbh0zxzc3Qwbd7MQpsvG2zTJoEy
c6v8ySh2bX/qfwtW9g+IEckevoGR695zAkmFXZWwOj9e9r9IRVq+k0lm0X3QuatfHIe91c9p1jWX
WAnKRtLmp1wBwCpRnXB5D36UtHT3bra9zyLQmjDgHxF+IsOHCZbj/fj9RxWshb16K361I8MxHOOm
fY0QJ+QMJgTvbl+EuJ1HkY6R/IIfBmpITtPbuDUH6bo7wBttyKtDfZIEi7/NpvWMci6tX8QGyG0L
6fQGVi97URhRCXEvtdflUC+F4osMz4K+sLcYoQqC2HAJ4wjd54bEkDp1L/tLOcCJJ8ylKXtGLbGs
Evi3DfFQ7tkI49JORVG/Mvlm70NV3aWXNCMYkwLtHi+cRgNre5x6ajyta9hZWpnKqO8ZrlMaPRAs
R5AyB3Xjkal6z1A8RX3gzgAr4q/tfLxlpscgvrlkM7W442WhDwMmNl3Z3ynSXI03DOJIAh0iBSKA
kLAlKsaIAT2ImcDYkDhzsDK2RoxIa3Ytp2xufZhZSUvdtAMKka/LSYoiq8o1YIalG8QT6Y2svuOR
mYh3yuSNcaELg/yBL4TQcipBnXUA6MCS1jJeZQmVtskUrn6BRlvVl4e2PTjiLXVSXfgT8pGSx/AI
gFpMadZXoroa29WzDK4HzLxJzI6GBr4B9L9M08tVnOeJGpQxAW7FbjwVq3Y9x7RlOpcJC6y06+y9
D7bxvtCbY0wXNP1l7ACvRLIwrss4+oD85MGC26mZ9inKMoHpTDExCC1eRtzexLWlZsCDJ0jtIDw4
7vEtKg5venTGJcnsCKPKhpgriBMaO+2VEa2SLt533MHayDGBIxeJPRhLEhtf5GSeAjoUwJIM6DRt
olYfgITPPW9t7c9Skot6t+ZE0/W9hNzKsB5mjpGwOYz00MsO95/2JVmATspSnZ7S4pYOfZQZJ4ct
/5qlLh0xlryb/bq5QawAuk+Zjvq+SF2SnOvaNyjRaVr2vzya0YslusWljBUi6iGaAMODOfvKZFVK
yE4PWPdhAfa0NRNIwXNTl7l1RtsMe37cYm3ZozXcKXr/AVFp3CWwWyAyArPoosB/I3ptH9EyoEKJ
teGcXdXehMwK2w8w+UDZdmk/F0BViZzKxDh3//b1VixX3STHe26OXNxCicJu7XkHV+C89o4b3fB2
U9JZvG3ExHWGw+rMICZqWfVuThYiYq+pfkMym+D3tJjb6MKxKvbhNaicRV6MovQfFimhKBOk6esA
4B2ErCI2vgbwTdsOrYEGEw1JFdy2thH9TTloNYXOZp0/HxEtthFa+iBN08t2+tfdJHdoNk2CR1Pt
sBHb+lFHkJuHhW/pED33VDg9mRgMHNC1qZyPYfJcCcpNwQaxQFGVV6HR/Nb7W1Dw5OE3OMqe9WxB
bPehpCchVnALqHWaJNc9hiDuNECxSEf07zwlID1KZ6sAWxZf8S469G0Xi/0Tsr6d6vo79CW3q+3D
0crRBtNsZiwKn8/YIxDhvJ5mOI16dRUEE1AfC4krWqWR3lrA1DcN9mCNLMEtpeXmrDC1WasxkZx7
2QZa66VBJBc4iZGWX0xtwRtYmjt1IhIW38n7ynqWmknH6UqeccUCiSSVKMXulSnJU6ZMGU9BSSy8
8MbOkB/CTVXOx4OW2+fwmQKQutAP5vtNPgrsiUHtbFakxTfMOYhhe0LmYBRtY+5kfr556WqInUic
qjob8eL/R99waG5f9zWo9cOmSN/Zwua4EFZCYBNjPY7FK/amfzAmTyJlia8vSjFcHK1+Nu5pDPOt
w7PzTK9p+dyjlcQK5V41K4Loq8colAB61kxe7vw5JWFtjT409+DXqcHV9KOb96639Oo7MhFofP+M
GfTzMWv4MZNddP6R8FVRxLeoRe2P8xM4sHdPGlUVQE7AOwle2Pd+5IV+B56Syi3Catzgq1TB1t5o
/ju5TnW8I6MP1L+wSkXo9lfjKrqPsLsgTwEUPDy4A66bgJIDsJfLrgNu2Q/hxq8bI+cHcluS35T4
7aqyxoXO6y14PbdF6Ov07kk467j+oRFbrRyRyiX2h8zlGgkdMNiIs+aZ93Zhqv+wAMCQPS94ivxq
MChESiNycaXeVMTjLiRB6yMapeLh865v6DuImopNvzVM7CdHuVqnXgwJFRZM+tZzGZJxTLBQNh2h
lfcxqREbFPdYCY698tA2vI3NJKo6fa/vSDFTbvvo8xkR68J59nSifrMaLODUFRxSsbvh1Rqf5skY
aNn58/P9R3Ke3N5SRhBuyr/vhk99r7Q1AOiNz8VOf+kV/MJqWDyyeB/DIi+PWan37vSPjcbAOoWU
NB2Sq9W4QaKqYllkP/aJu3ApgmT2T7MBJDDkIf8e5c+2KzMEIaK2Lg4tWcElDf4S4oi5Vf+Fsi67
jCsf94n/S4TZIMnZMCSedMbR2aoJOV8M+YmnIzJa6CFpFTbzdpdyI7RzyZOHEtLaZCKvb3lbuud2
kDfswL6ooBo9fLlFHR4qIkWCsdjm2INniEhWYhu5CJF42EDT98KyRm+S8stkDMu2/AcjrA+1i5Qe
IOxvaQgoqxKn8uLMr2vkcyQa+CsVRX9lYAobBhrlWMpjzDViEmYvWNyS7ym8Jg7yLE/eSx3uB0ap
DGaCDdn5Cben0EinkxrvWW/iU9qhhQkaTVOfoyaQJUkqn0RrxCOFv5QWcYjA/HsXl/GV+zW3Amym
FXP8Vk/4z7B/JTsfkLieLm9hMdL+WXapiX2JSiE+S/zlnuXSd2iQHzxSYcjw8SNl50W3hgK0gXmK
IfZF2XgMJfoj93CIpmmr1EpL3Cx/nC3oAdXFipdZ15JIjNwRhVyX+v21wwVgna46/5b2/yDT5cgx
zGMYFmDwmxO/Fr1ywnrRpcAnhvsO1KjqQoFtxGxNAHfsAqHBF9AqjPKM8BkheMobo6ZvgmRM9MMv
kMWRko9oYD1CDKBTbWvGV/rlyvtWthBZ29tuJKKwEZBPXX8HP4xwjrXEGPQNxWa976f3wX+SzlxE
vKBQOu2N7WxjttRg+sPtMNn4O5JX+HSiv7gpe4I7A1P4aNAs8iSF1iuCIa6uVAAW8xodYFAyG+94
5ElL/OFnn5oM4kt9rwSF8/0gqPn+Yh2Ea8cq1V5F6Qr9BgRv0Fi3Nzs7JSYw7m+FuOsr/COS94mu
AYR2aiGssHqmM4Fq+wXTEgAGjMpK5Gkb92xeeluz1kDzNqtIyFYflu3oharUx/z3snPl255gVyK5
Dj31KyFAb1uSTDiIbRDampJRdyz5lwuy0n3i7VMEh04hszV8X/O1RoQ7QmB56u233FkfcqRsqrtJ
f2ujIxCTJHaWYVqtkLaz2Qo0mZAEFWWmFeDTuxDX9VTjtxkGKGoaFW5a1QQAwgUy4sok3lxP9MJO
UnnknBdbD13gEE8sKzF6PYLLGW73T70BGvdZhpoYxrD2TUMeLsV1lWYxZTFV1mlTYhVwghDi2RcI
diEPm0C2UWNazAg3Qn2tgp2WhuMA5rlfE32AjHnPllSqPb1Y2wlrjXFWrlmaGxr8uVEawR9BJf8T
Am/2HH472jvWyrZpKXqpv5fMq8+KUQfjKEWeNOgpKk12VR+MvDm5wXOmJX340S8kbQmT56R/K2t9
Cl4IS9QwDfTBluoqyjTH1bs424tkYeKsoTThvVNUbX2OQnirnV9QX8SNoJWtR/1DHwiEhEtJXpU/
kIRSSqYY47u2oCsrrdnk+QKJOjq0C/IllWD4myRX36mz+FZO+HoyIKCeWu6MSATfkGA0OYJiFlqd
XoU2UjW1WiyH+VzRenoE0wKI9iNEwKE+ukVIzs2dHa+WRZgy9K0DH6yayxg0Ur2j1PUgm/IB83/4
+yhlodnvRFszCPJ1kjKM7J01Q/rdDRz11SLdQky8FO0l6cVpX7ZpSmNydmKYM2/m7FY21mFbSv+K
hVmEwwBxZcUVS4Aa7lKAuFypa8iFWjDjsy/cLAjCGVs7CSIcHbfvdGiVisNa3ZZRejjLPaOAR2hT
f76H7ss4XCwNvy5snbMAIO4AXp+KIIC6huxoOAZnSsLvYoarQ28wEfwDWxlM6Yxe1DY5QFsPE5vT
R5SVAFcw6ffZ5+AOEtxGRof6WgC2O6Dv6oFXEFYk4mERWL7uB8xnqVPe40x51kw9VfrAj61mBDks
0c4SML+fkpch8f4NrYG0ppYeYotisioD9cIFe1xcVmo6aT3Cv2PkUPvfvrSNjPnTgMnticGFMLf+
JDQdJgukEe9qR8FJiMB3z4zH0P29Cy6sxa5YQ9CgwLy7MwIJqqw4PPvuM1l0X479LL/z6LwnzpxI
zMq5SRcRRSOjzyk6p9VdRF5vXdMxrA1QVuZsVcJL0DEcF/SKjt7AceGjPOsq7K1/SJp9RcwCnfuL
ifPgDbYWKrySnfockk6ez1f8UkukzgzQ8WggARkvw7jtFhwg78H/zyInNsdVWxmQe1blnRKWIRF4
0U633ty0sifVJveBLrxGTxXIcc6hVPCA1hHBEIFAh5mshc4LeYEoD2QjpbR7a9WZzT3wl+kUja23
faa3IDOwHLnMERBjBRSni4QLOrRG9zQTrN+6qW6YqZtLDvB6vx6YvvwL0RBevXhZmHqOdSIv42yr
mwjrkvR4EI7b7QnbqJB7QZ07/IDRzVhqwb48weX5bCL5K7CUMihfftnoTDHOGDHKnbL/13K3WjIB
+3wBn0PEATwz6H29yFOK7V8qVxZJzP+jPkRP/WuD7DB8KNxwJBqESgpNFrCDb2IUnwq2VWV0yu4M
naD3cTm0VguwAyX/Klg8iVNWpwAh2cA6x0pkgRrWMHjVlfLpnL6YkgM7EDHdjGHffXCy9WHmVYYo
2BG47ie/UtOe21ikpHN7VZWohaU3ePPgACJIXX0ivt73H6F0cobgOAPii7D+BEHPfqdBYk//dDgZ
jmdT5RdVtbVKHqOwlVgZQbs4lzJinwsbmR9lcISG1NNJKkJBwgO7lHJZqLRc+P1EGx5hMTRt4/Rv
RHSa5gWRASdsrVIQzfZYVlK4KOLAM75oW2KfGJayHRwLTP1UQWHCsV6lGxeIIDSfPTaxi/UM2AJd
HDEE3FHyJ34ZBMRyximppaB+wVl1N9eG6uqPX5iFDZkAhzS8LSyT5V/iPFtXx5gkiaHt0wYl9BCk
OXH76i9tKOgVE7kuaeTT/rAkK5bmsRxo7IX+B1HcjEZXZc5r+X3L8Wu+rgEwxeHusymAfo+k6X5S
JuyIgB3AN3qdm3oYPB83kIGCIAIxnUpVp3d8gZYrQB97JtknigK7VGaMT4MKurpLqigeUmEJ9Iqk
JhDSjgBO1i72jmmITy2RxTlEWsbGhXgklxw0f2OkdazTNlsXnuunfmOFO1YiIW8DgHKQ9il0zqrN
KCFfR3HVfDdGCDx8VP/gJyDW1+3g1btrfh7TZRiFpTpBBwcQfnzj69UZIsZEq9mXGxPme1DMmTDI
+50rJ7/X9GfXkXvUzIBfcfCDC43RKq8pqGzSLs383vKPLIreB1y5q86BP+/LmGVDD0v5fzvYpHhA
yypZNSdEGb0MEkH5g/f/DLG3kuD51y9jxhKOCyVBNF6aHZK6BsOQAAXFDw5ladP+sJsYJEHr7mrS
J+TCLj+EOP9wDjF10WypNtNGZ7/BeAGdWsdQF6Dyzp1xmQsZz2mZ05UrolL4cz9nHda8kOjQxLs2
dV8zSbFp2gEBbHK+o04SMYXXECag7WYlDo3cE5D9Ka1na1RQIVx9qtd+pZB4n0WH+ivfQiyj4Gel
T0dNr6lBEONS21FN2uRx9cKfS18cWSQ12trLrFt9h7xXrXvtfYTovjWqnCn6yn9rs+dYiMp/qsiW
/y/5prfwbIFQafp7l6QYM+aMVNVhYJOa0KoE0MUwHF4jRmuXl4aV9p0eINhXylcu9oaPrhnmtjxN
bJtls4B5ws2Jw2/KCtxXDy6MNC5knm6m55C00ROX4fj44rF5VQvJRw5qc/5av74STUImkjkOYI0C
r9lB1MIIvu2TBbZzUethaRKqF3+y1cO7MOZ2DfvNUo3CnkEmAy9pNZK4Pw3AMCViljriuCBpFH2j
huPLcHzofsMctGpgvDynVJQP4I1wBKVmCTPAeJp81kOaztJmZjX51Wn6SuoQwuKXEM/AIgcWy9vd
vfEVR5aSH06gX26DZ012XrnIfguy0/njOIu3U/vvCdGtLbKeEVR+fFiK3UWVq45xJQ7KQtW7g5ha
Cv1futwoBQzh001c7ekncKCemdxnO9lX7L3bBApQGdOIyNvqBrfsUnzqrmWjNeOyspp3wwJH7WAq
FH3NpMCVSmkPGAiT/EqPrq0YyhbHiT2S0naiP9vs6bS0SBKs729IWd25LCvfqjgaA+PE8hQ6P9is
oHWTZB8F6qp8cxwSPJi6OB9cESuoHzQEP9IlPE2TDtEEUYxVqInT1XSQU9O9gyUEilVSAqfqnsGj
8xXAFHaK5AH0lFUlMHSxsstirafwE8AueDsf/3siA8Ct/sE/0v1Ab1DikciK1a2xzLEfxSBNwV8r
dfbaHXL/3sMVWkz0JOQ1NaRyloTMtc9RfkWEDnFsnPVxHDSPLEC+4zy3r7Z1HdZaVhQmlrwCugfp
80LqBIUek3+CQAbdPkJRQ+wbOM05q8SIIs0AwN9NWbozJm7cvoa/ZR6E1/jl0fsJ/MH4M7njrp4b
q886IZ2+ZcCo5aNXbVzZtT5VusQdQNvBpNPnpHAzhxMOtR7vzKCnmsLNbxx8xI8mqTPRfcsieI0d
4VKT2f5GWC1toKGU7mhywONphE7C5dlDTDRZ6T8BhDLHXmXZYtlIntpq+W5/6QnMvJD6IktT52Cl
IE1VXId8XEicT2qXnYJEyzuPo+wPF9fHW5ZnRn3avAQqnug3hNt8J+HFvEdqiDZY2jqLuUwmSH0/
z3/0bCDXM5kOuLCBYKC6F4mFacazenP4F4mND4grxHQzC+Sh4I27TgTSXzERbQfJqSxOQ/a8J7+M
kGhE81/wRsUczWc6HJB1jRo/3CkZtISWB5dB6JgY+4Lqb7B4XWX4X8W0KjVRbzwQIvIk2F6+3JsN
/hD/gTOKAydZW7rbGHD5cIqVljI/k2KpY7WwvHUmPxp2pBbn12lYobR9tEyhtjp+/vULZ1/vTdc/
CJiaP1JW+/2f4xuV5Kd8vVFw3My/E2aWz2xbmJpM146YfvyOF0xJ+NQnlVzBZmpKdLnUbtCha144
ePcaHOtmEVIfevZrqTRFoiMDrFvYT96ZNdN4Jw3BqInRCtOqFIZSOvT7FIQ6xKpfh5C5e/qd43uU
xLYxZ8xP8Uyxyo1g+iVbMcapDk6dxVTFIv7uAeWNyw0X6qJbIGr/cFiOND/lyyOLsPcUq+jRYXts
04hjQxFXMlcNKO3h/5KaOGSqYc9tYdO4sY5TtKo9pg3NQCOh7GOrgiyPx2R4IXMDBs81jbEhIqrA
z1mX+ksP1W9W1tf1ndnf/naKglBDFArgW9vJvKZtzML/2VLsyAL6h2GGsBw8nOlHn0alaE7dP2Hu
L+7zDJb6f2LPJFYx01UFOM3AEyezYfpRK4WGkLNyCUP15hq4coZXkBFJSBqZRxFrh46cBQuV640A
zUPl9KPEFD/pLrnGAvriDnFuVpHWlffVZZwWNWIU77il2ylAh1vtraR52Tq8zGfzyn8/wf94oV3l
2M+vlbEiaqEERTUcTcqL5yIUdyp9Gb0RigBdRophqmyXcpqaqhLtGu5FZVDeKWasRlL9UIuTek5S
JX/R+mhZI4PRWT7r7/mcJDNXyPKHOboVWegTlNSsWqjCK5EdDGrb0Ckfy4M38CEl+X/eSU2CUCcq
65898RqqMhOR/hlugpIEjQP+HWFTcFOEY6NvSBFjmyElufhAmLbBL/Nl83We1ByMixY/zEZnyb+R
3WBtR5GVDIOo4HAHLq8mi3UAgFwAViCYBNU5O+2Rh8FjLYDgQbMKZWyn0/9O48N3CoX2yYvs7EIG
pnZ3PKFEoirMxgcjgr1AzEH5i9MPSTMQ07J+B+oPWa4MQWNf4ww46ML3EhcohmAfK1jP1I+0NOv+
26o17noPNqTrU88ACiFOlV4b2nW285KPdg9+hC/KWmqtr7+qcUGbLX++qFKenyq9fT+UslbbBynd
E0C/vTqwXq9FgdMTLe5OXDLUdsBZBKo73ENspc3PJU2w2LgOS1vmhvunKT3GhJgcFaAoSl0aLdH6
V7QyIpvgGY7rThkp8Ahf+213OskS8Wru3kW1ADZvSVGFUa//M9HLILJ+osJrkairI9K7D4osa2oN
OE6YIb6iAzeAn13sz7+3nWSS/JY5Deq/r/y6de29j++MOI8swZ69etghKmZBTLJ4IY0NUzcOaS5P
cTuQ8Luggr+dx8WjOImeargMD0puaj+DACu2fN1TDq+E0FQRPsVHBxFhZUp5IyFd6Ej5dXUlWvwI
n/CTgEzpQsgrhNqbHJGY5KtJnjafiIvtC2+GgZ+59XGG0QfsUEB6e+/7Dw08l5ZtmWozOSL17b+X
ch4WrhIhXiho9pSQMHHYzM3nffen2jvcyRKIqhNRilmTJ74KeJHC/Xr0urPFaWCyjKoceCjiGcuB
8WTlLXB89kNJvaYzL4Ecv1oQH6Zgg5BUV6hkIHNx4zMe7tjF7lQxoGFevHomZjX97DLYQMuau9D4
sMpYxsgAkvyjSUrEujB/jWEjwT++V1GgM40f3yCcZ1elrmTCpgmssrGXAF+5Rf2STcUnDNsayzIC
oXWw7rOCLN39hdoJyjVwIdHH8f6WJAx8cjXTRNdan4c9Qg5YIRr+1oQzpCUKktGF/tl78eCNAyX5
QD7Bvy8cuQXYiNuTqxZkiXbbPVCYYIanEsE4V3gN5LSAjgHV/y9A6hG75uXabKf8Egb4aNwE7TON
y5McvBEwGEnbuFhY5bbacSy332FLbPaxhvJ+OMrmfiAjXeuan/k3pdwF6QeEbtu8EQpC6PY4Lk+J
bWEZ41Mnx0on1OzxJtI4EbxuZjLok++cW/T4vcg+ksDjh1eDpFs0rcrz8mJwGphJ3iNnv3xiXTpz
xBXUGiKtTxbDH0Y/kgYtge+9C0Zi6d9c0L6MPo7PbGOAvDN+sXftKKx6RAtbFSHGzMDUgdXdUqtc
vwuUN9SDVmj+GhIJMgAfVSmRnv3dlkfuYfIHcLTuw0rWV/RsMdioe7BMKjwstdZhRZO2iEUD07UI
ia1vkSCeEIORV2hCTRu4jEyenWmUKCDCWEekdG1BxCqZpZBK6uVIMxfsudf34Rb0kpp7fiLyM1A3
Kn88hWK/790aUtAAdCzVP/4uVB31j+0MTYZ96KbI1qll2w3yukTidIHyVMrpuymBz8hS2n9T7or1
o/3Owz1ODiTcB+URL/Dx7q/4p52yg5VO/3+CfEjJV83/uifumxnESQU1w07cf1PDpGo0Dk1CifbC
PSKqKtEUuvVKE8I2e+T6cCzAwrMv7gk0JiFTD0wpdTUCaPihK0YfbPvs0TxJRZd2DxGbgnVyTY38
Mhhi7RijnOG8O5yCtXuH/v5sTxxZCSDAjmQ4xLBUngcXdUJdMa4l3cSqFYr39JPGzQ2w8eghLAEx
liVrfINCYjsIjjojumv88c7eBtImH0q4H6YsNVv2wVXJcx4rO60pfoLbVE3CVRLxSBVdfNSPFNCI
8QsFmrr4ETtNR1VoLfSG3lTLAOLWXyEH+Io6vEpTTHq4y3C4+aYqSBkK+T8BUNimK+NAomN2Owdp
M7lhRzZqSKY9HQxPiM5S+UNsU4MYvUhEiyNEiRKO1CvCndO8koJRRgKHJdb2MBMR9AVNfjov3nTN
LrZxCyIEp94vRiTEp1yw/h5oJSYewyNGSS1nFqDxsB2We5AcxmHj8NuENFWFDnhgEOuShuVW3/c9
5e5TLVY41QTE4rbElUMywt2xkbwu8yl/AmV7Ks3e9kz9eHW1VTZXQF6N0qxdrWbgy8xVh3cX//Td
DpA3sW4z0FSXfQjHZOOHOOMPY7g7C4DUdXEPfcGu0dVhlLwWmHfa5iy8ViOJRi1l6rPhcmtJga2D
HrB5KFyKcxlStgdDEj5ExCPt36EzKqRh7KLHOtfljQbW08rtRtWvCGHtBTdM8uLu/9Fkmwd33dCx
vLb9YyGtq/nhp4DDSVTVtpy0UKS0Rgm/GqwZHYupGHNbyb5wd8XbdPhlvl+xfyS0SA43cFhzLzaA
N7BpGxtNwD5eDscOqPxsYUJpm6A7KUCNZlMcE97zuBj/kv/wvAPrRgynALDFb8ZfK18CqUbKuU72
J72jM84GxAx/SHiKa9wqzarK/lWoDzLO27tg+gu56ow3lrX1JmaQeu89kDRtkIK2+NCbD3h5fYE8
ifQ8HTvSEitZbWeZv5BvMpgp2osRmCZzZMQvOeqCJap8mUaF3uyZp6OzjHZYWxt+Eomwa/t3/8tF
JC/RQxvMvqYZn+KUtdG4h22XgrrSJ1xE5qLXifQ5lhTCvFqDqXBJc4dPd37lyahmrxO73KT40j29
Xv+0wUJD8aaYp/AUFKoBNA+w0e5sT+q8ZGzMBv3rvszgnt3ZVcl1MB+Ccz2jCciRxB4G+jJXfrg9
6jBwUcPQq27auKUDxSkLJLm9JTMuenUD3SPYutmhaUXrs+pxI9HH4jZNpNnOmT+50kuP/ranolQs
MkZ8AAqVA7vy2NCImWeUdzmfmB/kEPAWfKNqimHi1YgiogVIj6J14DnkKJpqvkm9+Ui5Knst7MjJ
X3zNdQ1ssJ0Fo1mxbvi20TJPSBTaQKxIRvw0/6OPNTk/dcUr9mq3XsI+YM3LlZSgLGaeCX8b8wn+
/dELg9PZ1ZEsbIUqkxM5/kMftfgq0TbD0l9vsJs9LX2QKVsSZwuTibdE1uw6VRXAcVcXZoLi1V12
6xs0Wp9ZFpp2rj4sHZFX5pXd4TJux+T9QJtzwHFWV3chY1frasCjyWmUzjCxWr7DE4NF/q37hR3s
vN2VZT8eSLyPauIeIQAtISd04nX4EdCbL7VnEIJkkAd7j+BVplWqQrmyAB7b2Z6b9JmO7S4nBkEy
iaj/eRf6ZpoQg7AmMqfY8q/fyhAEhQav6i0jGrIG7tmlbsGBDXK4kjAjH6XyEluKLBEAX3Bdudz2
t2ppYOhMxZD/bEODJJoc0G70QHkSLK2aD8XLNSr0is67OBXKhGxzbFTRQiyx4hsWLH5SeOdvX54K
8AsxEzMbfBbon05xQihCyRhLmM9caqfMXd6/ef9bdqdWz5JqvRFPl4M+MOZd2JtcTegGnXJTOtMF
/EdMP2y0bh2LroNqVJWmN4oeBTsk7bYDMQpAE9xDOLBwZGACNC3LkC74mIWRj9NXwSBYYtdPKMXL
Y1G4UZ4KtwIEGdfNPao96h5OhCYJ4Jeyf9DxpX0DlWKxxaDtUJP9Ak+rYtaW4xMHSob81lsyo+rq
WEyZQKEEXDVtHxhE904FINTGeCrzQhp2ngy/zrk/e1zZCMP9b/U4BnlSLzLofsD1ekMPaPb1RUqj
ygDTdkFkv3Ci9tDUNec35XZRS628TvD8KOaxCd9vSzatODqi1XqA3IK4wrwtscBPcVe2kMODWpCe
MI0MJBLO3r0t1Q46482b+lETPerHIy4XKgvUIQkdxuq6009yRc+suIPEDRXWV1GDStswm7HErq8H
NzeyPil7H6fn7ECYeFi+5g2PNOq6U7oB6Sm7uZKw77xrauLc7BHphuyPTvgodwYWZO4As3NyX8fe
8vOp4eBIpjkrc7qEzZTi1fhsfCIUxKb4lrj0uku44m/23SDJK9/HNJUONzPW8PaZe7ErCG3JhWta
IlJKV9hdInOJpdOVoCDpVO2CPvlJPedVVkCE2x2eGjt97KM8rqmsbkwxOCR7f5Ln8kYBdpUUTkk6
wd2YbJ/VUy2OL/7y3ojQvhkMeI9d7I4pgmRI/G3xu/+quRCV/I3nuqPWd53VlPgw4FWVf0qk2lfp
uYgsRsRCNNJBA3epKn3+AidqPUCGLF319vDhervazddQDlFMUKV2Ym1xm6l/adQ9c/P3rnCFcy9m
CmLn1fVqURT9Zo4fsUE8q9ObkxhJzWh5NVUOu6ASEmPttKzIjFYkG/N9s4HVjKiDg+c02J0d9C+S
oJ0BRX/D3OZzSX0VYtrFavqZhz54rfzmEYhtybLlulfrj7dt1Lc3WTc5FAabktSDzV6lpuuWMwPf
W+F51zZNHxIUYKKQaJ6i/QGV40Kr0K6e/trbq+aGmAzlw6GGlxSE3z1qf3eRbgh1nuCG+1OA98JI
d6ZZQZfSrmzQ8YtL4fPKODFNf8mAzUZfqcquDb1Vdj0IHKUX4zE12GNvOLdTePMIfpjn8D6/WcRC
x3lp0GGSeFkri9JBtiOUUxOm0rLlV5N3lN4DFJqJjchsiEAMdOe+OqPtntl7HCkPB5yLRI72jR3h
GWDqxJiXMkMvK6qGFTU+wH2K0/WzoErA005ENX/vOxVAbIl/Fg3NhQEGO2yU2acOEdaZNK/0T2Za
kNvSq2Gj81pFw9WIQaNhuAoalXMQJGXek+0TRfmj0isPn/AZxUs1erThWA9/Jo9XSS2GYvxldgF5
Io5sUgjL4W8cnvOcAI74b8CPUqoAf8dlMuVkqJ3+0xYSWBTDGpUlxG8gIS+sXncIpNmaCaXJcn6E
tlrMlmt18wfCSo3rTgBLuJxjVgDoF8VgfoRNwS+l08VpunPD27pSjZxnM0HKMUaSoW6zw7UyBnyp
IKAavayjOo96/L33GL9Zu4Fdir2OuKkNO6PVbhXzxjUmamlDIPxFqcRrdRPzIPfISNX9M/iAOqPm
GDixdqM94WH8Sa5pNpSeF67Gzck/U1SsRjDMKWkGnj3UwqAKxCepM51dRSkZiM9pkXK7yeoiKxA/
EXIl3ddUXZ12LOQ9CC5o5DQb8ndCrroZ31/OppIwPjZfg4Q/nTB2jihy199sM1o8HQmo5wFoRxJU
y0gSRkwXhitFOnLaYfYcaExoGWGbU5ipYtzdMll594zh740hn8GFsxBeJIWqDEe7ubIG0pANBHup
u8JstjMxdXBxZooaRlTPtVUSH8tVvrG34a5mvztS1HD2594tS293F00hnIL+y4eTABPWmUk+0qJB
5rIGP7Xy/Skaxqu25IG92rdCikhDiRhiaNSXJWVj7QhxNRrZVl0ZFdGmdA4+Ndns4TRCKy8lh/dy
RoL8pjvnVVTe57SeQyjTo6yUvVr+Ggyn9V8Nq9JCK92W9NF2yBM1/MGKtvo41vVfDXF1YPzLKNbt
6FTxJX/Q7lTzuEpPcaWRwccRyriH0Kwr4VWB4bZ4on0aGSpRo6c+LR/QIxGiv+RIcVfFBwamvg9K
Tz1hNKeaFcSCHmfiXYRJeqRDj4BgTmJMz6M6xAyugOyKzDDvKB3F/DdpwaBJOgnTyGnmXmF3hN/C
JNsKVOhysR36QuA3TD8WUOs1eAHDI6KGch2YVpW35cEZokT2ShnCsb01O8zJXJZ8PREZS4+DGArD
oTrOZYLi4nJQ+0PrnS/FLiF51WbarwDWAMwvmD/pH07DhZ76p/GS/B+DKzowusaI8RO7Gnoi4gCv
MpJ4K/K61ATBeuUD25hXxFnpjZQZFoEvM7xNULkBbSGQWxeHAFnuJILvXZ1ATmM5FAAHIWf8AQCe
nLddpnscroAc+andXmRgJam5gSYJ2XV0ivcNUUbejIOV3zbeZMJNUt6F1+jPMjl7IhDTHKR2fssW
orT30SvzSSxKT2SPXIKqAmga2hbnaLpNguM15YjwYc+5nQ2khEGCF00og+X8lsq1uPTBSBhRKS1A
Ic4QWxZH7HKH976qTKBwl4WgGqHG7OsuIfcGjquekiBdBP17QTJ7fe4ujefdisVWJ+Gb0ZqGgl5s
qojWCVSYxApkmAfyackWYG60h28Nrd9wtcgdIjYDruq/rajBRK+hs9gk9lvvKFRK8eJPZU61uaFo
iUazidrVcJWZMiZ+P5P3+zadgnhmnIE9wsVF/TyrbI6QI+QJ4Zh2hZNdBekg4XM7cmw0Dh9hDIzS
Ispeads1DKDYqrIPXQaqkFJIicH6glfcKf9+HAjPZNs9FlXyw00sKXwvuR8v1ynr/WtKKJvXWEYk
XA2tfob9yAqQhsuLLLs34UZC5iJb179AZ837PyYSVOR/KOXUilOGDz1+tv8PCVhMQLrXrh2Zo+Ft
a22kKlRXCNsbEg0J9ZBXpwLq65YJ2XO2bxeprJPD4fOfGtf3nbPreqJJjK2HfuajBsrhD3ylybI6
lMkh4JcmvNqsLDmBaTO3TK3PVPxhIBL1QEvPZcxfol1oUTNbYvdURw+krjgprGiLyai0Ty8ZoKWx
60a555ww/zhSrHJJ4n8cmNvc05Hs+u2cFC88i6gWg0R3Dpf9iGqZgjeVoCHsNjl35LxT9iS4qfEB
ELoxcmqXq2jhlrZ2EdfJMdzj9ZjOcB40/7JgqyiBam2TzyqBxf4p6TKSWO7RFfK7rQP3ACQdDz56
x5dMP/6PhYPsmJGdFmNjdcBzbKYaMwKt8+P4oNEKR3iMfBGurRrB4jM4Y59B02CnmJ1EKEiH8Vpx
CYdGfUgg6QSf71GZpy/vpyg4r+B3AmS71+n4/IDvu68FR0ZtTql/IoZX2EvdJJprLxxrkrz4Hpc2
Y/ubB9j0mAeosQ6fgU6yGcmXk2or9Wik7Yaryit0lbeb7Ywh6l5mGTV3AATtaEp81SxrYWw1AfJI
jo6feuKIO9NnqsLhAK3Rhm6ZhdiRr4qz/h0qXmWG7/J02pKVR07cItawzEd0G+844gvTMJ8JJEud
6pWF52tEyF9J98sXpW2vea1NGI2YxYwArq3EaFi1o4EzyTzTsH2oWfhG1umg5i55fUX9dtUQAEEg
NXcnI4onIZso5Hcb2FSzpwTMwIR2/qDTbpH18rIbBuF+/HlZyCzw3hFvwez+3vjOWkRdKq+4uJkQ
/iOhmiYmnjmTM1zQMWbof/7JVe5JZDV52mUsVNMefQNbETdIT+/2RH8s845HiohR7xfCEXCrucxZ
m2vhkI9wy/HU43PayoBd7OIoYfLaqYBwfuILjtdzWcjXmbABVu0JQSO74uE+4S4XZqfuCAKySq9L
jMpbB9vKAHXuxObPkt7XdoTcmpAi+DYv+oRFaJUciQpERrI5Q4GcP6J6HCy1daybfsuzSqimqwjp
efoFUa4YYlnQqgF6pTMWR1o+lySEYY+cCv3pmkeWCJPfC8FpKA+njHScV5+LplwZbVhOG5hwOwYC
sLtY4sFFm5UIuwIknX1xYqT96zUjoOI1GhaqY1BU9vL01vZXwC/aC/EvWzfhrpYPJ+ncbhmt0fRs
TJhQU1oZsMsUIHYE1ylhwtqTQokA7UtdZiuCh0WTj4gK7+Gy5l+94ah3KKlrshQoFj1x2P7PYlnN
QkZtl5QMZbNF3ZPLOx0WGw8oOc0qQuSzW3N/Wb44fPiMN+bH4ogAIh19YkJ/vlsNpNLC+ebA/67U
VT79i2sISYibz2mg4BRwmGYqWqDqDzdljep5EUq4//AFSoZJtHRcMsqKv7MWPY364fjcLSNnC7bE
Re5IFqeLDmtpJHX5ZS/r4lOJl/nBh4HbraWjhdYLRxy/0cxOvlJlYj2Pl/XqxXkgKIH/1jRG4FDR
5MniWCNj939OiylKYTY04aSoNPXYSwIfi5yCjI1VFe/ObseEmm742TItV+k+p5PeZxwhcTck53bS
7FO1tJZd2kvsJgktB+2Am6BhdY/PYYiv4aXaKRU9t533d8TKX1yEcf0gADgZfDJYbzaAychZ8tQc
ppHBcJekq+TN7N6Dg8jcrscxd+LJE6IUwLbCOD0EXND4rh10okcOP2whqtts3BQjgzQPRucEDfPj
9ONQSwTa6dvbadnuOCojQvr3Ky/K2LOkWovCusAPXGtqABMh+Pgq/J4LMGj+S8hutyCRMf733x4Y
9WqR/f1aY1SFV5+CrEUDns2ggl+ZSKATqkUi55alORh8VjwUlALjv8NC+SzIrLBRetEzOlHLspCn
ETj8vlUILs/HkAP4NJVie8LpIiOJ7zKGiOuttyPRB6CHUrO8qg5wLAihM9Kq8lpBVRwgnmt5wyzj
JKbBnVkTMmRAn7ra4X+9JaIyA67E5ojXdytd8N8o404RIADmPMhBj1Jol4gZ2S0flL2DVed4Ak3N
qSJSPwt4cVSMwzl5r40W2QOthVlfgHzA3lircIgQcXRlnAMlFLCmo0eX0lmGqRocPSWH3qzAxaZH
RZ+YMm03hH2dEbDLZCIgg/3gPhbL1gk7dgAcznIMOiACDgmYv4I5D8xXP5pl8yL7juPxIoqW/lAw
r5DpMcidvJeZFAIJMCp6olKk4eKHx1+kJq3tJ8Y5aMAASDkgfpv6jECqFR4cguxf9GwLxrBLqGH7
Nvr5P4GY3hakoERGc0d99SxUDxMCe6aNukn0q7ZMPlTeYfDhFiNQf2zu6tUrYysMjoJ29DbQKO/l
/uc278ucWfL85RB/AJk0YEbwcXCF9SAN8xQ+0t9jYKI6jvVZ2X7TLHH5tpjLg1DN7yu8G3UEBZpZ
raJcc04UoOKFTGW9XUutpxWVpaXrhSAYNFL7AslAyYqAcCCYUZ7GmTKJZKjVb1LzW5y0PkUMtKdK
j8720ywDU+gk6jzBA27X8N1hgsYQQYtMEA4wvjCMAS8BwbzZn6GhrnoCFD9lM5K6M3i+q6o/o8Gv
aSiIsR/D9fhqmUEodtdwbphHjWI4D3HTY8tbN/C+vam36o8k/WC01WKQUQbAwIwwIL6AUe1Rn8X0
htqC8dUS9bwdxNSeTIfa/uqLvY4o1cwUmLgQOaQc9bSKHDxWSuS98JbtfrV+ZzNAIfz8SPVkVj7q
uBaYeEFXs9t/sGKNPOKgz9KdWeGnZ0B8sKPhOWv1PmMXfQOZrcV+ohk/9zBeWvIPT3Jl7/jDE48u
2LCHcFQ7bY52Xev1riF1ZD49lecjWzVi29sqFsmqUdADbEGAPOuQn9IYGKtZxwRnLsuwdjHgb4p4
X5BLvOcitK+tz3qeukPQ/C1dXIpkUvNiaN8G7wbUc7LfQABs2ZAJvZE6JkMXtsZg7lTDRsxqxBVW
eLVId00oqJGQKQNzNoDZP1pl0Mn5dqb7scpxCr9XRI0LlFco52S0aJbkQ5RTF9/QPrdnH+Lg9GGP
sTIsDwkTMjnTNtH15P+vHkaTWMvT+Jv/AZ1UNGr8buoGfWsb2qkyKf+cyHJdUtvtdhn9VYrYtbns
zaEl1IfnmIJmzhfLWOmFdgDSRsYve7//h+WLfwPYm1MIapHZrRwqUmRdpvcWb31UMqBpVXw/tMky
PKFg+2VoiHWVv8UADVsb09Rvx9bEhZCy7YKhGNJ6vUu1ytIPuZ07ZN4PA4BQzBcb3lZO+cWdOmpp
xQrHjv2AA0+QHU9IC6RQtvos2Sa8u3NGI98Q/LRp2msGGG4EDQApT5DxYyK6wNdPIge/ohMyI1pU
dIiiEs8+ZVZHyX+kno0ZGPRG7CTbA0v6CuAIQtoKDOAXZyLk2k5I02ofKVMtK+s34euhsqLX6oxe
jcFOGcWaVIpOroF+2h4TawXtw55fqcH4IfdQJMdKcdUOxHX/lPP8eIEEY/eQk7lnTQFUgUY0BFnq
LvSuKWhj+O3AjgmE/Rw8RGX8b2tQtrH+anRJEp2lTW0cbjBMcLzwKg4Ked618QdCTlnUc72GDvdH
JmVvOR/lDQ7aS7madq46syMFBgytKxos1xy4KvUbEubiT7llixiq8EIO9ZJti6YlyLzVCjVnBVfw
Tc6ev4+UJdPIqHmVdlW5JRpqKt0eJkXg3GJhp1MnVq2epfX5J15y6yHo4rylm0C3MGH7CCT+jloY
Riocxa25DC2FxKQFlAl9UxnaF6u15Cv3R54q0CnFfUaUOGx81XWPMS3//nIJC84ZyLunVM+5UGSz
2bfAgHjIz2/eZI0BkczeCUc7g13KnvHNa1w4SaQFVFbg8d8E8U8hFvvCipDLrxvmjfak4JJsSXyt
C8dCEYp2KWHIOHIB7iP5poU8BVdVesOT+qJg6ET3lPEDKzhjd+si+rT1yhiIj7mqTcL1Kn1xyujX
/9qyEMLLLDagSQRZqZrX867G50qJ2VRa0FrC3lmdijCXF9IVlfWykdcusn1PFe2uGqrirq1VYOE+
4yVudpB6UZzlVaZttJQjnx1hOJ/+gvVRPyXZiVCZ5nUvsR1mKEG7d+Y18c2wha+6kRkoWo4B0l4m
tqnnd8zoVkX8RQwQw6UHH1z28v/iEKh4+5aFns5LgTJH40Z+D45hMqd4iDDMQklqoWlM7SzrsPm4
TgPx8i1KVgC6ETyG/UxxRclVKMzBzyvaZRDg+aLu45iGSGCEIbGBW4w9niG5Y9vaqj6cNn1j5Yf7
1rM7X+mu77AdOIz7eLRKOKg2m+c9czwyM8N47fJd9hfalssGwJTcGwQxnL5HaNlPAUjzc3La5k/C
tvSZOZJdSMkd01UiOvgm+SbgH8Cj4UQSZRIcvB8900BVx1VESFaKMvaMLR49WvKsXD4qHSvI8ZuN
HG9YvYm/zJ/2dinEpYqHBGmeVGcDhFbDmryB0ADw5aboqf4DRSRAkUrK7IESRXWiZ1OxxiCosO36
d8Hi6NQYvYq0SJ0dPf8iY+bLPGTHyOfx7i0mjh0k5kBbj03PpLSHMwyb5OXR8RKjSu0MxBx8Dn/V
JJUI0tuQrggteRqAWZo3SImORGFGRhVmd5K93oYB7AN+y1gEXa1uenXmq3Kyf7EUZIU6B8KiX1Er
7fmgMyCYWlPIW8k7zISNHN2olZsjuso3CeYV8NbNor/eFFs6lfMI7Bp5KB2SjhViPS7F0+YadIGt
HkqUJDnsfmBEDPf9QBNyTVc2uZ9WQNQy+DT0Ni3M/1WzCRLM8O2CBgDBLKsTyl3NM+EstqNxRuqp
4BW7zt4kQsHJq2keLbOzmjGR1PeMrhLZwQErpLcVNEca11BIgNlvLRpi/9impMwPjTa4WR0MMo/H
gTDneZdqFfkH0EPnAsGJmzoW5zt1KnLGS9YY+nXnG6FsMvnfNCIEi3TMABZd5MIWVRFmWTvBQ+kC
Q55Nr1i7bYDWQ36VioC88oV00lMOEN41+l/PvoHE73aLctoJHoztKNzTHYT/NwIHKkBZPyiDH190
U5FHhvpH8vSj78F8K2XPs96SYIkULI2XaAjD5h0mAL7CYBBqo07AxZG860yNaRcRfGktPBTkgqJZ
gV8LFNvD/cHS5orCtaXDWGOXqsJZH2msQAJttpb2sn5unPcrYJIXSFSCIOYld683Lshl5Ncvypbd
ueHhCw9LFsJzZ3px7DZZ+7jTCENGhpp146B/bhxT7O0KjfVgoFu4rNHQQAJ7fMnj1QSs3pfUoMmZ
BmLXsR89c6AJKr5TVrg7Ev9iapPF/tLm24jMeM9HaLztVbGJGiA8SCfFlGhAGX15pC9U2B6t8SSV
eQAAK0gMr2gYtmSaMGNLuRubGot4wmEpvG+o/hrBlcKVt0EzZIxBqxEk3rLEANXiRpxak4lUAsHF
H7/cryB0ltWdAHY9axLDUgFslFG0FXAUptiVpTin/MjgFWAb6I35+WT6c4Lm7s5GwhnEd/yabFQY
b3p53OgyVnbDJzRgZzIByO3ydyAQKfIxJFAxF9n9hDSSdh+WjNepXL83ElA2F2/kvg1HQ4nCTsFg
g6kkIC4bm+wkqkFsg/ng4GQGlDXVFdoSWCB9kVTWU3alTZ/c8PdO3R5QoA3/5Q+41cCZv8rOeTD9
+J1ytNZJXXDEC8Xql6ZGq8ji5b4Em8dPGB624s4Njb8kwhqqKXb3Ojx1Rom4EBMc3ILq8KEz3jEW
Xsw5bDxLp9/N5/7GsIuzr1tX1qy2n2efNVat0ioYoHVYjz9fiY3UNtkqHuvMoOeEO8dIso5cUp+G
gFEMiw6T5npXwxRlO0V09kq+yJOacPQQU0gt9xLRFXB11ReVQMzU+CeGR9vARGY6Q4gvDY+MrvmO
2gMBWK31Cw062JJcFBRHGBWSckGRGjohy2veYiah5qZ4/qHP2e2joJ+ede7aOW70+JOpy5Zle88t
JdC8BaSkhVZPKjeWZiQpYnMIB3t4vpIwC/Hm/qqvtrD+TVNUBrDG2EurzvweHXWq7+Crr1wPyXl0
3GxslFw8AqE3JLSWW0vCYC/vlRmED09/VqImwamPmPhyyYxK9oGqaXUg2rHSlgSrJ0B551MEn5E1
guebBVMR4+52riJHOwQEdyUH8wIJCv9Tnb0yTnLStnYjpwpqd3YiPPHfhUngeKm73ABNck6HKTUV
ojgsto37YoMaGJAnhmhv886J1y7JOawhH4hRVzvYxGPQ0FjJnpI8lt5dYwpNOtgFfP2vOQIHW2dQ
2GvWXXqJa8idD7DDXZW8av8UB5Vj/ZURZAHE1qb9fQB3f1Pxe8I9bjcCSKi+so0d97HnFzhi480s
8fvTLoSEMqJ3fx3yRj9Y+9/HMaNkZ7aNPHnXXLMhpkqQb5vCXa21rHqXP0eNW63KPYbzitz2NAq/
a6bcssIZ2y+tREGqDWYIupRzo70xQSGj6Sc8fGqkqQy+ayBsnoEzePbxx78tziQL3w4pk9HH4cnF
piHBK/E9uQELwTqoXApmSqp7z8K1JiK5bWQoR4m7e+gXb5hUx/E0M/fxVaqCXMmZzdIXkQEBrr4c
sZpVYgDBvtRehxdCyJEJQ1riaGzYpmNsicij10Yg0sK/vI0DjQbKnLFsa18OxGt9h2L53BvNVOHK
2GWFlXIb3NWXygswHD6aAfy4SesVVjTbsinyXE021QHvaM4nsM+BidyIFA+nPEWDjuchQVP8C1Em
QBTez0uQC2jNMf1ohwSxCfNSVdBq1MwbrIymPXfSS66Brne7FkUmvTsi+I/BnQgBKyNwicKvl1I7
KPjz+sW4EBrrDmLBAkkrdrHJ3CoAeHfqbSYRoTtHoGvfG1aeIIlPwlSN1txEd7EZALxaPWG0O9IO
kJ0vhJ11T3Yd8nli6DYrFbvXVDt7XwJfcz6S/J4VKgTbro4fD6eP+BZVupUjNcdqKzIhz2HyeVWA
NV680yp9wlxyZslKTZBaNCseDLOI6F8KsyiR0F8p2a27gY4y9Nf84uhU5CF7CJLxE2ejT5PUS6r5
VHrF7ZtqW0Hxb6R+08WI50fJ90XaDY5j3qxW++wtlRx7M0Gh3/brxiokXmdb9983S1vy5pjh9KXh
EeVPFfwR+O1T5VUNCGYNLWXOvLAesq8WOHzrYXzWeUWaFvctDPBinxf40CdcaQ5NDqNwg0i7Vjy9
49WM7YpCH72kq/xAmG0zjdvhV9M5v3MyDZLoOKUdyWh2PZu/v6fHoLd/z4zvkDGFPE4Wci642tYe
5g4W2/fclKkYUUlaksedLAckXjENRF/bpjvN2TAOyXVHmBahIg6PbKQiEMSGTzJAjnHcH1buvoDL
lMBw84umChs9ZlyQWU/KEPBpXEW+R9RHp2GzueXXCv2Ovw/UrEMgFcT+/QHqBxhZVnLAO3GknCW1
rBA9aI3Z4X48YtPo271g4A4txHjxuS5XEYdt3NlcKV9CEnXO9TiFc0BxZpUio/kSciiWb4OiIpo1
4Qxv0nwyqXSj6k5696tk2RDws4R4j4lskwMB0I+h82NKR277uDiccHvuky1bD21nHviFXC1TGN8C
f91BUfSAUTSbuzHK7t50Ay6nGn5+/hpmcp8GY0qyGx0fFj1hB1yaTBSGXgDAztfUydRjqIWQxWT4
IGfgs+NOW940Isq7BF1DD2Uqk5d2AiqHNbjze4enUddoMy6ccPSQFJ07Zk1Mm24/yJdEHMhIE2BB
15EChgMujt3XtYGnJsFHsSK+rgG9RFS6TP3qa6A7Go9yg4BCVOWp21yk4VmuLxxdm0GHsHaRq7ir
IOu1oQdbOrWrkES+bjZfngLS9sk+duzJXsmZLRnqslwchLpVwvSN/YnSD2oT7TksxBytuv1TxosQ
fC8t9ZGdrcYTOrl/PjCansSxXsLokKIcr39AE7iYT+QloNivqpjhgVCXjQzX5iihxfomjmpAj+Ly
EaTrx6eIvI7XvELrNe4/E7samkMWw42WodhHhkn1aKEg08gOsI5c2/33QBpo7ziXIW6lBHqH9+ca
Y141RPFnUY7qu8MSOjIUpW+mjyNL68j0fXA1S8cioAx+IzV+yxDJLgWJza+s0dNlq+2YpXZ/IgvI
FhOO2fdt6bGw1VjGQqgHKUFE58SbVhNJ4RHyop8VAwRhqRjGoOyoF74EpIVPzbtLaOQLsYDiM1yc
7ezOT0ga3JcLmVIcG5cfaxSkeq24oaELqxh0zFuGalRmqtY13iTrbWHIxzJCPrJu5BmH/ncrPtz2
YyVt9E4AtHRguytCZKsw4FkEr6StkZcUquP4VONRNsp0D6Zjivj6IvbDb2h6jjz4cmHIF2FkCDNg
2htpHcR9JD5+QF328vQbe4nRDc4rrJM+5W8GVkSVxe3mhI7diVB4XFuGTrMVM4I45/c/6pnYsG0P
rxQmEVj13p1kN/lPpHYt0zTktSvPWxIQ4LLvNt1jTzGahqBaxswRlBw5wukRASpswqkTFJkTs23M
WXHJBGYooXUtLb2sMs/j2Se0VT5avYhlDWx/pxTB26MKinHv/UMkMUqWPNo9HgWezBUs+LC7P8Og
B51P1ZJTBIpKhw3uUAofoMzVaGJ8akvzvQgIXrj6lzbPNnP7hnOzBgV8P1qFINXaDnaD2cWh/aWm
HKH/59ef0Bgq0RlmfBqdXwKSMJ6xtPJGCj9AW/a21kxB1aJrQJBtR9S0JNnrLJPzM31aHv2mV7Bk
UWwpYIBZopW8oP+Fl9lwOvoaVyHLmzmAXSIBSAY+VTCq9Bf+1vmUrVxe2CL5Kuh5FrdeeIIVMDTF
xlOqYOwGOi1dUPyfeVMbg7rXW29wzb5QF9smeEbnvFAQ9t6lC+Sdc9OjbPyH00j9O+yxRYo88q0i
20sNQFnSCQ6/8acgsDCPZvmVP1lEh8ymBUmNVo1MADF3cgBiZ9LcL8NS3HpLPIG4LH1CF41G9e+R
ZFoLOnP1ee9sXcLo/ZGFzqxq+28O/1fguMDceEYH0ywuScIgR1jd/z8pfJuJYCTHkOzuhTr3gM4l
hwZUFBoHViGrqUFWnXPefja5CCAt6WfGTBsFJq9jH9ajlKDI6LSe0CbYhzHSbSaxMHUdzwsMZVWp
V6cK5aot0oJLtP3++ihyyyOgv4Hk9TzIKUAax+9JkCTsqAlf7Ys1iSZCSt5BfO24FvmJu3Fh/N1c
hiYbOFZKmnH/TCsHQX4gtAHQiswxkRpBe9l6G65zCKYKnB08hhDHIgzXg2z+wc9+8FRt2MNp6jDO
k2oXJOuZ4zv9+BCq/MVONCO1nSiVfMZwDemPAZXEmdUuEfpF1q+XEmn7pO85qgz/TRRI2O6o+jlI
SIawnrJzpdJDqNumsXJec0NYQUPU+k3l7ZSYRhoj9Voeo6Z3g+CI6WxT9YpTYrsjkQQwCaG4C0wS
Fb/GckjSwdCHQhIl2FpecV6PbFkcy/CAnf/dho92Mm1FyqILCv3Dyg3lvnVsJX2wfPh8/zVollI3
Pz7OfJ2fpjflaFboub+lNgYeIGLjfs+5tnmOApMgyjrsB606Wp8svYKrgPmz/4AnoZMSKH/RfOkv
I8xyYORGXKUbE9ILCgVtQ1tTp+km5Z6yzOm30TuAiMvL56d7WPdRkOJSRnFGZjKtYN+KTDsIjQKp
taEQNdUDIUYNFzehdPDl7yOnP8DA6KM/M5HpwMyDtI1UiS5b93UWHvFARvF0PfNRPgc1ZbPCt32L
zr9tN8bVnJ5FJMiX6Y01X62JBpRJ79kTubAmjL9/9PKyx8zyMjpOw1SltzFmpwpVfciYKu3NmNF9
uaQWG6XUCNnkYTl5BW6mxvz4g/IwwiFBGvk5UC9dJ9LzyjYdaC6Aojgu5tuwH7uFkaj29NkG5TS5
kvQQVVxHLBwO8nNlcK1qhRceJzpP9M7Kil1ycfNiLruLhaWpC4eWdnijaAPKZfjKLLtmwMlvP3T1
aR9pNmCrH+V+otgorDAbLNLKUiI6Lqe8kWvHUZra9KB2jMWma8/lCmqnlalqMwFxeGNjbYgsK2f5
iNNlg9OM8zDsdWCOPbQO2I764ZDGEKCbToZTpEWP6H0qlfDbpSK6gFkv3IQyG89g7VSdzzx5POZi
uzhUiZZ613DPCOUTQGSOLjuQ+FhI93pQgZ5PpPqkwr28Iwto2gttNd4BQ4yEa+nS5Cr110CR4++g
ZONo/LQ5dKUmGilmDy39fFyNpHUcUVachgOfRd1in/cg+AouXUQkgpDo8yd4KElzjdBjZ88atBMG
Q9s/1EfpCI+IIJeonuXOExCb3Bgv6ZcJF6ZW3xzpX/r39kuAFzZGxOeO09W5FU2wIknVkK/trp+W
dnLrkDBFAgr2DR5Hcvqx9Jof2M8hMo9IO0GmTcfMjqMjXws4a73MFyK3C/W8BJDUS44tAhNnoI19
/HlVkHxzZefzfTvnbuh3jvFSBB3/L1MRfL8dtFWozNCptAbdUf7/PtB90/J8BBMFIa4cqdTXdIcu
tH10Zz50woim3nYbsclXkrHsVCATOCCNpmP9d0FB3FiCGhovMOCL1oD0RMqolGNASyaLDdjWNaeR
oiSmcASyQnwWdkowKrqLiNrQ428xo/+ykpD0CeehH6xYQAnHCxA+NskyG1EFlhIPgEUYvS9XtM3P
rbK8nUo2WpmEjQWK1N9LfsofsgO1xaIeP2vSYqhktx0o8EFv/Uws8oHZmP54EiZn5FBw6aF4ap3U
kzZ9ijMcgaXlb9Gh2mdbuIJv6+2M5nagJ5KedDWBrrGUrmXpsbw7u0WeY/C5mZLYyHuXAwmLB2jZ
xT3NjZb6DAXnz/xMaKUC3Ki55H5ZnBJktnpZBR9WTbth3Ebrkn78I8Vjp0vB+58r++yN3Bd60KI6
mN+DJSQA0ApfNGkgWJfEgdl7JQjTNPHJbAyHR9sld5RcwTHtHr2FHf2ufdPOmOEIXBO8tInp7xig
u4LRBRDegGmlg98/1Lr55E5U726OUYZyLq3A/mbAI1pKu1tMZfhxBSBZTB34cXV/Olb/sDjHIGCB
Xdb6RvdU9jQrtolHCfb4wEeruTwFlGYMXKUXmD3ELVtpRwh/yuSWXt3OljAlclCKM0oFLn5aXHUQ
q3cYFZAAWKIgfDvxk0R2dNNwTk/GcHneVVI+eq5I8AlKZaBMbIj8zWUYD8zFk4vEoAuyPQhNm9Eb
HWG2L6B444lLxNGMEOr3FZNu+jtszhveUltpH3o08Lo6zc1T5e7l3h7GGEiAaddeXLhpQb7pDkxl
FKvxyu1/94EHKLI1GPZJgV7NlAP9zmHCOhV6+4B3XIzjXJthKOnTAM+oyRO0trk/qbRmEj6QQ9q1
WoqssudMUAiftAo7Fr8W7JHzzTR+9JiKUoZn/ewspvQggkTZNan1QCtSIMBfaJk72pAM1p5/7yoP
lyp05aHR8TTKZGEJ2WMUM/0Tv9prKJzz12FBXC73lRgg6hQLTHT13MJY8FquWrw5cFliax4hYnGr
jBhjNFowHs2uQrCv/1hlYcygbibK4B0Xulh9yWzcQKeFPBrXr+EV6H/ijdhSRRkpzmPj4NrIvZS4
irKNZ0zxmcWkBIBds49/sXXyAjdgXcI4A3NNVZSVRpR7z+0YfKPhVsxf3/Af6jz3/0+mqTJEWdBN
W89OxAbv0aM9IYemslaJ5ujCCrlsxjHaD/5Zf4XJmNI4okC6Plb7x2dk7Vq3tmn3zvgIG/DMTC39
nz7h/mdLM0NZ4Qt0Csc4kl/GJSwM48hEmLX9lDaVZYtRGBJAhqkk7xvGtCIy39wBCt5h9Pa58CxQ
iSaJDhdFpC3k/Wsc1lrGg7LXK5LJPfNPVsNtGC2nNh4G1I+WlKjQO/c+GQrZDKLK8tfmyPCVOFEs
fe14cL1Eyp8P7HVUHASX/J/VP+THWXI7K9mgaEtyevjLTG5EW5YaaLb01fXZ5Vnm+bneS7MswPmQ
MPPK3LnADb+nLHKKUs/AI7FIeX7N6Odv3DXtoSrIllXRIvOxGAZ1L/lfo9iXoLr0PrzhkPrYo7vj
9prKJjibt5k932M3UKvDdHMzg629v1xx2vRSbmYCifitGNaGcLUrpYmmyb4GAoW09ahJQ4DCsbR0
8Q2R40zwD+BGfngBVhKYtkX2ccXk/8adK060kmfJg0ahwNTIL2FVvziyTIvolaPv4ZmheCVr0aop
aAPLWgsAzFwg6GFK/T5Iu63M2OJYVVrb3v8t+mwGpTcsf6fvBgI3inMdY+2DU1hsojqURS43GRo8
boEfgvWuKub4K9fpXetm8E2Zl/72wOmRfQyMs5y0v669EfzdGKdn0niH9OKfu4rVOe9rr8woHWPP
NgjxXFJiPF5V9DB13S8eIAyqCrZBkHtkBOOpPRk6weCmJNVXQVIvwQODRkJKrchhMnpPl8vVBIUL
hEBWdLMTRpA9ee/V0bZ+LYlUU0AXdeO7a8RWHuJ5nl7s2e0xJVk89qT2ydth0wAFYIZs0B1Qar11
NXLpkKjgadxmYMj3bnoAX5RRGxlIwg2ZbQV6L8YnyH83J5llEM+d5F6u/auqUetkU0nt6+Le8hpz
Vdh79fUzgklCc+gFaFTyKdv+adQo2HVKS1CUyHAZS92jGSgd2uw22y7VHEqe17h3cbgWFGR1xtmL
yGLgLYbzkfO31Y5/z8n/Ai6cYVGgbZ51FQ8I2pXOtXp4QQHVnFXt48rEcvr28zQ0Bgi0SKDHP7XH
8oPoh080uNVEdqfJkWEbW3JLUcoRP+UG+VwwUY70ZDVvEbVxUf/4WBUzcW6mkMGLSz2wD9dFpM/B
BWrIErsZ+0aFzKfx8YjDpQAb4AfXQ3T5L1Y2QVSDCE+TJbaDZxOu+b0SaTDbNe6Atu6j9BIF0+uE
hb2BkCfO+Mdnjl6WPWkZx/yV78zsBK1Qil82Po3qpDXO2JpDwoLEkDxWI82m3LlBngtlQYdkKHBk
X1Ljp6rtEP2Wur25axWK7HetFyX4w+j8/Ic52v/PzLPfxmmZmpDkpprV4ZN4V2LvttvB57Ozdqnd
hkI4gxUFOjxgkH66seuHWmc24EtnSfvdF7Zt6zzrrq3yIwT3p50kP9sKTPJgIij0KMR2jMd6GNie
Hxg+lUqlkjUGZ7dc1a7jgJEx1sNx1Jcf3525g1d8R2PrjTnQNtS9gp5ttwZMSZxEEvk3KZintMfu
bmVDDLIiwUTYGRRaTdk7J+zpBHmYwtdTsOEpHiYITagNaMdXMOAAOfxO5x7OvxKlhImUFYEEeoyn
9NAy1lt6oMdVHE5KJQSfQ4+O+YFzIPMae3un2lH9jD2YKZl6iP3gJ8dDG1q3OAx+Rz3PYUcJErXa
ZYlLlUFc4+DwFWvnx8JRHK6PfQdmIq2nuOQgaSs3N3ozLDN91QJdntypBQWutsQ1z/xp0bhNHO2S
xbre6W4sjzc1iRbfO3Vp5dwFuGlWv+Y+8GX/JtVb7XfOZiD3/0vrw2+wNo2PhZ+eP2IG+lIJO6Wc
G7NrU1TrQcA0Tz2dVLylTsymD91wYbSUe6OcYB6oOTbyhO9MxB9h9CYIDDtaRDggwLJDC3RWkznA
QjutVOSqTyHKYaXVb319nfwue/1gz+m9wOGgqS4yYqEoUtxtuhbfUvZRHfTsuicCSZKAA268WhD7
dyAPzbln6uIEF4S1+IzpZs7SMQskOrzXsifjUNybrN0OhLPsjJBpWfm6tdpfGlEfhTvtWsMMt/Ur
wNAYDJVKc796YzsD7bSyc5rP9t5u7T4qSfOyVrFNdvWJRezJvA+tNhE2ONT98UREveAm+FhKwN3v
cNpgr4hi/X0f+FqjU6oqWQy6rbl7djuD2rZM4b51CiDjX7EYj9NxQ9GPFuReCdxsnYOggH5Xk35S
wgSKiHXGYL3zcO2JrP5bJZ2jnH3mGxeIGLPK8AtYLOYIaWkTmDD6O7NAV6UXlIpEaucwhU2zjAKP
rMciuc6TE/66eZbfoceNVQ8lCuiar0VVHHeEUETzq1WFE1tf9gM7Os3fBZr4+czplnwwEtjJsmV3
v5R8hZV/z5uYszVS+VN/IYNoZSWbyvD07Ja5pUX5o3cFUqjDn4YXYkeipZhAORZOZIzLdDkk1RG7
lmQni+HojiKd7VTfP8ItNsBFlAfWTWgCOXdqk2KRGiyBPFdIeF7XAXLu7s7zopvQzgDUFfx+i3u2
0i07w5Xq0VN4cQp6xGPZvXhdN6ZNTIR5b7RBEhlk7I+SF4oioiNHiyJ2zn3HYy5zQwrk4lxz9OjN
N3uVwyy7lQqx4mOL7jEj0AS+Psc/u6qts6DCln42CnAf9ePRd/awpCJrMwYsFgC8B+qzEQXGGjRJ
iz2a2xhdCvveKlEvJJ4CKFFiwwZLzrXByOuc0kx0NdEJcUezEM9tPeqxiimvBhLAhz2ZeMd/KUQx
B3jtOM/puKPHsoe76btyYVXxw5KQXQtRCbK6612xWcS7QGFpbxGVyRoIKe7Ps5PxIAL3CPETz75V
xRXM1AxBMnKJi6brJk6ciWBOjoP7AUdZkjOhdcNPp8FMN4ioiSTiB72/iPFzV4UkQzUHvtu1Y47j
9g2mri4XA48Wf6vFru/HSdv44eK2zRfytXmer8yFYvBlAaU9qdWH0q7fEdRzM3+Mzs0snph+0Gbd
uE2E/jk2MZKnCc0nhraHexx9Y7OPBoJ0l3FlDsMofKdGBi3Tlhihnqs2oYOl1Q5emKHTT3siQHg4
vkXp4lPfZl+gyFuaPO4Pqm5t6lET67yhSI+rYQP/1VxMKLGwzGl81AeCgVaQ9yAgp8B3hyUNkO7q
7W0wYhTotMtWNS93tYwbjk8xODMJ23ZDj7kS3pZpbvAy7Pi8t1S8VjZmH+pnxrJWAXQ0wFBIvbOB
hxG1Tu3jIYooPy85NPMJxz8zcy8BDD/hCJxtBYhcnUlVufh/oGvgvWbNizBYbeud3gqZHyFxG51p
POX8iAe+y7RO1qWsAo3bgWCHLUd2p1E03/6JMeUvINBfivhce63vmlQiR6OruqscpfU8rA7YwCGA
Fp/PMpQ7YiZ0u6ZZn1IQ9/DlbxeZvpM+FeViIEP+MdlAc69KSnF3IhMIzvtaO9LOPrRJlUfSJn7j
BbOv0EypvXLy3oXtUWHpES3Cqq953asCClj+S9qlcGm+wb6SoK1nHQ7jEubdsSW0O25JsgAe6wIt
bZo7zLY5D9ftCeDpYLoSTAj1RoekzGvEJbxTp6j3XwggfUs/y7kJgOm4fdnnxmfJof+tuUfFQS1O
ut+/IdBQUy3mj1VExr84q1RncFNsUcDIyssf2p6Rb68NhJkp1lslIpPbZjQ21TuufEPUDQAjr9eV
QXymbjfB+ktHgWPzAcbnG8g+I2jX9Ar0ZZIQET1PeHtm2aFsYiYZESAa/8RkC4BxO1htL482Ggti
aTXr7KDO07uWiavZNKaVukd+4DJWn5WQS0+sXAN4/YrdtcCL5l0LvgqCMGiqp0eQYcQhT5y1k0KV
uZ/ymxp7sJUy+oFEXW6kCG5l2a6Jini3UZmsn+mrPlREZ0DBjjIlkuUDSYKCBHvz/G/gB4vAxjoq
5DwhExsdiXZjdghYh5Gm3X6+CdfdXcH7AzBU+ceRGfLEpbgfJxnmXXgeEQtQZapZJWgtLzcTAbcl
7iK/ul/G5II6ABG7ZAvcSL5eDDy7EsR4SjfFJatIymagwyId5OpofHkw0MqLcBQGw8xupTD8Koo3
Jvreoq+TaqLEnC4LTVQEmcxtiwJT6Udt8hpb4voQHCJxj1qs5/QlOteWNiAFh38Bw5zAwOQJeveo
sDpsWWbUoiPxHQxwydJKYbxQeUny4fBdin8m5VuyN/ITgAmAwIFT29CkaCSe9A7+y+IZqt4CQZNM
fEYxm+cncjvqsBHenLoM2jE74ZCsTIolS1beIdYjzHTap3VN0BEfPYo3gNvTv04ncNHOXrD89MIc
nj218BRdWrcg0/f+fp3irMMsBr+QMb7SmQHOdSi8y3fsixRmq1yddYHRrFW+1XopZdktJpZTlUnY
X+CO7VH6ycGzHuraoldAHwS2uosFF3HVb6hRwiJQT5w2r+cQR2aJY27X7a/w0xRlLafbcKkvJRyG
2fmWDcJHmj5RjwtkvqFcM4+H76vrNDuW1d78AxyZwzMnRx4GSKeta1507ws8VZEO4AqTm8GXLr0X
tP3pQmBiJWOm8l135tdtaO7aNfY49BdNnzLJgs76oFSAythnUQhdQS5lTD5DcMwIHWlrKqgG7KnC
oznWTByo43twlTemtFFx7j/klxsVp+SjX+3pRB4Hx+SD3GgmyQTp+XXiuEwT14qdG8nT6/77+aXj
1VpBFll4j3oDpLrt9lSF4qC0bdKKl781Muzr9kiOCkWqbsSNA59ugPKO6Kmo6ZcG0+H/fVbXILGQ
1D8+UipfPJEn3ZY+x1hyt8TpZh/nPxycdoN4ZO89PN1Vd3gsP0rj3LWpwtE0FkgfkYWBf0jg/EPn
Au9WNjR6GxKIqAT8Dg32qWlO8I1QvpeKBSmD9Qe+X+qQx8njmkYngG1x2gyDfuLGm/rhUBlsea9H
dD/UmabNrfX2lJWr6ZVYCrVoIRwzuQaZ4PxUvbBpKPwOvwVvCSqDK2rwtQoB5aniLhiVQrMEC093
f6DVi1NUfX4p5ou2cNmPIW5TDPUYZBcnC29RzbVxZI3ag/+MDJHLJNL0rpYJMbITGqcsgnJCrIz0
oyDQMpq+GlyBXXbM06g+zYNdeoWdtKG5q1iKJT8Q0b3uGxyVe2wVQINB0Q3wqZ7nrvHk3hu4wvkP
mM4cqZ3fB+AvJ2ILtnaToAgQoGhiflswy0zuRLT8+SNe3onk9pkCYGanUXlrLplSp16fmQ3YrY/9
79hr9i+jsUtzh7YTWcoEka4/XjrHIvZ2pAqKsLKoJB8TXLRUdp6gdpMcWMn2xaSSYZPf7qJMQGA8
SrO7rlxx1u0ET84VhpdaaXsYvQFU7gN/BlCg/y2/Jx4L/sMW3EOgoi6rIOyxhS5kiAX+NwBsIDcR
x7vjWtv00EoSKVDRH/tCc/Zz8JRFDVFFzlSWSfxMZNLxENUtVXpc5nw0R4x6ttheyzg0mukxTV48
bmgEgApbqGkytKj7jj8uHI+PHs6etLpTzKv1ep+xCRXtKyG9YgJorC7f/8/13chznJHI8ESkknux
uFeZMBSaB0Zu0lwefnBEkLH6npIeCLm0xMXOGlrAUBfVpYaLMNLkxKz8tp3CFP7JeVaP1kKN7NFb
ZLc9fbukwYdCW0kbZbmuQoVbkdNlMEIgMTn12Xz2pBYG0ZwKvxhu6O+Msa8jhvLulsuPI4Y9oxrF
GVfkJvMoMbx0m+IhxjaCEddCz68v+VgLlbqbhlK7eIlb/rPF6stu36fbRyh348YqAPB6gmVv9m2e
uw0s82GISCjrhSKDn5qknKbpsXKuyhkdZW5FnpW2J6/xL19KCMSTQ9vovuNWTvlcUrproy1fvVnX
msK/LjVhbZ4xPrmtCS262pVm+zDuT3RMSO3BAUvFvGWNcukKKLpvTcGw8zy6Ys+rikn5mPoyou48
o+AxypP757iaUbef1tirTRb4cUSRUNu4lzyaUCKPgNfO5L7xtdl3YhCzJweHUaVpDne2UIb4GGZ9
MtC6GAD2/HEWrNpZ6bGc83geoPPjbxTBFZDAA3EPESzsb01NSwHb/9KgnvoOQDdaMraBdqK5zOgD
tRQIwDaHKNOaoKtdlxiWXJ3k2AGx2w9MaJ7BL0Ka//XYqYHEqavuAv3nAv7dfNfynQbJK8ptJk3R
y9Vzx1MiMywtF0ogocqlP32+Z7yge//x4XAeKGeN11Az9dqNZIrywXSBU1OuOGgNUkw/3t56vsgU
mN8GQZ5OkVahRgLWlElf+Vvl/FSo447tosyjDLYyp5EQsYvlMYz5jvkOBVqRieJp+OWjovKSj4pv
ADivteTrk4Hfh7sg0yxk4IdjycveY9uT8aOGCpxtFNQ6e78IV0+UmJ67aquAmaMXES/y8Jo4H3U2
DilDWZWnVLjuQyHwIlMya9izMxFgfpe3utt51k2FxRJyi3ANLy6/oWSvufDpHZa6a9B2BqxVgbpD
x8AJ57IHsGsOxAx6rBbe/XZimV0XxbzvPH+018KEYiUEH6bEvHbtp4wl24tZkpVu3k9OnNMoLeNq
FvSH7Wp2U6pp53w7SycdmVLoCS9iqJKy2+oEgeKC76s71WK7JYZtp5CPUyAkvhvbUFdWQupZK8xL
sGOURzkZULroVxdI4UjCMvyrO0xJcSYzIjn6sGhY7U8MGbtlTdA1rbRcbSuljQWPZQCa4VjlHDun
BZRPVz1/Zb+u7s9hKsvqAoMopR9aGXSbPAo3EICWwQGaGf4zk9JZc1d1rzibXmGput8ZGe3XEWg/
odFCHqTcQlvEd8qUWbSdnUncwxSpCqTGnmZiustXsQd3nDOhmAvATtRCaKUw2mUpXcEIjQ0e+YkN
ArIJ2vu6JXFFd2yZe6Jx5C45M04SDSmUOmn9gHDmgnlNkALpT3J+R1NxsnjwSkvRa5sNcnKcrkNN
rrJObmHtpHnVjo0bZm5F9uA/woP+3RCR7uCjP6TYtighbt5IKLc8okrAW1WHXutdXwS0i9l+FuSw
0jaZLp/nQxZiFqMSnTaWLCYWtlKW3JWmGTdLvKEK8UMVhCqAbk6rtXpFPLdo7jlVD26/ANflZNX5
kIcG4760/1w9KK+zl58QUdPhQHdKknnE1YAwhqIGH+DiXZHV5of/pzr8ttcEjIDwgLGpA0pGcz6Y
EOBSQqW84gZ68AbDIbn0ZT0u7o7w9mhwxAlIFsNQv/AUqYCE3twTH3D4o3TymXSf3RZZYQlCakc5
lq3Ii3n/cyr2WL0tXxJ9HKcTk8MHOoFXRxwMxDDzm50ltL8fSzqW3bFRHo1Ep1AO7oS/NJNuPr5Y
Magoy195xPnpRxGL1tD1DrxrVlfSZeky/8Qc7T1nPmCya81aDMeGT73OPp7zQDbe5pW4KujuwigN
pPG/IprxpdNzeTJ4+a4JzG23dEiMbeOF/xwz+1/ZTPpUKvgVuT0cCjFqWr7lp8LYqHXd9tLVcmOP
yBeRZQjN0Ix8OMzOIZXa+fcwnw5trjN1Wns3ECuYUxN6Q0QMKhZelouhvLDsdC7Wo20JNOJFO3Qg
uatx5iT7rPw/HIBI2M9PN32ZOI4P4T4Xfv5AOQ8sMeR3pGgK/sk67gEZR5jwng0c9MYp1ikITApk
G73tDVOB4+qi6PwqsXEEBzEucSIrR04XG3YqV5lUZWMgWyMGOaDzlNJ95KyYrT9jBn/TLoPgfSmV
CraBdkNKNtXmMyKPxTFXaudX4uP3R0HuLqQL8bww+LV/li8DzdNrNfsuZyAnqZ6fgI2Rhvz3y0VK
YmU0hXjHzEUd9vVIKJNz6WBODHF3GEhKC8PGQe665gcpCOei1GktWGfiPdyT6ezTxyF0EpSKGQFd
N+jMKPXb1xZYOdTQT/loIg0nOfLnyJZlj5fSe3/KI4otfs5EKaablh1cZwJG5LYqMuLp5tJ1OHgV
Ri42K3w8pLKt17gk+dUMbizu3IkHHN809DQjzrtPk7EsL8q9epjBPw0j3N+o9zw8lovExC79+d+t
n6vZTKSrgybVEYrXOE+ZlGslvb61ho40jtsTSzJ8gV7WeChPqySTDw2mq6NtrYy4SEdbPt5XlMw5
V0efvaAsrZ5hy2auI3dzIrxTNgtA6NtGtJOUECwJcRkVpY6XSCX5n3uUrJWzHtrAqtyONahamGbN
W9+J0EjIo1VIYPJXH/+Zcn+HNXK44IvB7WYoCFADFjPIN0LlZdBAk9mNqav6sQlW7Xje3rIr9nwB
RMO7DJGgf9Ltdr2U+lmtMB+HVCwy72zWPvoBhYVeYHYFbcMqOu34c4sOyqrSnA7nr53WlOgidIYk
LJ40HoTPODuuzzp3J18MpM9t7iKJEGzggo0huLM2yrc5c7V7ncpjNcEO16jtW/knVVYk5NaCuxnk
8SZEs7/3E9zsIS80xkDAtLLbn3qDCfANADCkbNxxJtKKqNZCY1dJ2XO7k40QaTOW8VGD6KIgOq/A
3LcJqd9bkfVJFIAx4JpYfNnN33B0KcYtsQdZoi2CO/6U3Mf+xLecOwBT7PCEXijOHUDvl7FCPiZp
dAmVQ6XURrrapER5fKHHwaOYWpGd+pnx4xNQ/ljVyXhFmmIqvjvDJbbDIFJ0BeYjBMlyCcJrfFrh
Tz2ox51Xhj/TUAJo5rnS/4VD1GE9cmfGz8tfqhwRKVckrIkQldyF+Hz8asCseglke2iCbEfmzOvd
CGJT7a6BQ438xcj4GaEfhUg5TDBxyHjRc7UhEifzZGX9SgjBzI8dX6CKQXHAUbqATqNs6fQ9s0aT
UQCmBWDDbY20hGJu9PvzlW7a3fQ71XqG+g/DZTlfRJ+VBRXlSYHY6Uo6xv/9qcOg7BRMtAzAn2E3
o53/RYp37orKMm0YIsZwtylYO8VnbIae1uLLYD45PhZDW6rcTlf/O2VGTx8H+is0HwtFM6ODRpS1
wAwtNs0a8XSk4dx5k4PtGWIguo1NXBtZ2msfa+2+j+9I0DJ1Fmeav3t1gNedIrfiiSamVU8EmfLV
Y23iwr4rfUwjRiywQJU78JpwHejxEaUbmB3snfcW115Z92ANzx9ifw/hKZMfm6UzszdRsCHGFJwl
84zumsGZJrWO2UcsXqgtMlMuLzM5r58OZpCBiu4pzh38Y+DJkHi4ZmV1jN+PWPo2ptas8bSilWfG
FLOaqil2/onBBiKJ6bUJ7XqWgWtSINmFi8+GnYguflkzAlsgIq0RjAgDnJ0CCvcpo0coEsvluSD7
srM4vYM/soqy59D1PtQ/BdFhowFXPld9FkjIdFOX0svXbL6thGshfPmaqC23ohEmdiXjEGqnS2PV
tWXx6z/mH4gg+K2hoUv0GAyQADdCJrFZEU+mcvnVACnzDh7iH1m+nqWoCyLat2KHy4qWhi9Av4pR
ApX/1MC5gJXrdameZ0AioAKL47usB92yc07imqRPG2mSojKUdmE7uYtKzWNc5iUfo2m4+C6AuEsp
h78dR+wst2mQfVtKEb4uH3qzLjh4rfkRSMHaodBRMUzbaKMYPSxhDk3kpORZv8cR5KLnodkbvQtF
bxjYS01t4v7i2Z3f85ddLaUWO27JOQjSKkRrbREd87qH1YWc7pIvY7QgZu1UkMB8eO4jsdmstfEh
fsXbqu8JoEfoIfLrMo4tmVA7BytX3GstRG4Yqgchs83bvAJdbdrMQxR+Me9NCYjBYULASns6jNYJ
rw7fFQBwDR5ejmuAjXWWi2cPeqpUmp7dhiqIsceVkkMLObHLC11LSScZptKZuvkQrx4C9t4/pxHX
Dj7TFq/SAtMkyDXAdHctwNzjRr2M7pGWBOv9QyzXmcw7a/p2R8suQlV4DFijfIbQDxXbUcLykzSi
7dvr+6rrWThaRnEBkRnEuWnP9xo2Hmpk6Uu5/jQuCOQ6/wEZBuIqntsBMtM7wXO+9q7wUhfPU5KQ
YHXeJGK6PcRd8eHzYIlxJH7rhNUTwRJ43BZ0hZtwloTg3b71+zqS4t4S2G/1qf+KvZXF41Wc+20q
TerSk2tmXPySuwAwhkOUhuy4EZ+3clH4zlR1kUE+GgCkKo++rvl/CaR68Miye3W9rOegNq9Hfp2R
soTy0ea0Huq0Zt3/pmujt5eB0gc1OcLx8gFaaGQtFdEOe0NJAxnCEfClkJ5Pzkc9j+YOBCWXKtEe
idE1yoLlbsB8Q7nEkX8Al1QYctbuHOEhr9yQCK5Px4tKrHsKd2Rb5Zg4aJiB7KWtjpxHTuLXHMHO
xXVuP/7T7VuuxZP+hNVwFLAPZACazdZ7eFGrdq9u1yy7PY2sFdx0aBx9Pj509Eo3byCaOnX6sQc5
fiSvtEsIuXmuAqLHDZE4iDF9R+IxcIBlbO+VN6G61OZJHu2k3JunqItDC1um4QeftgpA6yLML3iC
L3qxvSns/MPVwpunmCR0ks3lwvTHPLahI5xCJpWklFY0QvlqpAwR7rwYzZDTY70M/okbqKl3+H82
AK9mJ2S8b6Gq4qYkWduBUwkiquUkeZeA+x/n241F24gD9b6nMSD1jf5fzF2FC88oI/uHAzzW6DuS
8nIEVu2wLYCMyz7oEQi7sH1ovKFC1GQaJyG/vF0JxfC3Q3AkbkSGuUCfqi1HlsJTcNKG89EuzetM
3BjGuKKdbLpmuYiOzoqSt4w+L1+c+CozpVAuzQSl2aWyZsXQEiLNToKafWLIl4C9WvFUBWwBuYfn
IOsktsBbM9nO4dzSpc0LZLoL3jTJ83M+Fub4iF4cCp5bDX1HfrCF9/2cUkkoljzrFpnjRzlRIq/x
dROa80uO8cEGqNA5iRvM5e30Ltj5GhZ7otX+W+YDXhEFlpQVUyCWM2peG+HIItX/pYVkeYxR27Db
mtdMVXyvkDQYqf9yZfOq13WJaD77ptPLlGUFlf37BtiDWv5Y00BF3aSStEv/7sys+LVoU+OuOrIc
oQyEdcK2W8QxDAPkzaWWQ6rHd/w4zC1KdAfCuNv8m8bfESBlxP1p9F4gMHkmKEJqseqNC+nB8Pwk
9ZGz0Q+cq8pbxErWp5j4WvccMKOuCMlwzAweRmI3EKBmc8bihYRDeHhaVUQoeh8m4fmG8zSbZ8zj
E5yPRyUo5+Qtxbk43KcYGnlchB0/mQkg9jPG05wlfd8TI0lIblG0D+q4Gd8gRQ0dfzTuc9yBr9cx
eejkrKQaQ6mftOWLOaFKsTyUzEj3ffXDlmtiiW6XjW/dSPAk2fkS3BX+qauCALK8jix+1Si+tOz5
in4zsYVISUiztf+2I57D7WhLcICSnyY74scWtHltK3J2YyrPuPYTTpF8CsHTBrVcJOTsnvVY59MK
wJCwunD62Ps8lEaL4ISukW6luouEokdbOZVpezlNa791FQkBMKa07FPw+X7e1ENs4gRfp99qnR7y
c9yQgBlHMI6msgH1QZtSAWr9OIvVrL732/srWMvcUtAuoAM9/oZ/Vh1NqJPOdRtAyqx8ZS76/VNP
7R9RZ96AWkZSKHscfe7h/uIZAoGQItuZQS4sEy3q8lQdkWmpcseN19LdeS0rgw3pyeKUEhQasMJ2
LXxJK742kiDcvumDeBIPMWhv73kDijefITO5202fqZ/hPG3w2yZs7CQ5HL1YtUG5ncPF50RinUT7
pjHdl6pn7PDNkzOtQW2Dz3aMXkmejhp046GrrezS1geP48IX/d+khoe9eq0bgtfdDYlzGCjyRVmC
nvF3PB6AJud7GH2MovWxAwyxE4Wp6Yo5dnUOfFCAHt0yt7UZtbaxUgI17aTBh/WXE61U55Hzir2P
fg0Si/5gwJRk3c/VD7toIB4vU5dtB4Ph0cpPktKMURgZ3CeE+CjHx/HQR+Mor2B4xttGcjKppZ+T
iadZWkL76nSQUy3P/D4eTXpaeRKYXTadcErZZYCXpTp2s0PdqgJoXZjT4v8CAMugUa45Pf/bDiNl
c6b+57RaeA60bb+nU3HJyJuF0GaJFpcnKkKkXV2E5XyLo7HVbtpUv49T/jZlvZLvFg0w2BN0Fh4C
laaX1s5QRJjUPjkIQhIRRE1dOv+36tMmhW1v2jRG+9Flit4gkxmXEWis/QT47CM+ZXwGTUxdsp5w
S4WCSMhVfQCWbqX/qs5XoHdH9N1yV61RbY54NIDfoJpY4o4lNWmuycXmOhNviY676pB2tDxbX7ZY
IVfnho6UW/DJ0IdKLDwQERDXm/Ev8jY21p9GQReg0OBGRQnPjeHAEbw9dhqsIVkrdUJYB9QIeXVD
dcD7GkQPO6Erbw6utzULxAKsozG5TH64lKZDAYCoal/pN14N0YmrsR/sdhLXjjGsRtEyvEaldoKR
sr6+MfKD/6ozuxu8hjyjL7HCOhroKefzS0c8RYdBcf/ZFDGf4CzMzd1S+GRFcsI+5RRXqh1i92JH
EfqgbrOcGbAYdTO/hlnEBty+gl6oHX+IUbD5uCjLWYtF7oyL+KLM56esdovUSkY1s+ZNDmwkEIKQ
SlA1rz5E+WmL69D4qPC2zhm0I5Riq4V6X7oNUGb6z1DwXrzja9XIHBpSfR6DN48lWWyJ6dF2pSgD
u0usI0IRYIZE5WGNN0QFy3c/hFPgFmHWNJ2ApzL0+c2HJCIJc+T3jPNwtKXa6Ys+qyor32uqztYb
c2ppu2afpmmkxQ9mQID3bSC/dZiWvt/2PWHC3KlpurrpUNm1ftqP5y0mNLn+6OG4a5NRvkcTupK4
YitM55ZoY3exX+sKr/ckRl5XDIjdqEW4mnh7UnXCdIH3yNucqF18ZmJucYWYAzBVz8xiBr8sZMNY
3CroLi0vZvBYY58AiufIWFjRQDsOBwAGlN7Y/68rPCRe0/HsSCkMbjOmLA6tKeoPHjRtt9sVTAYD
S4rCHR3l+41Ard6yhvWpayKzA++h9K2FIhRP0YKmXBy9ngHzWnSAqP83YrNA5DJjl0CPT9c8XdRp
o9rvpytdOKUF7UHZeILo0EYHe65V7sEEtN4NbNijTdYenmUajykWvDBDpmq1EupyJTy4VSBJ9puy
7wwuLHPVuanAlzAHE8RqMivknBP6idS1wFsYHFjcu0jbAdF5bR7+orh8yYRZ5CCddOcqQd+ujFfN
3Ze3tq2+jLg5m30qFc81Z5OkGmxwNjhbqr/VD4IMLfHPIn2Pa9t8lh0QcRQZLjkRCUBDIZ86fpyn
yWhKndHUCQ5gBHVOFAaTq6lZgrUxVHUjYLBE15v/aZJEAkPfzKz6yS+ZLf929VcyY4xIKURZ8+7R
FO82zzPwyW1SIqCTWVtKytNw7c8UuFEtHaCrf2HsEvYwhnLFG+NALcW1lGYKcH3jN7SAyuWv95Q4
wQ+61vm/69jHQwcPEX6XbY/eH/BTbFRrN6nhS0/K2HuB6YsEmPSlO67VstO00F3VqnsSiQQngaqR
MtQucG9fmXRbC+bWg9JD+TsT1X7twT7ADd7ktpc8QmY0sGXLb/TUAnYQxCzvkz8aTnKQBwzWcB78
7DERaXabtwz6kdjcTk1gij6xUtvfYDc+IXyW9SN+vXFycWyVrR6ezReOnxeukf6H6Xdp9+6Asov7
cOUHaeYgThhq8joqK+Fx1RUOtuZEHTYK83Q/YHlacppyEze10kuxrP1CLf6ilUv/YtO0IINy56HD
gJ9S92t4S43N5mOGL85Nlsaf34rbxIh1N6GPtgo+8AHhUFZDIiF1VYb6j8wiK1HYZ6NevcXbMmeH
obE9QkjW7Ontml2jvdzzYnrSy1bQ/2d0FtHJe7LIwH7ZmbCyFwQdlKZEJOWxuc5+Mv4RgPgL9jKV
di0KVYQyUiuwek4j4pCGaIVENdPE9NkymK8xA3ZMtCwH/X1JZPgHoG7wRT50SMxq76t0ZBeWruF1
ZKC9KwUuDLmoXxba7G/JorQppSrgTiodckXrsDR3bzWMRwC8nRvhDshZpJI9WSXTHPd9oVSnpCsP
FPh5O1tXDDso1RCW6a/H6uqVpGCuNb0AMtp3fLoBKv35OYkTWMew1+I/6OkZxxyHo00l8jF4MdX5
Ydz+TmN4R9kLjU5AfLVKv3wMQJVlp72iAB21xgoo58QadcEyowBaGhstU/tTtIy8cQ00MuUEiRuq
yUhbAWYpVJG9QxThuO5lpPtQWbe/u3qVrLC4bmwOz3MdYhW23zrKz0BOQNg/wtfaoN1IFMYs+Eou
04aLhIuPdjLLzvMKEAoA7Vxsu/gUu2oDEgXPgMtoR9PMir556T7eFkBmCm4VbycIAqUqvraOkGAw
H4NFtctDGyhnFwdw0gh/YbUU/o7Ilove5YusX3Xocbto+6gCu98103Q8loXLawiArmGrhbuTt04t
tQbtpPxQ3YdNjUgaOvS/91l7moqsL8o1hx5Nf2Lr/WzFXY8sgHEJTIm2RikDyWL+fG5I+PzRJQFC
0mlVyUtw2/Dfd2sGeewkGtZuNEAZsIlzK4ZTqkdsgQdpv0vZHhSP80H+teFvzSKo1JflE4yfVyBc
naMJ7HMBn5WQm/rGEvO7nh+2AUMhLcX75RskzXKIpB6SeGsX0Tt4MUST76/ruak9fkB9aLSYQ+Ex
TlFB6ny2ZTE+BuBKpAndxDXIUYmUtzo/lid3VilXPtcaePUfnfhkFwrrgq4undpSvR0M4pzKuLXL
BTRAhNSW/64qbtm0sJPAJARByhKvnJJFHakQbe7T5w0yx1ouqCYqLXJLNlzYctGVSYCIB/N14/wW
ENrHL9OrX9LEF1ZhWLnw9zq1Bxl/QYQcdcRHzmoWadrq+mWtLM/kFwsJdsAZdBit+Gs8+dVC+/ia
6j9QyRaU/6r8JohEtcTZcfwYpYucbDInI5v3sbQSpNpVJCwuj+u5mFrFdYgNFHHMlsN4zMtSVpry
tnnPUAA7qstjvtrnUyxs97AAZiV7mgZUoWH/IDG6MZEMa5tuFolKm9LhAiXL3JZh4Ia6kr1X4ubI
g8H0Qu24PNrUlmGvVq37jQHteU+08iBZRvgzBMOgtVlPpI07LwkLBXmwAWu2C6iAedeJqRoS9Dri
avALlybgDEvEjNx9kCfgHF2Iap5/EMOTD8Zz4Tx7qcXEmlgh/UkpqVSKgcSb45Q5QKv6UxHHDR45
7VY1/upQsym2rcmqLY1zAqZ0fKZw8TD1vN5Tp5Up4LUaPpwy92tYjk7VdUr74hS5W3nq+oaAS2Bq
CpMYMELILw0a9El4b4VtwJPmx4csStBbHkoWtOH656RWcCuqxw+EAzIxvgZACAR3vCFA2UVUR10T
gbIo0XU3HQhmvo3pTg80Xz/WPHQyK2SSG1sASAknRS/oY3tYc/oVuUNkkuQBcbGhTKYrzHLtXTAN
rncqtSTDjWg/MRHUm1kMkGRSm/sT6olRU5YWQB4O//K8MNa35Tl+q45Ed2LFb3pk/waWon3mk5dI
wI4T+oelIqY8sB6F+AObvCvCXBDVVLnqDjWTi/LuN7TJGeQ3DJ1ids441pKuPYzjnjtanvGWaJYH
ROKm15XDkUf000KvkWxbUMe+lSmrwP+hlJpYAqmjplNn7oNRLYNK9+zIYiJZayVnLFlEjLbYjXRV
QTMdi9RCuGoWaLmQhWf6qBqFTN2xd8p5Lz4+LJdOkUv7aE5B0bKdzn/hNThaki1gwhHC4p6XM7eh
3VVOkvd63wp2lJUbhs7MP+FBUjTk5aKYcOK70BXz4HzMXJiqEJtK/wW5Goc8BsM260sYClIgrfu0
VRN7J5yrg2VkB9Jf4Hi4cM+9wJjKwsaF3icqM/TH5V3gOukucFVT2XUTlKXRzIohS1GbJc1EE4Vm
qwvcfW5So3J0LH4gaPPsURnUmZwOnhvSQ8IzBnXWZWgzj5cQLOe1TnhTeJ3cS1C60dBjCuW+dZgi
qQAFRUUYCY81Ri/PvEYDAXEI5thbTwgHzdKK5kK1dRbk1Il/AZJEhk5X+u0LhZ3BdD4yUt29CT/7
eNjRh7ooi4xP1h1Rye2Aj79iyaBw5tIXdJ6zA5+OktD37SgPVia55vBLai8Q5PJj7Jmh8s1e3WQA
OzKE+ZqSwPLraAx/Ah+v+Hd4p+9pB6SENMDaOzIZrICk4cPTNcTAlGZLdFalWF1BwAUX/qxzX8La
4/G2Vs2S/7znPldoipwkGWf24uG8IZiKPeHz64xTf046MqByV9NwYJ6Vi2+/yRjL+iKBk31rbrdx
+mwFgev7Ml+6Qduu7KWwCwpa80PNq9KO1oglsjDMHnUDhZFqML4ozOAub/ta2Q8B6lnC7zax/snV
gOGSt/CEpQ5pvsy7znmjoN2sdZxC02t9/NU3IondpquM00vFZea22Eg/5HbsNW4k4jWcxBZW26Uv
Y1fT+yS2uQUuT83iqR7EJ0RRQTv46PlCFqoRaNtjPj0HNWeRAaFS8Fr3TAOdTHkehnH3QMABO+Ry
FTfQErFzuy4AVabI4kVx1zQwx5IckfW63glz8Zvwm8b6+gi87n/0A5IJRhNFZG+pPhaA8CZIbH4j
DYwD4fodDe5CmQraX7QutCXTwAPErVz14exkENSPDKnX2gGU8X/MgRHU3DomxxK4hJfGXA89Fw5+
PPqaOMQxOL1gCcu4UTTaksMrqsT2WRig88O9IC2OaS+9q18PvbrsW9P/WB+kiXeyR+Mnf4nJ3rv7
L7k7hxivjl0+C3e8YIfjGbBONQ6rYhJu7ZMKmt2thbixJpV74CkjSqqT1+pLyR1eght0n3BmHH3d
RbIwJry1Js6WF4Ug09EmvaKkFzpXtuThghpGqzEvircqYEDLGHvs26kEmKPkHAIDW4402bSiLn4r
+uMm5kRhhTA4RYwZvGd95JZ0pWdSOpgQulxz3STAA+b4RmJu/PCzMq7lZKKdf+TLTS3i0Af64HH9
5P940GObQPDhf8rmPLsYkKh8Cd6PjY1MXl100VuOuUScI8hVNlGmBrnTC6I1Id7GbR7p+w6H0+aS
lbHhyp2FPklXRp5vgB6uP8vJpuszJsDbE7Au6upXH8Ogw0S9OcSktJcm+V76v+pQdAo3dzcj+2gL
Fde4AlLh1aUAiub/BfheH5UAIr6Dz4hXLbHCOLaCFYSD76ImXzhqNjWaPeeyV+doS4Q6fy9UW73p
1sEJKb+HFbdgwYFY3Jysm/pBpGQuEtHvh/qJ4Cdef6EVA9nfptselexNAIQUpgD0yKZqHZFedVky
8hljHxeR/OKGuGvW/qwtCkX45TT0YaLtdEbxrLkYbGo2lEiE3jEbpNyvCZPH8Yk3w9kYQOpcQfRp
7ox/G1YpdOzJHGxO9R3ilzQ5Y2aTX7oksv7esDE335qbsO+PJRe0ZM/dCsD+UN7d3ua0/Hvv4enu
nDOVPuYBHHTB21zza1HiTB4KxAZGSvgc6kRiAnOziR93cItm5mIqvWYy8Ar6FrycUMeH5KhSnvHW
kAuOJ7POfpviwEWz5Gn7ErlwLab7fXS7/9WucbCULIFolJEraHQe+Zb3qp9jvSRu+cLIVntGWLvR
V6Q89UPjokr8PwJ6igtDg6egH0Dgctj+Ehw7S1bbj1cCtRvF6iXE6BnhxCfqVmJams85lam+FR2V
w4W6A9/fpVLVxqbUoeP3goXu/bqj/NXbao9QcApUc5Mvz/tHVr3K7umvDGI0u5bR8TQIM3HRIIQz
CO2JMyDawF18aoJAiUrFLUdz8nxV1sDG3muajXGevHnnpTK9f23bDDI+59XGj2Bhx3sk60YR5ABO
YaX3tovoMTNufS8iVXS5lZ0Efpymg5MAak4iou/WDf/jLKgfCEmA1skiQbtP1Mw2eLTr680ot361
5k28gEcm/2MFYnAa0XJyN6ZjFulKmTJ0ZaRE2k+lB5/M9IKOASvKDDaIpJli36nIInwQjvSJ6G0/
bJ7+jqab4u1NZSD0Jx7uHwSQZ0ESFQ9l+9d8WvHZ/Zj5keYFon/rH4tA0iCWyIgc/tyUWCFSb4xu
gPGQfHepoy/wqFUe4KIEox5KWpLV94HtHa0mtk7x+EA1MBPpm4MS3sz/94prgdzopYS3Sa7JkRQ0
vAQOhAlJJdrBNjw5+9pT/2Bqe9NjTZVtEpacGhvFlYAMN7kL5bUv3CpfmcvbvWE1FxvxTOMMSArT
SjYqWkb1oO0Y0v6g2jsK8M/EE3/d1ZRbuHZ3w3OC0/mnie/MTZc8MKiyhfOJZhe/CFM+MYsq7mDY
a6l6+LIInKNpk+vd6i3N/nP2Upms+d5Pas7b9Y6foV0hsS7YatG/o1JRqabcD6oxW5O9/HF/6jJG
2POxD3CLt+8QIc/KSMMnW+HoKnbbdzz/oBaoQF7GhjjCzvBlNkk9WyMiqtQDILJBOmlUp0dPVCQp
1pDaV/S6LGqB4xl/CFd1/GfNDBcfAuHFCye1TyY+0E+fcc5kBUZhhjq1Z+/bJhGhobDqIWJzrEs4
1/cWY8QIjABLVNfXXvrf6qUUIulodSuVdGLstn4VuooA2mCavk1gfwhYLnR4fq422FSy2zAfqjLQ
gjQKm2cTGQv8yCO3FAsQ62ny2/RxFab9U0isR0P5VEMKt6lTu3pF0vLzZFxoDMH6z3nwhjL27nYq
KVPWdDX9qBTIx8niv8bLvE+pas01zl/Qv9YlYl9UcH9aMpWZ5FJns3b/Y+wI/uKtQ3dj8xivbfOZ
pJGgQznH0yjdeFmsj84L4Nfn/MlCc5HP9ErVRsBRyLyVlli+PgXBg183QKxUoC8rwmy5dtg0I4i9
1KK/wB/HOmpUP7Z9DXtTZ2OUw8EZERBImqZ0Vr6Ao/dMHNY2+pphmV2fcifySG4BQfbWXJadqUkU
BmXpqhcVm8xYNScAUgqBaYQ4iT/z40lMgF29OrPdwV/QRFxLjfrpXc/vDRi/HrbOzvhmzWz3qRRe
X/qmjO0l+XUJPt7QZYoCV2rUm7YnyRaC0tRuLiB2F/tZrUQF2ywRNODCdhZlGMquPSI49qsbdGds
D61J5Hhsas0K6sdIHZHeN1oJwWiBJiGm19nvXq4ibHAiTqpZF/wc8tc2yk2H9wK16sav29jtHUbT
ImnW4PKCoWKls77Lsx3Wsejqh71qpXqiPu+oShyA7xr6dGeQptNvT+orZHAIp8mqlpPzmI5hxl2c
aWFOpKXXMU5XqzXgtHqRRISWyRpDldY+B8IZ7BiJPf13g8vAKjRt8RisGIm3kGvT9ctMZ6ghEAnY
O9prfeUExqWCYqU7ixbpPEIxZ3RU+mfd6tt2RRlE0swSVVMhRF4rwEcnoYskhopQXLoNE7w+3pNw
AAFnLi19tl6MV0IEjIf8Y+ErUODL3WsnPAf7BIkQTAmvOHxEJGjO1MwIRr6ORJvCypB1vW4yG1A8
t8k5kmg/MyXQ94wv1hnITmeR+jWVi2Rl7xS2BFaRUIdHcIFz7fa+OjE6Izi0lcxsTgjA4vGKpcbX
ZrMJTyuiHcu86+1vtSPpDTJ4c9GQUKaLWoPUOlzPIwqNUb3feyzoNd0yhRaSlw8LQF0HlRbnv72E
d55+QXTv44tCuDV8iU9IIL5o/6ix9XNsxDWvO9GI3Vg1hOvhVcWw8jw6fnxBsAA0T/suKhF7gS12
BdRS+qpU7DfAjaeAaKHJB4s+nyNgo77rh07M/s0pYVoBKaJXPF1tcK8KQzXRUc5G5DXL09HWH/tv
jQhGPRM7n50HCi3brEGCXACXANmfFm94J/NheyZMJqH7IRVbn8bqtt+KpcsVtSwNN0ixWP8NAYqj
rBWL6T7ASk4IojhKzqF1WBVr0RjQDqgv0duf0SWenehKCiT9Xi8NjH4NvTik0wiaqMg/3JcNukRF
5N586zFJkWhQGME7sry1vF8IKVCTLdB9k7gTwLu+t9ZA8kxC6RrI6SagQjpHPkcmiEmP0OL/3aog
yj8sJ5tnQqhEG93mOz/bGCSmd00HqO692Sp0ZulTFuFBvsK0vg/f9Kx8rf9GJ4YkcaAI0XwCb8+C
vKJwsEyxV3qn9T/0S2f4lv3mzJi8HcQXvXaFWIgZEcLUQ2j3YJuTdAZMC2kMxp/74xZzOaVc1UUQ
R2J/iDw8R646LE8ZdlgByVG+/VB9ne2+V8eIs4jDl7nTDEhoHDy9ZXBGqmhOzYcMDdSmZ12VKhKS
2IJyQqk+BPOtq1hkeYYFB8xTlmR0JnpXWZy70TjAsFvy96YwiJSzG0CXbnAJ4EPD9kxY9vI/5oO+
bx19Jei63/hMLwuN7nmGnBvpRmEdK5/5eF1yAD0Ekg9xjsSND9nCX3SN3LSMDRlAZN4+dUnnokQy
rZeTnfLzmtZNyhbN6hFD7/nujqhM16m4ih2yjiXAw7AkgVFvntSSZtGQJRpQZ0/6cy8OAYa2JZAA
u0f/97tyCaoTsZyoQ8He9NjPXFU5QyObVWO7MDrbpa+dXQubIZ3pB/FX6rtnla5+xPUNnaaNGG9A
+LtszA49BfJxMfnGLARE88xS8SiT/qdec7A3ux1mu4vD08cfu/WZqm6HiAt3Sg5g+1OOQbe8bSkk
AmJt7HGQCeoESDDP+Pswsg0Q1gxaxc+OAIU+irO1SZopR/aJ7+31Xvj63X3Wyx4uTOOje5NrW0lB
+4XlyU3WjShVlGgSd9lQOBvCsE5MH5tQCmF6bDPrH97B99CkNEGIY/KHupV0SpVCxhif1x2lfToH
8IpwoH1tVwZTYxZLQ3t3Fpc4ysQXmhZOetjNG4ZTB/QXPad/S67con3xQVr8Imk/aXLEUdiKUjUJ
a2GduJLLP67K0CpDvibzhqORLAJZFK1JqX1178wptC1ZDNPO7en6uDBh7mOF5g0K4h120VjaxVkO
RLBmbniHcNw6ePJFNRTv+h0d0tBDYM3fzytug9be3rLaPODqcLHlPcasfiXR/cmp5sx/ho5xsCmg
66tVeMcrpQxtKupBgGk5vxyq4SVgnF/AxkJAjdVcG5mibnj6on3d5WjRtNmBdj9SwOagZ8G4Qd1u
zBOooIZ+SBMrlyfMc88KKBaqkiiU1qqtxJwbmxNuR/GqR/6pKVRmvMppPnRqDW7wzzn5r0lXxIoN
rrIs2NROLJMIR5hlWTshWYeYe28zAfABm1ZaW/Pg7BgxuMPZnmRYsM5dqOXh5Ue1yqrhtuBVqPc6
BNgKX0w66/pgQjYaqtWMZR58MK3J4xyBaKvj1AU8DRQvmjpaERPQn9e+gsjRTxQEEdkl6+5Hyei5
Z+dxQbhjECa7uwJKA8lu99wU+vbeLOezocSsxj57J03miWCUOpv7GolfkoBb8i7t4uYbIOdp7yE1
QPxcA4FbPmtrsnUgFvo/seBQGzLqJwKmhOlIPu3HFnFK93FQVmtjoLdcECCoBFTAQuH9l/yXKvXy
lYH7kA/uBPibaD1csNlDU4Cl7vR4+NvCivdxLf2tA25PDO915xTgX2Y1X6lKwVhma8lXzmo9WAU3
kb7cdNh7priLkzA4frtgwIKCHJtl0aWjS+g1hYLJqOe4jNvg45rRPlOF4QorijpS7pSWfGXxGxQd
J33vbvAGarFof7gadAhuxmoF6kLpB84LKWtcpyWif75Bu2GFqXJcrAuw1tDvFexto/N1yALt8jHh
YW5mbguBJHL7a4tSKI386xhSfgHxATZ/8yvNWsj4hDcDbgoIDp768TR3fH0ot0FVfbGLtSWsvxbE
jauq4Pl9p0JN2AxcnrcjRvDWE7aaGuwBGaABFNQco1Y702i2uaNotuuJkWI8IvH39U/cBxU3GzGj
A+KDHWCcE6N37pNr1VbF86XZdP7GLdfMo9hlWdAWY5L+lDLIDBddmsXXJ1fwlD3DWfkIOHnExk3m
O+9rsrWyvwCX/A7sgPIBZmdRhNvUxE07kRHhEfrEMg8QmWoUveGYSN/x1X8+Px1LRpyU/MLomtw8
vB24JiNYPl2Oiuw5ZkVYD1U5BHqYpcBkzPKGxm9yPS+xxi95OFVymRwOl1m6tvEwwLDeqCT3Wdyj
h+roJ4NIVIaIB2/2IFs+L4OOiBaTKwwDv/LzWS+4/rQQCcMx4DDyZNju0V1Rb6RD2iMfO6fixmu7
71bWVBLf6O2GAhOYCqxeysFCr2Plje7fQSzEkpPp9gB2ZUmaalfk2qAUZ7Mumx14nNWWKhm9tHwi
8LVHXk/dJEQoGCLwfJhYYBJ01C6vN1jarxDDhEJ2AjNvbOp/dgMfuTsp5iThr+cZ0aVAhVbVhFmm
ndxbkfiLDUvU1K3F71olDZsnNXTgZou9d1xPWL1oJRenA83QNSg4Zyo22F1afb0ldF2xRs6noBLU
x7f/SDoAYSQDPJ5y3Upo3V9ODGEuT2Q4X47XHSvPpXuiKGOQ7Db41XAeRSalaAvC+KzV7aw3Etdf
/tUh+btUMZw2eYqQNoG7euvPVtqyI6+jXf89zm/bYhvGh4kjePC6cuBV2EU+HuWUWAeVNmeju2gE
9xFUY9KyXw6aBjIF3sCIy/8ZF6CeZokzg5cW9NZoCVisAqDxgtMMuF61wLe5xFeXU9KwrsZUD0T0
vomqqn/XeJXVbTPS0Hrb/LofXDGs4ebPN9j3OteSZpXQd9w86KufnjeBcLGjMKnibtyYjG5t1U0X
qgyonqJRZlbo5ZMxHpwy3IxIWTJkNMaKa1yvUb/pEWS2yRQ5fiKbeoBQ8M0gBGfIc9+OxQR6V/Da
0LPRT7sb4sV/4/cjenMXeBqHEc2uWUoedzgqWgSnQl4ky0oSXah0faJpJXaoto84p6nuAxtM/egS
p+XhqPCDGZQ5gyTVqhB8DOfc0I5swR6j+pdWB/+fcKPR63tTo48nSsfDsI18ezzGedE4MAdNrZKF
wAQ7HDMmw98hwyTWG2EiTIHlSN0Fm9RokL7m0AM1OlmSyuMWf8lxCYpWZntn9Aj5ODm42Hup33Kh
wuj2DtihBr3VccC8kfYl5NVR+z9dqLEK3ex2tVU5DVe7nJJxXvZjoKI91iLNofL7SNPrl897xTGC
sS2jTBQ+mLRKkVRfLWR4Gf2niL9WsCnNofw8tHlfLvzZnYSUjH/dI22Q2qKyLvkjAvA+Sj0tBON5
7sNyetW44B9it2SMD69LXkn+xb9H5jnB6mZyvko4/WeY+2H9dKG/1rACuVFkOl4L0lPFJ89N/MBs
ySGCL6xwLW9N8De4A6KHuvqWoYWUo6+W05cmlNDuq57FUv+6ymMXW8fjAB5dQ/e5TqX7cpOOxwxv
BRdGVVniK/0WlhqN2CDiuL3x2LKOlhalEoCzytgSm6n+9CS33WL6SufiS4/5RwDSObVJXwfqYugW
vATlYADGaReQwJytbxQppF7uIs+JmCJJqL/a53SsFojdHDy1+axvQ+wHK5CqRfOr+6zg29Mtl0//
8t7hiBjs+/ZQQjuPlq1uLbjjE0xTSCryTwGRACmtZ08F3GHwJAdCp6VkMSOwz5jA3uPSkcfdO3kT
JC9+JPdfy2DVvAbAuIK3NFbASavoEYvp8gU6YddfIJ20y4Vy0DloXygO6tT4wZFw8VH0Z/iuxQSE
/GQtN3DGTqP2ApVObCjj/4l3VVeF2P8hCy7ZDMosrV5U1/uGCJrYrUXnCUsyLJLtr4Ga399AGiX7
+t/OfKn7Drv6QvPtbhkZDEyHolF0oQNUgv4Vnn30jXrnd0nZxRYGvWISpu+8U4uCmcZXRwdsu2Bl
I7z3yYWSNGXoybzWp4PaGYWoTfjWNzJ7xFOF9rx1jAWamddVOKAsFcgppJBwEz7DAi6Sqbymg7YC
dfs5TjcV/FECqK7b8ZVEdDRErN7afLMXFDyMAGOSG3tpoDgpGVrQph7d9Sb7Cvwm92aUZA3xf4/+
8zySJb5+Hpc3k7xj0jDoFPK08V+xjPytuVlUtQBWHReUBF6FVH1NBnDb7wpqb1z/uqJ0VWTpit9Y
nX6QfzgbcECDka0hI19YjZrt9n6XyiWPotpw3AcfKcGxftGbnICMtIwz1SVj+AI9B46aSUfcR7DQ
hgSkT4RWVENoy9+y4FKcxf9xwUP+Uns3lvVbXQ1j9B9M2i37LR0Ig+QGXAXmdwZ8CJdvwwnFb+4K
mc1PW3JlEiXp/ACa0MTjG4iYdqKiuAbOLk55/YtWDuaT3nABh/XSI7QiEmRFuQwDeN84QEwU3q6J
8TtboGTxw6DOWkWEhR50vDCI0Yt27stvH1eRBjEkIWlq8hN65oh7oYMrpXcxQ7zHtgzs6SZWZ4bB
yqyn0/fyd8KWIs1qbJPA07xoTbOQMTOoyzxwWivInTRm67X3NY456jGx3hddhZNejXJ5crBoYPrk
+00tnWZf4ab9YLCE2R4nU7MY6QFEcRdHMuZWpqWv+YKl1UM26ozK/XRUG048wBgIrYRj4dFXbceu
+vOz7FlCBj4oDr1GyaRHLy6rU7bs1LBO+gg5WPbTwRN7RcbjX6j+ITG/A886kp/rVjfs/2mlPmfh
4CCqw7K/e71+I8nAB760fuCvihZI54yNzGnADfSv/9LSpm4WcF0fDiqoarOZcoMBpkL7eerMFky+
+W1pNmSxpb6ybiRL2CQhCTbEShRpAvVR8wiTSn9aEmGShiVbMJVGj6Jzyxpmts8DPDfqHglu08O3
fQD02FF+Wk2OAM5sTnpabjPWnxYmnEyM5ruwYSU89nB1TG534Mrcb9wJ6bvrPcdx0zjDrAlZJ4Is
LRO7mXz0O1N/reMl6bNvO1UTmS5J8HIoHPduvENBo2CHqRtM2fj5Xv8jNEf3WzyTzU9ziYx5ycyn
8uXsnJcnqxY0ridI3UABS9u0JrYCPJxUGeCnYwWmLPva2wk4C00tAkoVZv0VFHpbwrQrh1aNlOvP
MWND3+3YFc3XJA9v9qMVkIbIZPDOWCYtxGRvoThg1hRcFw7cY0ftN5aqYU3Tn1xhvQtGlRkrbdAX
h5PK3kSqc7k8uMzPL+wdHZ2JuhOVfYyiTxaGtKFSaVbystA+U4DiuSESSfOJ51ixTbqNZukvNCAG
ya0lezMqwkr7Wa+/CDHqnL1uf3rNQM/reMVblzhLrGCOCq0bIuBsNdv420xqJdLmBBX8jZEFnCxh
d7XSKFlB0doB+XQMMDsIdZ7QuQYOeGkzDAX28Vp6/9N+Lzru/kDnCD4FDtB7Npan5j5kuM3RwfHr
FTKRgeOBvOG7RYdBvZosquZ4/0CMuZKFjLtALnbs1GsRY1Mi2Of9K5B6OpGzyhGZROp57hUtqlJL
4dqPXzFQtVgTEpkS8Lp1W6i12UMMUFgu0cShHjwFelmX7w4pUJoDj5nQACTPJRGaFkFZ2N+wAnJZ
LdYm8lbqD61gQ9umGsWlB8g7z0Hu271rYqfPbXA7riD9F1YVKL9CynEJuTcPePSQ6DVC4wTgic92
2omX/6XyGLOLk85vwugFDIX3oG4FWuYlbkc2GaO4Rjwx3J6Qbkm7fsC/zpiPfJ0G93yvj4fq0CHs
lOxmCTZ3aWtrM263C4YDOWJgVyeJS957FPB/2D2Fd20/YwYh3Av+v5LczmL0PbcdU3dVB6JSzvDW
jWV+xVRF0cXYpRySWW/ksZS487FW52uTx4P2twst5xFCkcezBtXBMdzzew3Sx7NIUeroAX276x6L
OogE9cCrPAUfhXexqG7nil4/p40UFXxPe9/liX27fyyl+USLG3pS1orX816Oc+ZRQ/OfswScZ5EE
S9auX22qEPByZzqbVZMWabkHf33OvhabNv/IbZSg17BTABezsiub9297/ljSLem/xWkz0PiZ0hh9
yQogOt2sPQyD36nbAKM3XlEcf+iI5UD9/yVVbIVYKsWN8yl/PGEwnf7jMbG5XAvg+PW1TqJisAmr
8w9NpNDisCajf8XE0TEZnvI44nuQdQTpPFGgE4re033lds2Mf/dyetgPAkknip5shbjozMIc8DYb
5OKc8IDJPNy4T1jmlZao+QJ/6ou4qXcJfAC4b3+DpZhQMsFZ7+HQ89sdCnnlsWzw+7+w9oSmCOHz
Cj5ivQbW7Zgtt0V8OARB4HuCMpatlrBc/op9b0GmB6po4GWzB5cAcQzdRVmOACv8fXqhDbL0tnwe
CsVWE9b00vskT455VRkE6doPfAD+k+sYAc+hKvh087EhTXeYaFh+om1/r788BZUN0ePY1l2wx97R
l6eeyK0lRAaaM9A9f3yDGDZsszI99eXkEYc96jDMvIi6Q/XjywWievWF2mlRT5FFmvos0bGNlOhm
YsFnRAfuuoM4BA7v0SvoJt9fuV/LuKXVULEk56W61PewXrKJ9fRjXgOyI0AExNmWUEA36RnnIDSq
IsdXjUUabQBGGAU2FdzVdTSWkTKU4yBIeHwp42Mt1IQgpJTiO+wWsTNq9m0ffJRGfiITfb23ecZB
K3u/imi0xUp6Z0WvO6xWZQTxY5r6+zMTjDEW/dQuP2xGkVJLx9InOu7Gq+WyPbDweKaVDg2E8gGg
mVkEaeY8wHxIFTzzfARhagr4/hEELhuz+ZajGbAkm1e6WMBrsPFK77l064c6TmwNqaIg/yhsbv22
IGSNdKd60YJjyb3OmF/j+7RKpdMfVZJupSZTGqwQIz5U4xd8NfTPiUdI6zF0bIA6KbmuRp52T5uT
LEgF9Gcwt62nKsrG1d3pykVxIcrOFdebM3dXzNXbRf+pODFI0Sq5kiYUFXeW+5J2EAk7u0/RD2nh
1yBri3lL6b9L3mnboPz1Jx+1LzBZ7WVlq0Rd/Ee+YmDxAy3+qR6l2n14rlBVM1+wmj/IiYJOsspu
V9bhzBYWKvS2wyw8oysVw84PfbJkKX9tOA4r86oJkN47y6uV6FJN0R2UIaCR0zZr4EzkLwkr56sR
g62Gve1u9yoIB7oPmPuiZdHqRVJJu2fe1HJfXzImfROuTNiudRYbW1xo4PfeYkQ4rsNE7/McE0HS
y8Tj/LzlitnG7WXpIqxNAgY8uu8C29GCWFMuTT13QbhUcCHD+1vAezUNaCkUKL5JslDq8Mx4foLs
UWJbE5KHBYk0sOy+6ULHZ7S13ykAc7VElYg9Bml4e/GVMlxYEXbyX11qeUIljzFNMP/JzHYdiMmi
WbB9te5+V8lLR90h38OPCuK+7F1a3SfqiDIcpI/SLj4DndDJKNOMCw8rWQ/7eAhLNVOhtNlkEDu5
amtKOO8s5LJapjKH5Qme0pXMCoTdwxt+Iao1vIxXUI7n5zGi0xv8aSZZUh5Rho9Zb5eRB598lteW
q/ufdzO6sSze0vh1u+dLuXR7Pt9f1BDk9K3UwYcH4ynoyV+D+gPZOaOKZNjinEG/8aKStVSaHzE9
tXuv1NBbAYYPxZZSxZVsVEMi2XNU09b6ZSfRosPfoQreC4rShAGAgxkb20Gs2mrDigSSu6gRF1fn
AYMcGgbAYvnwhFLa1ZsJWcd+RAwjaWZMqC+eZLpMRPWyXagm/T79rKdG9+CN/9GnITgVlWLyJqsZ
hNuBO+O4MsqzBSTjs1uzPdPdkKC0mU+swt6xAvbcV8XQwuCsK9H1plyyVeZq00dMm4ZLyuw5J/ks
fD5VTpBtJdhdj0m3uE+0GYCRuEAgdU+X+YLJLPoUuc7ie6trAuhLUkMn7zUtgsYEPh3ejgfv+K1R
tkHJAAQlXAgI2HKfOKQ1SyfoQtRPD3HEFzZrxMKv2Ereuiy+xE+YbAXztXqncL4rUQDNnAtuaKjY
qlHSXTVT9fEL4cpVlMyFqlOQIc2NfL1J6ikyD7dOF5ltDjsRNQwumc82V4Y5M4KlIK+yW2wfaivF
6ylKgKPwpZh8Uhkl6SVN8FIq8Kukz8jgHrc5avsF8Tr4lnzayOt5HMmCkc0JbGS1o+oChvlZZwpC
p29QhsIsSNgFHmgf1aqotFHYpzT8uz4eEkldW/tT2XRKg7EGP+hTYuBVRKL5uSzjSaovqeb6sH17
0x+jcDXydW49JEK3FG+UoFQT6BZ2kBr/PqQtOBnzB/1dTHH9y0t9/C8pRoZN7c07kxSD6LUWNPP1
2l5J95yeaM3g1eGzRyDitmNa43B8g2r3aDWFCoxN//NTV5scOMbx6A4afUdGx0sSBSK9a8OhAlb6
9TQpZYs3K9drG8ag/G/ziF6DNgvfhrZsqSn2AUul+93X7meqSMfKbxW5hksG4uanyu+6abQc1ffq
pAc2NjPU0rfsMojVSbYbc0lBwlMpXb84xKtxSZeawZPUu+lxkS0V8EtKoRPQri8o8PwoJxxuuKEC
3jxDkh9tUaLDcUuFQbCZ3OVh9h5YKSrfOohx2r7YWKJzx7O5t0iJ3Yg6RlEPxWVqpD3DA0NQmAOk
Arj7nSLzEX0lt1u0WqblfofXBGarO+BxdLR6x1C+c0uLrD8CC+IG9zf+dU2tEAvzY0ILcT1CdJFq
FT13N9Zg+jQaTeXIhzLsO16blSsQYgm6GelSC3epDW5a/AmeAl5CTfvUWrdOVNbpa4A2hNI7mUgN
fBy74pzfk5ddKCa11gKIJUqERavOvW2FFkUQvY1WtRypeHi5qEkf6C5K6s9SkX0wwMKPgVyjTfYe
mhMNDTYPY8ZFyPcCF/2/SmYEl5tn7h45nR6p6ktUqGapKPGuz8L5eZAxIcXy7v+kQ3s45tpUTA0y
igg7mZMl8FnvGguGegYG72fgiSqvp2RvWePKCeTlbqi2ucTTmwv+svblPYULFKxggWM66QOLtgvi
Tn9m1SHolvrhA9U0Lq7ywnl1BnqQ4yFvKEniirFLkFEYraC8bVxojpXo9Go1pEeHa41GL8f2ieM7
YL0gxcCiBcz0qScbccnzc3tKtsStO2VNzLVjOS+cmGmJ83KjFCzT3w1s07WcDuUiGKxN7SBcS4a3
HO2hBv5h6y6vr9kFnJKgI50qLNoZXAyGCf4ALy9x0sLfl6MwG+1v17kexkMIy3xnaX3xAgRfIbW0
gVE5JQAfqZIelO7eirqaqS2sMTXife7XXY4VZJ09y1iJXEY1HHZFybKKq7LOTQiBIoshecNN+ZcO
TmUz3d3V0W1W5POrvmvQ4UOS1hrj0HzwE0q/Z1jlOtOmYF0XGF7kVvp5Fbb4SSFFwCJUDRtAgY3F
sMS7vEwUKafEsl8p17L+dP+iKIXDiEUQF+QIICuLcmAFvLJvOKuoqTQAu7NvTEwGoVvKXXx45s8F
oE2q9ly78H/Q0fZV19hF4LEI4rJSz1/Pnb9OQ+nrfC9CYZstyygUR2RagJX9insREyPHin5davPK
75Fp6+qflKqMj4+izvNavRg0K1ghVWY5e12O3DxnhcDrqDyndyPKKa4RrRzJpI3Cm3OujAEkg2B2
LjNazXn64YUTk0TMZ8ZNEG/K4VQGZLXTKgYcAx38JGGOZPpdgng6NAj530J7F7EPkS2MwBZRS6la
atFH6boDvYFM1IHK/BTP8a0tLhpSoUe99XWB4EiPcxCX9LIUNAAX503q5MpY301tBMaiqLIo4Um6
kZlGz61r1nbZ/re4lYfveZbWvlBLej9LFc3Qjr1sNi1bdLVvv2pY/SSrPEQCPHZhaJY32vKGikF0
ou07o6vXK4JZKig/XjIwC67vFylH86UGGo/oruwnmdDlVErmga8PFdyMovi1AjHL8+6F2jvr7CaU
9IAS8k4J26ua6yw4TO0Y/XdCAWLNLKnDEU9HIp8IJ8FeKKqavpYkAqbm2tNFCn8ecfPTMk9ixloJ
sAvxCd94BQHy/+umgV691oIFIKssnF774irTUvgRP+hPoTyJBFhd97QqjXlNSVqBMqCYkiOH8/c/
6HaJsSAoxSw1TkPtj4u+AbMuWN422PTPV2J5eXPlnlz3UzuPfzXkAk0TRSdHE7ubnyA0p2zsknrs
UGGIfOUBg6tWSMZ3BTJPqcvde+GQuZsBUJxI4aKm/xC0xl5Th8+8CasONYCC7UvNLtuITrCanTPb
vZrFHClbVmIT88FWQeK+eww/+fAheIBx74APLnitJslNhnvsQ9zzZ7VhpkFL5P2SfJ8dYHtJCUQk
Jh/dkBXiE/SpkkzVOIIqzKb8/NkeXL63GTPydiZIxLgnKYseIaDvdrgFDPxv9ACHIH0j5DTvXi4K
QwKJeZgMJDtYgyAHd3iMc50RE2Dvkl9MggmIF/zyKWrb/WQdpDmUnJcbq1tQ1pkqwrwt8UxUaBuQ
G0BwpYWdLtjWNOFFcd3XgjAICRInK7ocn6y1AYiOsAeHyRvnImijBEebG4HRjsw2WT2Pku3ujPeY
1vUs095XXTrSvJ7QarL/UMmgDmixzXzqSjDI637Ca5n2k6WrjKddce89MABtqkZ4gBy6f3s6fI/a
iRxAFu5ZR0SJLXCp2rSFkmOMYXmEwhaYLGEA2qipdM1bMpFvSRiJ6RSafrMc39cL7YR4DUHqykwR
87aOxiaiQAaywawOiAtFgcPRm9U7MVjRSdBP0YxBlf0+3P0Hgw6UtL0oNE9knVuaYsFU3W4d8Rgk
64LHyDNMZ75lT/e8uZAV4DL/OpV9Y8kK5ZCPYrKMhT68WqtV+ANTe8niyDu+/yRXFM6Vze8Bqo2s
pXSRmu5Nq5pFOnBeI/lssAH+EKDc3FT9iiEPSU5uYgtWgGdZPksRjYBOYOXncpbEmnqSqSYgX6oT
ouSp6EAAjapR/pt67ObcbyNoIXrI8XLrWTLDz9xAbKuFEdfVw4pF1pIYNmxbkIR86uUEqslt/MMb
KcVGfTZxKeNb5Puzox7lUixpqUAdAnv2+J22lQbditqaVqdaCwa7ulEz+6CBGWqqWqSPPrinDDpN
grRcaNKJ2UtxOrvuiIQgaCJ3neJtA2Wn4lHpB+SpOqAAtDdtFuFTfcTG5XQoFKH9Am4QqptKOOoL
vToTtaA1IhRxqMwTNqisJCdsC7QC03DfEuFch8g+LbSrN3UYEdAcjBrKciE/ztviGBzo5KRa+zqR
9Kwq67ISpzneAprxkL7P35U1QHSPBFDk7/KVnVOezE68OapIBWKKfqccpv8WSBgVXW6+QYl+70ca
IPjdibl4+6LNic/JmykCN/fpy4AMToCQ9PkL0WzbkhT2QjEE52K4te3d8nEZLMPVd5y6Z5Zh91e6
Rn3rudmS7rL44V+8NDtcwBAlWyNT1EPpDcJDj8z53DQa1c5w6JUYQUISKj/34ypX6LjfYbOw4P6i
g4vj3LZUwKgQwgPuQY+Z2g141INGqCxApqduL1aq9m2Zwnd2MEmkPtk3yPcEJib9oS1WQln6/7kl
rONl+gix7LLP8rgbui+va/OxFWDRZgxt9tqRS5sLXf0jEdBvDziDYLqTdxioK0Vnm1T7ub80EXr8
Kc3W31BGawthdFhti7SLC+vt1E5EBUH5+SqLH5LJTRCG4DCAWRocq0kSlmQ0fZ6+k+KYqOBUWrq6
nEFNLh7GUocuGMkWuVHN4p7uMk+NBEbxfsdf7TSjv8w7hCMJbDCrPlNpSKRtBQ5LzusDmWj/xgmS
2d8W1l/C6AdmV2HTefpwSNQiWLn//I4NxXhvPR/w5pa1L6AJK/FLYOZc8Gf5a42+EWx5gR5/yPAO
PuI7LUsuBBDwwZ6qQGKWy9y8PBmfaG1WCQZQWOJXzs2Z7R7DXUHOtv0QHybyN3O2iICc7tq7GbNp
P9SmIS5TR8su8VU+MDYTpLowC+7vzPcr3ztq/LoGc3tmblCxAcbUiSewWdiAQO+u7L+A6P7bNUbF
2/6SU5EhzPZHQlUS8vocUY7KN6NBCPQbQ4gIfl1E35xydociH42F0jJotJWP4282KF/htIiSyyYs
NxDFnGjrPenDRwNLHdYFJKPorSjWQN/dOtmUc4eMUkN6VV3wd7k6LQleXk2xu3QrTA3k2Uzxdb8O
F3YAgk2d67W4MjjVGLhIa/T95dUVDVWCvFrgHvqa1/YLFFgozITzs5OtT8P59/Dwl+r+XcPh6xN0
RTjkUIbZhXkEhb2uoHC/7sHkBBufErm/vJ4yX/IPlzey39Osmf1SXzzBm3jlFRiT0hmDTU9Vv5sg
MbUYpEPv/eIX8KcFZPtlN0g+4hzk9MMsu0+K8wOsTkS1vosGvzYLKzFDhPHxOj4BWxuWvLjUcKLp
4zj9lFzjF1emTe6M6Dcb6cBn8qzqnkaJIeuUL+n6xYNI/Pb42sndUVFNDBCbhaZ/boPfwGvon5WS
szOdjmaa77XZUIp9fY1jQD1L3/8UvutMaVRLr70uL5WM6haiLefdYdVjkK79xaSYW4J2G+aMdP3V
7yVh/bZZOmWWx93lwrC2qLGJXy6lvWm4mKBM0rHaC1QUKGPaqEavqgStGMaBoKrwjKynmh2QGmDM
7TUgYadxFpOJ/dSGpMTA+52lDXSinFFn0rXLWyqqu6vnRaoiugvZDSyV+uS01IJiyPV9Ytwy6EyC
uZtWP/O5OlruGtG7AGdLU4+Gfr81xPbrTeU6b4Dcw1BrRA6eDvUypupCCtUv8BfsvPu+CKVXaLR1
I/A6wH5sNKTf4S9hVuNRXAt3CfC7yz+2gOpSSn6yo9FU+B7wGF6B+q6qb6oBvGNJq0C62ECubwIJ
6jiqibKHYwi8bdhV9SblhkEaIMcaeY7FQ7h8CdPQTWyiPpQKOwlZ9KL0S2MTuyuSBvjbH/E47SXL
TTwrTa1U7XnB2Mr6AIWaQKihqJIr3QWa5nQD4IDi7zu3i+89bqEbqBO+xJk7VOgcyv8f3meNy9kX
GGkNgtYSdiBGrbOhZpNcpW8YtDdSZGrqCVNCmGt4+RZSyaIZD7yOH7M0dExMqcJwvIcPpzpSqR4r
zn3eUjQnkHgmIf1gobz/sj0oqOWZST/BlSMF8Z+6rsb1hAvUZaLE8N/FoghPvHFEpEdmU04nX0kN
OA/BzLxO5g0HY5S8cExArP8AadC9ktrpdFCQQdTeEqcbSfnQLRvp+9mHpooS2r88lCArN+KCe2cw
1dhlNCFASRG/XFZvyewlpFVHcgZG5lA89uQDXy9fOCoFfiGFogVcTaSmERlXSOCCmf6iIsYNdiWb
zgO9PLhEVPpu4HuakY8xeJtOu/+0YtLbsTTc41mfgj00PFBqH8ThZzpECSaBy4jbO3VMP1+VBo/E
KOBKljilZ9UZM+GVOLciUpPoVb0nUlCm08yDJBmXckcIdMZWJu2mdkjig16jfTQ9oTtmXOMttS/h
aRAn+q7BanAkst9eo9Wc+71ixH0WlUpPB2a9GeF/jonmBNalUSZ1MwFiTlNHol1QyNjxh+CXPzbQ
ChVpE/UhZUfuKsreMeDhSxoaEAeUD+Q+KSQMaA/73G+JC821dBpNwx0htHooDP/UprH3QVvUSiSl
mmEzajbecm00zkQJxXqSbrvbeV0U7pig2nE5MoJ++nrYiImDOm6mOZvi7oB6/LJMdKXvK3DBkbvT
vnGCPlnawiambAQKjvWKTAaddqkPB0bKbcyOBxnzws/Qal1Pj3m9zae2/46SoMmgm+loV9VjhcTN
D5jO2l6GQ0kagbcJuA8DZvd2rGbrMSITeXmiPODJ9jVIH8pls6a3OggyeQ3iFU6N8ELOwq9lmaQ+
D3hE0889v/2T5WWpU9V3y4v5cgAj+DQvI6vxVlKIjWxR1q9phrdVVErRGP5X6b0EOyH3dZGTeF1U
D7gteyL0WjV63DEtssWX7hAsV+7SR9yRAWP0QmB/Q8y0EyroCjS7V0+cwx+UXXeVV6QwVKuL4xLk
gdtkwH7XRjl64kzEkZtnvp607ixFR+dsTMPTJZIBThzoS62l7Qxg2wpx34NBNc6rqN8MGeh+1mMl
LO0Fd3vHSqkJSDlzIE75c2KaZXmoYXNCNcMcYaaaiae/eKNugixkZ5jdVE3Fbr8vXo2UmWDRbQgP
peHWRKC5+yNpiBjLUWsNmApfXZx/KvpEali/4UIYRm5F7UYaZBEsUuVES344yD/esSks17JFbSMZ
6keVyyvaVbY0P82MFQKwgxNpwLueIaCrqA4M3+3zBChgkdd91N7nbzcoImA5krD3A+RLNKUhLitb
7xa6hKfdrKWaB1umJ9XNwrzbZbqUbxI/2btFtnkIDt8h110/vGqTrvim81FquUcIUo8ZCA9fC6RX
TRLSjvwim4Fn5MzAT58JG25u+6CIHngHHtyY8dGEjbkE7EsbaT/UOY41/JEychbPP1IftrY8vYvV
x4fVxfE936f+6TpdVw/n7FyQneqlpzRkOnuphKAfTfXIyUvG5F5m2hJSi6x+Cbmhd8BUxVNlUEPr
x6//6DD0CpFSz9wawKIksk+NTZ5MqrL+vjk3d+wIlP2BCMLUGXes37lW7PrFe4BmNwO6A5SuIpKR
tlKPLDOO67kdF+fgAyJKprP7PPSuUfE9t/7gYU62aSqyA5hzss360I6VL+UPmR15bDkAZuKJgq3o
6cgHl+Pa/Npb13CNHWmVEiYKp58mRwQG4ILfL5jV9o5PhKZVEkN/HI21MUCgX/6WNfTCSBoRGtPi
63OBNOMZLiSNm8YkvArbYy5UZcmGc4XDDiLUdU/iN9C5U+YTCnyMkqBUap4dWOdXzlQPeAb+kEki
yOpgD5GCD654dhqyeum2o/B1zTEsTHYxFluLOFC95ehrUUstYffuRp1uetcT9KdFk6qUQAsRNtuh
Gx3kafSJ+3sqaAHbbQCA0EUAbmaj3OP1YZ9ShQ87dHpUI0TcHYP475+KVYq/zyzU9ZOGBQxL4bjS
KNEHhCm2RALvI7UoABdL2px67guFHVf6k62N/P4fxhJoqTuX/VhFOh7D/yUBjso3qHtAQykdd79b
sDZANxM4LIhopDIpr/wiEOe2P9xshIA8ZM7lKkNk82UMXECUjVT8FebN+vXQBzofdMp7RjZOBbFj
Dt8xG4bdzgiwnc3291dflbCplrZXewov++4gy3/HBQKaK0QAyIhfFucF6c3M9wkAyQkwDkfpwwn+
EmwJZX4l25PjhpFDUYQavP8/5kvhNVd3eHw3SU1GVEjPAfvr3jRdN2G+BIeoygpVAk1q3q6l1RT0
M2MOJRd9opnkm1HjfVr5td8XufVsnJgbarNBOOpkTD4m/rIJFJSPg6CcZZx++uErj0GHfU/n4vvQ
yVj5B1l/J9wXa61P1VwFZQw/m8X/KYmIoGQanlLG3R4pr9g3wgVa6czyaDWfS1Tn/mTY699LnI+B
IW+2b4Alq8U1sTOFlETW7gJgUWG+ZuRhzt4hWbiHjpkUfT5Q9LKHjy/P1aZpsUDLouuren/aTbEi
oZLhx+cMK9xWQR/Aqu9nVCPid0iMhNZyxtv7SSpzJmQdPP9hY3SAp/D0cocoGjJPMZjdtBpcmqE1
r/b60/RPdGeHpOwl+X/1LjI2oZFCyXR9/eRrZWHgfF9cbBHS4K/tOT/vfcviuSMsSNV+X0or2unL
2s3Y/9n7NXX1OuopF6fgiuSkoEpiSmZurF2AodIf67EZJXJAaDutvoY250PJnGjJGOU691zxoTvw
rjJWTpJtRwaGGjT3fo2s7bB1LfsT2yFzSnRJp+5pvCu4HSEK/3mNFNmTBp7TGf6bHI7SVeMmuKqt
kv2fJj6P4JiZRwwLF/I19YCEPT1XoqhBscHsrT1nIYiOnnbkAzaKBsTfqUmP61FMrDyFqLdkG6gu
zGYAESfM0v51PJItNnYt6mmlEx9aYrZSbFsNeGErpWY16PxlT8ksWmsMn3sX7ggnHbntWPu3uFDF
oG7FJnQ+qbahYdj7DRsiT3HWbVSo1OxliJpQi+rwx4Bu5yVQiiS8WlF5zLtyvOtIslJg6iugDMuj
XWucegEBP+mbcUEjM4OMtXMVsVDOunFfCbnNZ6H21fpeuzVvl7hfQ4FuPNJr8OOSDOAMZ6+SES4d
OoZjz+YOQwRB2M9EjOwklMr5tidOTc2r8NbxKxLC9NvLyj7bLCF+ltx43TDJKKp4Ap4Jc5PbA9iN
G7Z20gEDGiPuyYctwYZ5s20BDlXVtpf3oxgiX8H/MKujOX3rOUbvuSX8hmuKfhzPFZXZMlzyqXiP
54CcqkkSz/iv9IE0sp9sTNFn6V3sHKO4xpky32i1+pnOtcd//7+DRSID0KdRZTV2E5xh0NRXTiMp
+I3x6HVhoiLpGoG7S8Tg7vPKHyWLjWOiYj/jR9sJZXeeYf8UZKC4ojkOvjQCBPZ0W/S5kZMlyCZ3
IuM8eyQLcpUyU0ngUfUTHt4ySQjvcQtDMpY7xrE9tK8CcBD8ow8SGnOczt/xSc5Q2doVuxTTZUcf
sdmX1lT7/Cy81CydARiuWIlQ8VD22LeJcG5jZ/JTQP+nR2naJPDPS7OwSaI+bPgxMFL1Pj40GEwm
SLUFsp29hHlmbHZniDaZahNWEHYV6PRBtIgdAXKMW6h7eWSAD11340VaWs3FPrMsHgr9oDgX6qdj
YqFIZ2lR69lPYAWNtbZLyUVoQEdGaHDMHUV6vma7fkdPJCAvJetaocK87ZjM7uY8r3AQlgm/tZjb
aMIKOnWyYz5rla30KGetbCrsi/KphEcrqetO2P333cqtowS+EYVY3damETzNOvD+lXUiLzmvjYo1
1oFh2QorAicQchSPghs1NI+zbR4nTADsuFttlI/rtuA3cSUPwXi4qV022kXn1YDLzbAPhvv2MdQ7
KSA/BYaudy9bOBHZ96O7iIcYa02XcFxc1Dnua8TyWjGJyIUosYGY28SG5k383xVlAm6iTg1Q2mQk
d7PKSpJR6CEunxgU2uUtz4upTXzpT7FYYZu7xBF25WfhgvTecPtzkWx3feowKD2x+aJ9fNuF8yqR
oM52uYHu4jEQ1O0oVldoYwPMMRK2hkKsxnMCpQI+eaa9A8IR8Uo9VvbT7OFYOOoZf/p59s+MUeZ/
fjcxDdPq4rGO0zZ4FhskhA2q4LIWNPI7XIZRDAr8KgQY/fXZtGAkplPNgea44OpMPCnpT+ma8S8S
24revsZu+yhGSSgN7YzaJuI0Zzm6HawT5N+xy4a0WHhlFQhMRRi3SZYOf4WSHrY9ewMC+CxfHwyZ
i0OnzLx7U2TRZTA+jpjNydECx+bepxMFfZPKd8tORVPZUVmaYJNhHbrvp31MmaUMp/Dbw0q7raFS
L9T03pxDd896o7mWEUOKeNyDdKQrhlpOueY6q6aMMO4mUVBcnvGquI8/eRys4P9WzmJcfEw1Va7K
s+uDbOkcPwyYsL1fvbI7s8josZAVlS3c5cWninFUvoyGMXr1KI6eD7Q/N/2EYbFFqhPC1c8iuYmx
4ga/z49xVTySCphIR2treYsp00KXf89XiMbLuq+Joh6OOHtI2Kg/9kJpwEog2s/aLRC70KpLjCvD
GJtGB6RDfPX4BIsClL4KdR6JJXLTK1N9ThbKJweCz4tBAALzDDIIhuGQZDeM2dlM22EylaVdBDel
+BhTIhCV2X6K8igTGp2osXVbXwlRip1BptCZUWBMqU3/+Xrn+f26OdORQy0sh/0ffoixODA0BiVs
6ibawGbnCSOq71F3laM4tN6WWYsJrFhVlvuDhyH9z/6xuMHcnv/o078Ukmxtw/MLCbVVFLQ4vCjO
c5Duv/ELsbWglfeaz7ai0nWUHlyEfcwsZkasHowsBfGv39b0e27tMXX7Hma5tVGrp3ppBpXy8EVU
xOHVwAoQtw8ss/Mle7sh3t5cZBp4ihyu/Lsx3D8FTM1rVldrB1YuRn4HGUOCHkwmH0J7RBa2doYH
utugRNJx9jfmV4rV74wZ4j8TsGr4xKE6XqgB/8geoItPpLUt31boMPQTJJRyg0bY58YG2unRM1FC
6hRI5cJObVtmAjsSVlR7blhyOCsE0W1ZDmOg+owdF50/oXw4LvvLR7T+pxuDlbd1K7G4yUHXuw3P
V98nq/beiuYBlqMXaEg5E0CkVutO7QlFVKKRRB+a7MuU1fCiQ5h6JqEDPgy1rlv4oTVxBEu7/F/N
ExkAhcEPwEm2VRtIxFSr/XDuJoVpg1nzRAXeUNKtZuD6/WNWLBp2CCEnEvIhYV7n+8Qol5YO664Q
VawlIPUbNOspinxL2zrCEbc5R8ahS9UhwmJMrn0wcOY7ZQ+UUOkefbsmCh06hRO2Q84VaZBYq3sl
I/iunFxycqi7yZgchctgCpwbxrOiJHRRMY3p6HrNjD6ZEVGjbXyBQTHYYK9ecNlbFwRQm9XOyOot
cFq3GQsldAPYkTxgrjx9OQqYjFHOwaMN/bQx262BdoqLQ4Pv+4waoslnauvv3xHNXrRp8FGgZ/gi
cJ2C+SqQzLoMx/55yOFCpBf6IE/yZ1Rx+Ctm9H82wFyIXNo3uMejSQi2T+Z5eBC+Dl6z0YM5az6d
qzEzRSkIAME7zvrfvfZNcqNQT8UV6p0zjJLzDa8lb7WGYnULUXrK2+Ac1OdSGdxR1BKMKLRSj5yo
nSx6gyIheCCnaE1MSiT4BwC/1A9A63PIz+kkHT7CsNMimw5F0cEZfXZMGR6wAxiKek5RzAQDI1T9
mSuBYqV0d9zEgnOS+5Dck7sldlCpgNuWzRztw7E/OVD4fn+8nZJuwBaNY4BHlRurwmKjaLgb6LAD
Hk04ON9t1zSJiNrzXxzwmslDOxsrNAYJ0uEExChnzc7MwzqCHGU6G4gedKk0exW7EppBvjDyARnG
l0DIBrbSQUw1eGETGz6G/sb66r+eAI8klddxgPTG6xcDZpr2ugguV6MsI9hQkitytY3Ma4cmOf6b
Wuih2ahENIPe40oDLGT0FcZm0qL1NingW+kHLVSEk0YM4mWPn0X2n+/CktTh2HbrnIQLF1SKcjc+
ozly/yQbfCjoBuoYJeVpccXJ00vwiKMbLs859+ts8kdQuhQpGYJJqijhdNcnf3x8Fslz5ObvIUw1
VkW80YE+osuR61jsiAO7lgVfjWhj8xikh5MfDHaiVWKrqCBWhgDSVPUQbiPAPY9i1sHujEzxoGBr
2FywAKR6y5h10aghbLaWtm7vkk6nbEJlBicLryD5ILtV4thYv3mtxNyDH/fZ/xb256VusDpAJneP
E/KRra8dOlM1krNTzJ3Y4EHjvXsNpZhSNh3XvG+rahKvX+Z8KnLz2sRNWzu4aIiCpKOQhVOF5A/q
hdF2mSOwe2qk0l/By1CN1JZZugh8KbN04GpVQnfiQ/WMylmAxFIC957QImqemT3E07PqaFz/WU+1
A+aI6kOhiIsYsfRfgAQqBaT7YgsF2hzBaPcq0DC3zx0WxJ83mrgN+Gk+2va3XZoVYoek8eJDS/ve
+zeSApoMUotnM5pxKv5y65iPTK5IScaglNnabuQyMcGT449h6lGCX+oOT45rN33VX4bJk5ijPJ8w
sZ804priRgXBDaXO6+mooMDphqQOlv+xbJmJ77zc/lt8aAAagpVQfs1nBWhiAVVmMljbf0nq9wc/
2cSLG71Dcl+VYPsIgMiFIN7q05BE/1SlBuqoP1IhJrpyiytcGn6tsq564/OTUM0X1JRwxeNn5f7U
aJjEf7jvgtlsKjWlEgwTJPtfz1D83Dk6CcD0KMXJXiU039ZevZqQKyrmx06w87/EL+Ifk8a3GWE9
lfx9WhPR9MDm43tRMMQaqPowCliOznx16iSDLzln1TCXOD1eGB3bMt0Geu9TVynzpuvaOsZE8flu
nQgGZuppNZnHj4W21xFcId13APrS7Hi/EazSdNjEq6DKpf9GtxLHghOMBgzQB7b7mSqYMkCDAHj7
Tp2BS0cBxx+nTUuWEYUs9JUPPD2eDr3F26oE+QTfPy2jhHm13g9etppXyknSXOZW5QnNxoZcJvcd
q9jJUZMq3tMKTWQ7RYlG/W1T5TOBItDMiGB75Vu1/RZOE19ngWxt+6BDhhDz7BMh/5wAqcy8D0Z/
c+BHDWGxO3V9e4TAsBBc2re5GGWJIITiA+o0ghdV/ME5Nig3Bd/z+f307OehRZwbjr8bZ/7o5BGd
DGxlWUo8EO5I2Ed6LNgaoStKUk84nnwhj5QpkI9BHV9RcNG70xDY5aQrkt9LR74w7Mz185DjhZL3
A8TpJkea0OFJow+x8rMYkcVVagYdh07r3Sv7E5DhLQ4KKo0q4A9aBj8NRJ9Gf4DOJpd5ZCcELoui
qfMPd9V2Ps4KSGfNqALc+48O9TyjhQhw/otHhTMa04HSuq04HW/yk/ovShkcx7RyB4kWcc8AFHc2
aOl0kOjx0TU2UbfhDMFjzcM1UOWrzceSHU6d2jPHQ6ooQSiTAAwPGY6V/DOy6BpfDTCXiDxdO2hu
DtGkeTz1UGirUWwZqUijMtyfCOppgBJBb9KEIqCDVjVicQeF25sYWj6JqqgEb2yjGtAKa62hxvYR
n5BA4YvHdEKQoDdnJdilChdWtDtsSwyWGaIQVqkShGIzfOpasUkBdSHLSV9E8wjQ0ou6A7suIe0m
Tk2FPNeJyPcVhi+It9DFwdw1UvPhMb9NvDh/b5XA7F2lV7ZtV22GkK0aJbefTCtOigQ6FJq7XacN
Qh+5TQkF2aRmDKR5EOg0G76BAp/EkCBAPrIYEJrBnay+5IPwT4IgeZp4pImX5K2qI5qc7l2FmiOy
IWuNwN+AgwPtrRyz3laB+5DU5sXKCx1luLnRlhFUpLZ20unFF6tRagAWUheAOG9Q/Xj7wxhYYYFz
PLeGdastrYHwrM8xhBYMp5RvEI4Xfeh0NUQrzUAcGAZgOkBpXkB5CHs9TMPXZgcO8HRP7JKUfxGV
ngoYGXInv+ugignrENzywjC8RmGjpXNlWybENgPeUAd8C0nCbMIBOZVr5RjZPzoRYkfTDPBveypx
k/XLNJoz11qIDtIlwpsXbyUPqjt+rAo5Zl62IehKHletMWthN+aoznT4gvSCc4NqHkto5kIIV2WA
fFtyNOTuuxxvyqSLLRh73DmwuaSKRM8IbZzFx2vOb4gWSoajfLMPeV7bgzyslzeTL5RFxKEyvKNc
AnbnnWBs6ocYE1ByZTulKEMTB4PZAO25Q9PvNtF/s8GldpD6qeO1sQTdYsLCWT4tYEUY3Flad2gz
mTIPtAycykq+5v+usv04gKkW981gr/vK/IpoTRm8wO2sOcDgIO3zFF6KrdjRoVeXjVKmVN/gc+eJ
L+/N8mZZrC5xwBhDdymVn2AxX9Z65p7Ow9DwP3fyY91hDrAn1WwZov5bvwsTH15PWQQXn1J9dBd6
r0kdGiWvtJaYEafeMqQeh2BZ55IxuGgOk19ccpn6f2qoaE9RnUEJJ/UprcKKtt/q6+sD1hSItqDj
ZRQ5ZF6xtLdgPuDBCo9DLT2fCvPYP0wiWT/lpU8TzSYHj8hO/9hymRnF7ub+6vT8gOWcnHw6mRZQ
dDXZbWQYaepF/HMdRPgaHreTBzFV8vJR6OQFadeazASaFNv7Cr52W/vW8lIxgrj5lNBh1RjNUShR
NmIik78Her9dagMP4JF81DEuKS3WPxiN1Uf0kAZSu+seEqsHHP7dbJLETWuR1qzvmj8FQ/XZbzav
gQj+TppKI46CqnZzALCgFYLDWrUwDGmL8u5Z1EtcQCdFRw2itLsIZuUfYcsXJwjQL/RUMkyn3cQp
Ee8+3Y/q9LXBPhhf/PDeNQyE+/kVpaZhplcs1c4CCJS66y7oxgwfHeyqUIAYOzEoVHp7TnwmnCAI
Qc27ZwcrvYNaz1TCd7hLt93jeCdsj2056XvLBj+XVP1geMYFeQcCUBLWt8FqB0T5JrOigiFQ80BG
BxaMLmr/RYaonPe04UtFgs+WMagzolzg3Soh+QvgJ4UqmNam4vHvl/vkBaqeH/pgaEJC99y7CZrQ
uf3U3edeaUQH0BgKw4IZKdWUlX2PZeBf6s59Y0KopdtY/O4k8VYNy5kvFMyOVsj03J8eTMM01Rcg
vYigNj4ShR9TNN5efmj7YlQ4MAG7uiBCF8Tp56ReuCeBS7dWZxpZgOsHzDN7RW3QpV/2Rw77bwtj
1L4yqRKkI43ezWxjoJoAvbiB5RkcSno4nSQZ2LOGCpHJq5RWL4405qHVkLUeIpEdLWimaEYQOwN1
p9/CbjF16FVtNvSnx4Liv3ATnsr3KUYWseRNiZxfwjLoV6Yp+mAehXM1esOe+6/oZmMUIXnW0p0T
Mg3ucyq+CvRmbPJ/CaBIlGTk0HLYkqpVFNNkS1QcW/k/xia1gES20uO9th6+M3cq5Kj1U3H9R8Hs
ipk3lyFjFi8LF9ddpyoGJadk+21Pdp5PVzUrqRHwwlgqB6gEJoS3/KED+TyF5BQZ/I/LYkAnwG0p
o9fFVIdPicnUT2nJjpLarMdVj6VQA6eims3SLLcoOy8gqo19xxRt4+0LT2Efoe4JXgUPPE5/lTo3
yfxdXIfJVcLcoMBb0bfd2u5xDK80pIIzBHBzTHyCl4/tuzBoqKw/zAsjhTk+2tMNbixOC3zDwVRK
o5WlNULPVkhIWL2qdWAcu6ccmyDA7lkvAyNQJ5sZDBaO4ICmfubw+sV4/6/nRAFjTY3D9ktHeO/S
xaCyGvUCZEPCYmWJLLsAFK7O0qX8bYU5J39JHDQY6lVBzmnMycOcTKFJ/J563MmAP33LRaCIlX7E
yeLHOWcNOuGDISlBYsksfN0mUMSUV+xCO9ANKRKv/9XTbw/ZBvXk0SscjRJMzqx1SzQ90d2FIrTE
+wXryw7TBd5s+ETnYQRnhz+XVRFsIpFRD1rCbkr+AMfOEd0u5OECa+yXWWVKMRu+n/cSsOi3vLHe
BW+IEbnrpPGEtiR5/gsmGIMqsI48ZU0WtyA8+zT7/U1objwQUS2jbfpofcoPV6tKuNrashWFDVwG
2Ai9KQeF4V99Hhqb4WPaYNB56gQdpR40T9tBgIyKeH097y0GH2awf8AQ4lvgPJSIMvKQaTZq4V65
id7DdMSJtO6nuLaC80UikK31I7R41sc26JKAtVT6Fr3jEaIFHSBmTDBMB2wzrIfciw4DbG69VLvM
e3WG0dKupaJSAqetXMBi7Sm5SzuLpGBPYbdhZkJ6R0q/Mn8/IuDoFXUVqdGPuDGftkX+XzbSry7L
JJKXywNs0n06pTr3LvDDLz3Bl9TRdHHMC19xqFibRkGsWvALRqHhpVSQkRwx7x3sGWpo70IosYRt
UxODtWkT+R27Jah8yzvW4oXYpXZYDJxdJ19xrzeILnxtBhx3Km3uDvOV9iLytzD6Ju9xxYmxR3WI
fIdxZb1i+Q/PHMDnAy333TZlu3QMt7H8cAcYkFHbGquKbYLoYujDgi8gEt5HOtnyC9r/9pRqv48F
KL06pLsxColt/4hhW+7iJUKtp0Woy+NnklDOq4JM2f6lgZLCJnlfD3+b7VQomCg/bGPV9x9krxn8
XEO0tfw+y8Rk+KH1XP5DtAnPjZCD2Dl1Kuf3rwrs+mQ6sNWKXnESgOyrtOrt33PiXxEBHT2Fm2Lp
ycjAi68Xb9O4Pl2YfQCT1B5Tu4AfGq2c+/oA9D3bp+mNjYcDTDC7H2J75U7x3knH3ofbrra/yxRF
cRNBV3u0wFJssL1BrvWRqlmXOFWkX3rNh6/zK/pI/mCGriMejy6wik7ovAzq6aiqd//4yr/lOqEq
204K0ViAXtNrllVS2SdS5uAWuZrvj/tjRgVjjuIJe7krYKnxTrlJLgFUyqFNEvLRBe+fn00UiWmm
vKWdc6QkWf8WJrTd89ofbpv+pIremmFYLikLJwB7wo8Np6nCKv2bBb4ECU5Hl/oqtPA9Lwib49i8
2JFOg93A1GK/xD/WmMsf+1XRO/Csb/AZns5KjXOJVmqxOUdg1eizlhQpWD8CMHBAMlgHzachZB6C
O311QLC2w0XtmEOSCTumMpKw34eTIYTszPU/yiOhdoymgI530ntqJAP0mSUYnVVf0F0OLtM5BLw7
HjFEd7FF3r2Hs96LFqiPEL43lTq8bvNYmM8IIipFIvjglfFc3l/H8VXP5YR8k95w1rwjc76pY/zy
fvYKys5/Sn4bKRo2sznm7vU4MaTh3woRk3f/oZ9RDmen8ZpvNHHwtPkBwacemvPU+Aqjt8y5a6dz
8kXlugJN3q20IInOOuG3P4ApVaWCPrO8hhRG+tqYQetzJgOvtDXiW3lx0J98BRw5KxV219BgwiQA
fq4U6S56QQI+PmnbTVSqOkwtGr+xEHehj/1Q86N1mJL5ECDlKForcO5BzOFkQ4lRHYLV7T+gyy8c
nOOi6hq6W7HsencsnWrVUa+MtXMofIku8INEjwHIpYTQgfitX13yrL8e/yD9O7ZYLrzUkND4omSg
4upR40C58Jc7habSnDqUuvj41d71AvQDUBUk7D4l3iMpnFnZRcBBjeEQWoQVO+Gviq5U6t/oMyKf
cXhxlOjA4T6+nZKjxlQ07dIb04G8OyeuRhrcyCu1l+4yc0/Z/ZWeE5D6dJJljxasTMiT8NyqA7g1
+d17xJC9Lz+vg1mUF/kZua0kEC3Im8H4FaGVyxgzLaAu8BNJesRfpkIPJnSiO7Ye4hgwaTj4qDxG
aZqTk6+PEWtcPQVT80DooJlA2qTe4S67ga22qO0DBkuKt1YQ0Rn2IfuLInypE9fRMCsKPNF9zFpH
IG4uF4fWxFlrNi8tW93S8yUDPFG6oUPlzTX5xR1BuD8vKgivlYbkmfIckvAGePZ5JYw3vDPXHsUU
tw+ai/u9yrLd6gyVARfgMH15RaewvdawyRBJ45c5lwoAWqpftiCfA7ebtt9zuqNXfJMy5qEQPQE6
6hZe7yGELjpLY/cT6Q+r/gtMQ5BOGy6/MVNuf0IQLx1XESRsWP41tCrG/+Pu5TW/d8U5vYG84Wa4
Bmj75wgcdx355YUyvkvlCRPAGQQpRiSx68rDzuTqNOt10u91Odm/cVw2pzSFVnCVEg63djdDS/1n
TVHlDwF0RDLU/EzjigTF0i3HGf/eWbB/FbWCa5AYv0tqEKnOFMx0oLUD1imr/S6ZQqPgldMjK2j8
PyOdyaMgmzm+LH6sYQs2pR8xkS8ACb7JSuxyEzvp3rKo4See7FJEykwVqy5slQE1AFZk8cVLGohg
X6lGAa0nRTAMWHQIqBQkNYJaJ+EjpusPffqNxa+wrbwkV2/DBsOGE3XPszqZe34lI+aHM03CCt48
/0VPKx5GJVtgjHE4Rr22z/5YznWJhXxim+ZYtMN3PWhd+YA37CkDvyTE6eq/ndg9a8YBg5Zu8s3O
yxqd1qeHANa1NOUQUtv82/JBupfP+qXYQ3og7mOkDnE2eHvlkizw8t9Yy2wks/JXeO5Z9OiKCrGM
7E8VgqySpyMdDqjTmaR4ylNSbscATbTO9UdfVhKJsIaKPHgPCr5pSN+7S43Du9hwz6zxeWKH1DF7
Y88WH9ps79ZEI8Tqi4EF45i54VO1U933w4EFebjsoJGiGTrzW95ucKbUUwqq7exT8I7PnELVMqe1
ZNGXqZ7jDDaoG0gHFedKNgdM62VljKeARmA8ON1jhTHySS94ntRAi6532OoA6qFynLzo0sggyidB
bvroo9amBPzl/QFs8gK5ITWSnvvWdprnyvzGtY/6ibwz0N9bnwnLyRIJl+lO5ICcK6s9WxFAWMCL
CXc+LVeYcsx+Uj91hGgznamJol+ua36Okyn68nlhT2typaQNRmpO+CQKXHddzKwsjfmYExiS2eko
x7jHz5BdeFb+0wzrEI5DX55UgoGHOY86hUHF+8+rcNg3gk6wo4i5/dUgsJ2GIsXGAKR2QR9ergeH
d0nExXW0XxXZzOfGsirayLpOO5KE7jVEwBnyY70NOl2bHGkvMpWxTp4wBwG7UB5ITWgpjucn8QSM
9eP/BdLy8dNlqHtLRmLyNJ5z6kESnN7XamfpNaMg9mE/8BWRVxnsCNUA0RI3xCb6o8GfX5AMjMPo
AMvmt1Clj9EvxJ1pEBQb791A8HXiw7ANd2uZujd0uaQzb8GtLv9IbEUQP+DG1O/3FNP7J+5IDKSb
VDO8yAKYfB7EJ8OYcxdCiaqePobin8KeWBhD/XmzMTUUUWcqH4eYsBPqGeGkctvcpUTzeJYzBTOc
so3zIiTpWEvNi7GCktHm4eojPDxeytySLLplHxS89Q4Wai5goAshLWtMaXKtjDNzR0dcH+xlZjio
W6ij9zXcJC5OBj95Eq8X1C+KyK1/SLqIhXcr43xKZEAtvLCGLI8+5EnFhqC6OHA8ws3kc5BG01Kq
5/qEUi3F//iDac2Ph+NsSfREAYdngFxb5TkWJFNlQ0WYXdBodAm3dYhYQURzr8r3bL7dkDXT1Fy9
ypWFIpY2scDe5BaO/UvLoMOnSrzrBZ2+MyN/L0CAht/pF7TfTjTgOEQrgF/BXeE/h4zJornwFjAU
Torpt7l6uSBH4QSiP45DRneAzAEsNyPDk23QI0kLolm2rVcsDeoXUdRxbM5f99kFU4zpPAVghLk0
AsSSMSTlCZJGkyl8i3ofMGCqsWoGteOh1LHp5eDDdEVhDnbUnF1OEPhATvKs8BByCwrdm9k6wfMj
daboQmUAd1a8YEUfjhIZCSNwcTRjxidy+TvFNnXp+CT/65t40Zy0X1q8+PhIRzgHDMlW+6OrPcto
5b8nRCmulLPgNyaIObIanEWVWt8QIP21Ip2XzXjogTfTFTfr61/DiQ63JpGG6jTEUa757EidFZDM
fr/RD44SbJCWsmf6xamG76qrkLSJZFPv5bMFO2zp37pQJQD3Zqf/+pnmI82EAPk8z2VICdUvxfui
YTtscPb4cyBuls6pajsIsfNbIlsVTrug10ZAAahBXuDYW981uAI3NNRDNKBZyI4zIONNLKCM+APv
Az9RjYYBRCWp5xnFLczVpUULwhvLBlNFiyizQ8VDdAYlPGDPfQvpBcYPDbhUi2Qx5A/UpsqWdO5u
0wT7DnwqvsZBFAPV3A+NBoufUrYjWReRYJR9N52QTbTLAyt76CDW6MNEyxEF73ORs/aUOmsC0keI
u3rLBRi+NVUdkKNTTGlkcoLB4+lJqh5y+AEiijCDEi9WsOcKktvbBkgDezTJIefmL8/QSXGgaJv9
WSAEElHNBzZB8DaLruz5lgG/cpO0G1+MVTKdHToF5eQxBAalUda/mWrj8dJ9uvvvtH7P+fpIixXU
6zi/0GU7ouN6r6YUnzZB8DrpEYaHP5tdxeaRU2HmjY7BRrogvZJqjMD9RmAIwR+F8RH6l59O9vKk
sfdZVSlcVcSbHeh3dN6Ctt4prYUIU24M6ozg0JjJEohjPUPEyPcLGemPIx78qAT7NfMONReaI0kK
WSzjSzVZjHmIV56c3PtTWQ4xXDMtxepG0pMdRXg9bVuB37PlU2CU60scCmnsXlvVjOcCyUg9o/Cd
Ey4RbpXPbloQsG5uE6Gb6zEXexe3rW4VOy8sqOTeh9O3xl8x9UBI09g4tXjFHjfVqlAihQ9JfJ4G
Kd9in/UgLJCehdoDdXpNiUTCJxmqRjjdGtGEDrZd+oXkmaVRaqjN0InT9k7EpVzm0qjmUO467wBi
yjvWQZtephKk1SEg0DD+A4+R35GPnWn8rGaJXoqYbdhZtCCWKVLFpMpqAJ3heudRO5iAUoCLJAur
sMhVfii/KFvgM3SBt6rszg83sqtDuIEcRzEOSpphYskVz0TQMkKCxwojDouR8lfkvC39B+sJulkw
U4NNO4g8mTl9BW002RroSPjvqT4PAD0Ge2wArWlWhUrHOamdl7NCFZ4c9C1nAdGWDGkyqU7i9deK
G1iWqAPQMQ3l+vo4E0evrSoWukGfSOGgBual4/S6sOxlCxIp6paKTK/FZJr4+EbxmxHTHYN76EFv
mERIYaiw5Sx7bmIlvmaB7RG2QeSe/w2wSlhJ19fqv+nns/2D0vHk0FWLCVC5BrqGTSzGhMjxF1qd
x8smifeu2kNusH0X4BhSSLlTx8xGS5++Jv1CV54Z7Hs9ngPRi5pKl9jSXno3yw/ow7eHLQ38wIR5
adlHScaWQULRt3UAczZhJy2qmoxpkQzEpZ+gMQaxfiRbBzrs3zzFwikqt3D5cKxv4fXgMLiZK+ki
khTWGaMLkgPpvXcRZWZ+K6jS57iYUa5k+ZbOpRjUXFeRrvPpAl8UF0aOk5oIIs926p5czVFoEA0q
4/cIKMdwNDC+M2UHtwsHsXHZ3YmlwZilrmyRCyH7V5xBRDz7aAi+4qr4uFAlEARMuzDcuazPK/nk
vyV0tVI7K5zgUDvGda2kbNoMNz7fVMyiBx5XA93gddntJDBL2NdlUcmM0s/K22a1dccQ6Vu/nVaH
nCA+jMqCHO+gq+gaMb5Mjisfq/bsPPvR1dxAg7tbs63qcWAL6rvyL9/Ax4/wq2rf7+nlN7J4aYVh
Kcb2gOxbiCa5F72H40ywg7vxyQVlqWNKMMzKyon313nxo8wzX423J6eKLwGD8fVhbfGRf8npk3Df
BVn98lIOnqFNnz5cDIIvun0aVC2wgok51mSmvH57prMOak2YoMh6qAEyhQAc7IPOVtcuJABjZ37t
dDVO7OaTL0XkvtyZbjLSugZty9JV5bec2cf3mCI/rx4NZW9CPyqY8b/3r9hl1k61uNFADkOrQXQX
hhE9mWL6sv2d+ffw9vpK/QW85a/TWqZI6dgr4ny2EILhturZpPNkJiefMPxVnD3VnDAcglMfIAJ3
Caah5cW5PDZOCmZ12TsLdPsuxDEZzOlN8ub3mEp9NS+E3mWrmy4RSlukaRSqIYQ9if25Z8ZRSsjx
lSboxjA3Vdc2ENmSUZMvZZqpj51wqsI7Kzg7fjs4d/IKYnt/gD/gXdYEhrH+9om0UBPtJYkBtieq
84DCEu59w31l47S02zdyQr559BUb3mT/2KFl5HKxSnZ/n4h2g6L59ENHj2S12LLatVBVy5I8gSB1
rbbjj2QJzMNGUrRSswKc0ms67QLSZbA4RLDfeMcbCh+XJvSTXDrMWjtFg9FOQnj+s02haMz1yz/q
JE3ohArPCY80Ktz0IHBMgKe7KonK+6BKMAzYbWTO4HsXpopoOOwr/TtLCrQ2ya0DipcU5CZ6jFqS
jLNPr7OlGSzh6GXUryOqkkDv7aAjZigqEljA9j44kp5lyw1sacA/zkuC+UgXYsST3GCk7bQJ7OBm
A74SnQRMbaWX9bv94n1J761sTaBRnW7MnNpTgHbuDYGyQ/9p8rOZCfwQ1rck/0yfpRC7a4KuEPSI
b5I7ZfJxBbXSEUn+41fr9JvIaAGkoLnjqWXaf6CsE1578A8DxskV6TzVqBFyayda0BHEH6V1OMEH
imWklfo6+JJT+NbPn/Flt/ztp5LuE50cgxWn0H3R+ch1n9K0Ph9/3UCw8ZnMbZVD8dVmGYl6dzWb
uw/+xgXxdMGoG0SXRaTQMRMe/yGipgDkSFTjTaMKHQRxqCstdmry0Y7Se5KWZ+7h46Edq575TZPZ
F65S6C9SeWWfN2YshKYnu0M+G2CVsH5VB09Opwqc5yMuodLqrVbBkhoJUiaoa9UeRGMywl/mfVoe
waBlAG5jXMfbKngHcePu39o3ZNhBdIKbh4TJs7vLbWvxV7spsiMd9G0NWKiLiZ9gEsoiX2hTCEbn
bjq/zaCucRQBFtPN+liFK8zxX/Af5WT1xJ0jCbvjXR/mMetWrsAUst7OdaRsJ7h5fcN4iaK9bbZ4
FXbajtPTSodKOOb5gYD/Dr1B02s3hv3rdCOsR05BQoACDMGLVv46u1gcBB6tsohg9EC4Y0jf1my4
JI1Sj811UEm1oLZld0Ercgd5J1GvSXyVuuE4AgmlQfkQhy3PwJch2tH4rl/Uo7Wzq+Gbluau9W5l
8ft1QzbNCk76vF6YXwZSsJuJADDX2jfutDb1AwEtkwTElUMrxprfqzZB+qjxG0iB7YvK2i7Kg09V
8yEe7sejEPyRhat4NMMarz40dD10rjv2z8LBj0Fqs5jfgNIa7VEKMq/2MB8emrBZ4E/EktMcJ2qN
4zXf3Ad6o3EWihP16K85ZqWYdzau0Z7oWzaPIN2yZTI5R36FR7ro1qUJOHAWtwvvDJBoK32+/a4k
Yet9csvme/48i3OJVXTb6nAPoRJ6Wdto9L5e2LliQSuWiFrhblcdLsUz0w24mLloUIHuyhT5n5I4
byZDk1L3d4VgIMxIxkZ1EmBhiED+eUvDQVNinIm0MW7/0NCESAs91oFORcQLBmOIg59vuL5udZ/D
AlhKo7QCv/t5MesYMGoFp1GGFBhSVH1BxVy+URQutdgrp/vICpf4H0gUu6+laNgUl5xmUx6+w7yl
ZHfQCvVOBpRXKEhq47wgHwrO+QKqmcpyFz/N2Ub69l5e2XXwSzF62DYfEjD/Us0mcw06CHM77r3L
O1ggIMCUSN9TCWQu5E6TZVGvN4Q6NW6Yn1TIw9XqnP5LazcZ8dSeKadys4jjOaZesUh17MVZ8PSH
AQhVTL51mhPqEbWNk0fOjm0D3M5HKE2P5RYJEXGevGnHnD8Xwf18IcckPwXzAwkmLCb6EGp/VU8V
lZxQjn6OFXRMUhsh887PGhFOfOAhc1RmX6cAH32FTinDtNE8mRrvahq/vz3A/krnnLk1tn/Uaouh
nL9JXFvgzRGmqSLyUlg2poJ7HSJkYaKfqco+HJJwW3lE7pTR7j0t0imOd09Iy2P0z5xyXniRO5BC
4ZllvUvvqmx9AZTZHyYcnmjQ9/XM/kDZwqN2n3ldBmGTObhHY479sXOqvcU4/JV7l/Vqdk3yrrGo
q/PdLzLNZUpeAFQnvGKNXsGR53/cmfkqSxulBk+SvLQCUP9u7X1kFtal7q3Yp/5qEqk3ajWLqBt2
S2ZCaQEbhXnbORuqiSsaEnSEAQkGd0T2vTfhr5mdlPW0OWY8dAiflPozOidxZb97xYLj+NkvDma8
PmSIYehzAz/v0kBod9bTgLsTq7Fz/9nmfHC3ZXPaseP6zuUQ4nRL3hnLI7ivX/tl/ZItoBLUH1+T
JSEedgcI2Prm98ZzcuqZmlYjKznHmakQ8sxg6QaA2oFBIL3bNn2uPN3p42Bko7Dtwkfh4FXW0dKX
/oSMnycKRQS6pyFtblgT/UW09bCyl3xsqm0GMejyVg70+YLM2H6SbAfDoLE1PTu8bWTx1d2MQWMT
xluFrSZA4s8Fjq+dGa4dqJSiOJt0ubKngiwk3tmgE8L3Xjqf+P7T7Qc0k5T2IiX/fW/UF8h5L9t3
DOS62+Rj6BNtmJb/rem1h3tTBl3QVxtlwRKO/00cY0LUvfzrdgHEGC3ornafnjqNJvOrAR/gwOlG
ds7ei+cMrg8JquBYb7xYs5Mz7M7UPgEdBwJNdqW0Ckovl5pRgUPPzyl7CTkdIfqTCgUxgneDTucX
WogkB3GCIgGshc15QSvW6g2DgPoOSWRSqz9ZW2yM0LRANUax8FbC/jgxPqu5tlsR47bVf/c5huKf
kMO74XenzrfCtqpFvttihYTYMPDdre0bRbaDgPa7zloCzurk6yzdpJpW/wVTVfpeBDVV7HRJX6Gf
Ft8SVRH+7JZrXe24BJ2JNTefjC66E6wtRuG49eHdOm44SnTV//BssIoV8t6NMBK8ZRBeB9yEq6Ct
jhgv8L6iqOIVQw3CepD49wY6FuRAVErH5sds/9ZcOwMmsspXC/paU1BWFCyX4cJLD/xD7wHppisI
YYnvsY7nmQILi0i9Ux1VkDhX61FnOL5uiB7y4sXvckf7mh46+Sj1DAiZlt/puF/4XQzQI8fNwQSG
xH/R+h2HoT8MWUTC7Vchb/A87/uhue42dJBX4TOJ2urEch91dM8Fe2N+8N/oFsaSxWViwB1TJGNf
YE0/m+rnQ1JHgaeVeuk0hlwtrEX1FMxsXLuz+6L2vmvMTkWOmWmGaDvR3nmDYyhbqPUIc9245txp
qJGszCq/iKBypeNplPjw7TbVlQpp83scoG2uINngYt9Kfj8Fo37D/geYCHgi66LJRtpkyoU1Dija
Ea9/0hU7vkkD+Yq2SrWwFDtRQFIJz0cVKRbb9ffbwwefZezgBnV96k6bpwVir+xC7a8S4aPzpeuq
ZyfqOI2Pdv/60Qbfq5Iz+chDXX481SF6HAeoH4/ztHpzLlX4tKXd41QfxFKF6qVAy3Y4otOTXvO9
sf4fZCOzkhMW4d6JGwtP8LmeWEOdFIE/x5GzwDUdoNm9ejtZmddOc1xb4qmONAEqoZHH4OrXoo8d
I0YRjCBJK3WQ/JNFntK/v8U582PrHysjal+9SU/iB+FM6Ma3RNCawdAZ7NqXxTlvw5VT816bWGiz
lEFP3Zn+uyRpbUx3LFnLD5++nReE8l+A8A7gUl+ByT5ImgvNMb7Q4wYysRS1RH3ouhci4rrN6znS
UGI9QXZjOj0/SAz2bR8ItjVPTaeQb2QpfzA9LeFPNzNQpYxIxeDW0aT/UdSLcKzKfp3LExBJXtuE
YmkcwvLIAfcJ8PgDG4B3IDFGwqhZh88Uv5Rst9YB/pWFmANSrGcpTR+IrNWA8IGkSimtbGS+U2Pg
f+6d4BxLF64FI6LUsXFVrc2rCoTV+63LOy5CFKOdMdXkCM4eFlrkeUk0SJNWajDrWeHwv04Rkncd
7lFDDTEPzvkyQlEYqaWVfHc/yGx3ze0Z9EJCyOEjwWDGoAE1de6qovBg8fTKH2j/4kTg7dAfRdD2
7NwZOMcz5H+4spANJvKc8bgZ5RyEW+h393fHp8ihcxd7MO/UASPMFjcH49Kle7hC5pZdBItNgnSP
zi5bLhY9BdC9Q0LJLj7tTshjv9ezM5yMA5VggITRSB6mV5kOPmKdmW9NVcky8riY8yCwv5f+71Du
yxJHYtKNtuqR0pmU7Kb7f0bcVwgSNq1VLo5NpNNNc5RYCb5nf5A9wTV/CHWbcarCNwD8vXPB3DKR
5WBA6Ll5JNNrySbLihlLI/7hjU+z5Efj0wwf7yax2ld4GZHgD1qu4TYgNuyj9WFaEqOV6thh0jcm
ZZ0fergRtdWoEabIVXx8V09JGOIvr44/F1Ugrk1GNHOJbaIxWVaVzXDesBgMrjSskzCJaihP+KAV
civRtlMoIy9fjSh2GV9N0+0zVxGQ5q+AjqyqLLjr4u3W99jvECZuDNLbnf4e4Bm8taPOpwhYaGZ3
cHFaqLKKPm1qcMCuwQUtNwCdkDF44NSZ9w201jnh/EAgyCfWYjpvLR4RKg8ecAlnzkcBWXyr1q2q
FXdODrAcEL77ZQK8YBm5FHXYPQe+cKtZq/RgUvY6t2SOe4DwXtgC0tNx46co5YtNBFZKWTh4MLeI
XR/0plNhitTl3l2CNejPf+/+PB/UfDzPzSTJKmazcwrjJbqqs7oAU9cwBeeig+/uh6LFnt3gTHIp
BbHpHLnQRrk2cW1HuAgdFVMQGRBf4Vy70RUafzfvLztjXJ0/bonrJAUfdz+7mvThQJQ+0QH25C9C
08SmGB+qrXlssu0xS6NIbRHb10jRCGuJXkFhjQbbm3vx+rp9GqkHxZhcH+vfTprbZ37vT1z7JMkH
kTDq+Krypev8wpGUpQI6gxEs7hu+ZXo4nE0jSy/NpMVgd1StLNMUh8Duq1A1CGlv0CTdtj6GgHrM
AIHIYOJBOoN2fc6jc+qnRYhMKTLYUAY7GiblHpFS/46+NtHuRrX8EOOAsFLOGnGEb0MsKAPQ7Odi
EakhBxjIGo/dRgxbBCD8QDnOixZxPVKvQ1Tc5OJMjo/LJttEpBRaUixAIng6AuD5Usaun+bkT1Sv
7qFmPh20CV1AJJc1Oc2B5q94pBHJSzYTBvRJRKKpvB56gja8hf8h7+qRrq9xAkDEdUXBnJwWvMKK
NV5OKIBxWRiM8UEp2bjqbGZW7eAmt977x23Sl02M5cgtc0INJPO92hANEBCzbScOHxS8f4iKo7KU
yIXQE92Eju28Gmg0v/ILjppmLpSO4CMV3pAOPGTfjHd0tNpT0+kQpNcWZMRj6WOo8au/MSJnRWGB
WZCpK5wfYCb16EAqvPi7JLiWGKsxTwu/vAGKd3//+7dMwDgM6GfHTzUUZL3PjHxFj8XCZlD1JH59
Z83BXSaIMoHTCeEVqioP7SAzfCwtziqOozlgHfLQHCTalwAZ8dyvIOhofsSGqej4PpMq/X6KyuBw
hFCznBTxK+A/0My+3dxLzi96WiVTZ0Qppv4K1cJ9RZUFwBXkPReiLGk/K9R5x09I3m3aZlVxMIhc
PuVdm+d8Be9eDl8HhiQRM0XfaN6PSQoInMB3dfvQ5pPjEoX2wwgi3ZJz7iYy1Q14N8+6hIUzH/5f
o9Qym6uWsv95tdFn2SzozYGYkUT0WZujklMHAB2zN+y1P+ZjI0ZdR3sZxeaSXqOR+hBhTIqYWfhj
6j1lSDzA/A/UJqCNFGLU3bt4KpXkLalUuokiXbyZjTE3++YrsR9qwhnRLkUhCcW/MbZNW8Bgj9JJ
j+82qk1lwNS8aSa1n3dGLxxz3Lcbne735IzexgGr1uz73DkmePk8h2VaBqp83hf2JYe5JF0MKqHb
lxUUOKQ66oWNkZnhYkJqV3itH9ASz0XIkIqW3fLnUVRe5LVKRcNklIvbK6FOUO2cq+T075GSs+UQ
8sUDnyxCcUQwYuEW2+uqc7ohE0hWO74MnC3Gs7Jlr2o0hxsxN9NQaAmESBOtExkZAXhXpIyyvDOk
d1i1kTcg2KU9ozfT6325yVH8uMoOWAajDiiTMLZRWjnQopm9pxkIqxeHs4NhUalkyLliIK417llQ
iBpMeSu+6nXKOu28XvHIjxggakhdUdlUSZsiAV3v32ApVHhVTEvmpKKX/vGpEWAvXpj0xNbnGtoM
4SuWESoQuJKfr+TPjYGlPfuqViBXtzMBgFG/i26wq9twoWqv8BA7sZO6qsCDs17fx9oQI+vMTAhT
11QsOaJ0x6AwwLLNzD0jmy4Ebz88gCiqFJ/RRad3oZzZfkQkEDrVz2Q6P1/ZsXeXQ67lIZ3/wzAe
Cl5tyIVWfTCvgAA7hRXlOpvLXyiBYGTcHO/PQNO4a4XvIneep4YJ3Ie1+zcuiwmeD2AP1GGgw5xJ
0mrWksxPintUXx58LPrYku06oBNUq+HZaUKB5VbQ5PfOuUUYRJRHlqN1/rl1glr8O0NntkABGRo4
rLR4DwtxYWdI6ZhPEKOoWcSEhIhGJKJBvHGdmS/KQA1SRLXuIcy6wrEKImaBRSgjq1MaUIwZxVds
A8TNz9YYrKPIy7QuYCq4O0eMJipMc7CHcEojdjR+jYpVIvcFgQQPpY1Wj/eJfR+MojdDgkIioEkA
2BHCMokJnGPzZ1ZxUIWmwHeDRr1c8mM5HtExxqR0PHbidRlFVwfQmZk8JguvbsVRWQzq4msIkxsW
wQrlEHSkahQj411FeunFIzsRw0I1tYpoRAbyZvA7x5OIfoUrJz1ANabfUutV6K6XDGs2cEukVMJw
8NSeBnari+iUFVDSKyO0cDNQWzeO+844fSbh8Gz0GLZpPcz7HZRfjXqkr7vKgLqvj2tqLCCmMX+R
wyaUBgeWBV+wRJCNWqrDUxqBCbH7gmRcbQjGryxE+zkhsWV/Jmrv4K8S5yOF0d01w1t0wmgWuC19
RDNsPXdzV0LtvKGC8NHdRCTwTEU0hMXPihBXqOk07U5o0n9QFITS99aJmvX8Vw8TJbL/20TrzRhz
ZvLGgRh46DqewWQNkhZ6HxzX7X4DWVeBPh1LHkGD/z7+KpeHGUgfeZJz7WLdJEnGkCUaHb0dUAK1
Qln8UXKJMgXRLbf59S2nYof4TyjyukpPnOc7nKF4j5aYVYbO3O48K5ftAv8B6EsPaVrZZxAELLFk
2uxvc/vgSbanXug/rinrMIfqYxvw49yHvJ6cIR0A05oA6r8GizUA0uijC9ZWT1Gnh9D2ThSxLgOz
3K7Lom/GJCcetNV/ndKxqJ8B6pXYmdy8AaG8DXU3pg1DlNkT4m8VjA+LUxnKlqOvM3dj+G4QoDgh
y8qWeU4/lnN3ukRKBxL2QdcfcPgkkPUpB/JRg1rUTU2alELI8JKcFk2YjfnMyPAu4cAauXoOTHpG
Y5QGaFMP93p9fx9Ao5Udl0EG+KyFqkAmbM/cxuxCUlWaOrAlWsNk8Bf99GHClmBztruLR8BErmEU
BxVpVXdyWeda6HtI2ZoVGa2JM7b3RrBAguX9XoxgsKtcR1ENDTxbDv1MsHeEKLolv76KAEyx2BGO
BNjmrW2BKcw/ch/gqV9j/NV92HgmLIZPn53kHXcAjTvcfBr/hYrxkg4c5yklOOhD846GROk9r8DZ
qNeH6le2hG6vGUrznS/ehJ9F8BxiyYK2hPO0C9cCi4qgJISo7LYc3WNVYABL2mmkYaL0kqBDcGh9
6gy0hxN4ywFUdkCpHjm6C7c9eXoDlXP2x4SpxRcaCOB9Z+ENfKW6nkKQX2/ui3fs6d0sdT+j6gcJ
LWDz9ZouFdBENd1bZQhjPOB1IcFSJjdjuHjkAor0+dmIxJV6qq8d5rTK4xJlK1AgiqpM3oS7WGRs
oMZTeo5ksvSJr0TzUbJtS7X+psYi/fZ14d+6ONP2jy6BJ03v2hFcM5xEz/c/J2fZ6Q7PvKFqcSTa
SKJjGq7weDFp2FP9kam2CQiXAXbnxumJ+CRmDnQ1feleDX4SJk9fmpQVICOh4qL87oBhHIucifIY
Nbjn8/xcsn1GkUgFqPxSlzuLViGyXHD/NM5ICrshFr9NZQPpWhsU2nbXU2kwj2o3I3mJQ183322r
lwLKkbrKVHxDhAi5dvdbpzcywUz20m7lOc9ObYo8oKUDjUNTR8SfJozHIgBBChs3k6h5YKlQTR4S
CDXye3otSRuoeeFVqw04goEZ/AOZobolJ7D2WuRtfLoPjLk4Szyu3SNu90g7w10FW08mCVVBZrpX
a+gC9szQYhZmiZz9xfLpn0SB6n1p2Pv4vkq5bKGRC4YCwyI1RZuNw+QX9uLARg56AEtaJhh090Da
VhjeLhAdE+0ifUTxYgTBzDiHOUJtvO+ydVyCBGfQozkshmj+bxD/GvQxPZAgh19o93iOb5pClwYX
OM7VB6GBKsh/qUC0uIxtrqbkpwSCn5IsEERgaAMP9ALPNzHHkZHib7KkVO0fv2J2OWDWs4qu96Np
JhoMCqriEPcQK+6pTIzJIT4508lkXChNu8tzwMqS1ge+FyMPGLfkTdrs0O2LUic3N9ISplV+0EQU
+SXhOJ6h6Zvw6rvY3CR6c8305bPKaYjfAHfQhyhy9KMwN4BHcN/ahMI+/1DIkxGbo+7eJ5Qb16eh
Nm+U64+67/Z9sxpYVRx4aTzfNoHDx1p3d+5BOHei0i7hFRaRM5kJodVXVYIlk/0G0YlwO0geVWUl
c0fvSwsXXtCsEvPQYvKdlMVglELiKmPwcTCMF151jZrTlOFIl7RUkUM3J8NGOxTv94PAQgQSLRF5
zM/k0U9OtFVA/gQJRDldah/qJ3IXd6IVGRUEFcC82uGm2B+/tshMjGz8T3FUPmRh0+nR7UEE807P
gcrQkct3siGPSF8k8j8Lx27JVmdwUiKXLyoha271XPzyvbbVS31uFAjcU/01POGdgkzvU8KHVnId
OqhXziYlPj3rJGB8nutUcvrKMa0LZaclMdiqv3usgc65h7WHtsqOX2ugbpuh8+5hCwladlIqZd8S
qscNak61vYlcKwdwHRhzkk+ZGjpBr8T1vhQnfjYTOsTplMDmxdKj0LDs0i4Ox1cG7ci6BPcvhjLn
pTEL3O3XExxhNV4jYK/pKMukeoRaXZbIgYuyJ18CKoat5tq/zBHxAlvWDoxQ7BDXfxPqkogEHOe9
7I3gnSYdWucC6TcubolVqSGCsrHZePVx9dFONiKkbw1iqVbSMAe/hG2D8puq7nJLF90EgiEkSOeA
eqGoZdauVUQWPztWjeFTCpt971IhgXR7jBXk8ykwFGshwc2XotZJPAG35aXU3E/4uaO4ZOS6IUuW
uDNnmnzx8BcwUaqXTcblmoQMeEd8JywgOi8cJdZt45gdAZoOSRmGttepox6hB0h7960jWMowrj2B
GtZihsOTamvZnIY5+n8jSSDYEovUeKFTvYSksE4LTprS9wOCqX68FNxqxLsG2aAfFBsZc6yNul+j
NKr6gFexrCp3EAAFUw6CJzQ1MhfoBJxeN5l87fAKZ4AhrrP2G0oienBbmNMf5MBJ7cUB0D/0NwL1
Xc+exW5d0DiH8JefDxNlXGruo+reForjYSnJ3KxqzcwjDLTKWLMkZGuiFQXwJrpEO002VJXjg0BD
O/C9T1rJ6f3JBYuss+PQAUG5qEb1uhL4X0J81NfNhPPPpkX5U3Y3jHm6ip9PYbejqmzQN2SpnxAl
sniaDR0POa7KzXodbBr9ypMartyJI3JWvACsdZbMHzWpdXWkxFRmY4xjtNPYWWF5XeOV7DcOhoJs
Yd6A7xJX+T2uG8EBacZgZXMOyIRgW2zlNNMgktW5McjvNCA65cA5YF69IHwUC+N9KkNir7/DCOTx
XupNB+ffVvtykctnxQ+esSLGDEHR30JwDcMFk7PH2juRoM+QN5xGOeAcvxRyQQIorjAJD73AAT+x
bC+Qy1CbcBbGLLxHPNMFPc669QMqm05XO7YFPSfkt8jVYAJCQL6g349F5jL5+rV9yvJiXmmS3+MT
7xHSXuifqA5YM6l1P5msK8aXS6Z8i8YcEnL4dj3mzUJ/6SADDWtoWCdxzxn2QURA8n/1BQn9YxAP
a9lmXcJYDWNCMu5j8B1ApXDPzld8IQNPc+hCvnus+LnIdzPYRXz6oDJW2fx+HijOZEXWAsJEKDqq
6BVLiHc0pmX8odQD8oIaLpSOB87Tj9DGlG9wtfXMUpo5bBigfM8Uj9ItKzSKzeOof/ALKqDX+s6k
SaHWmM37ELePd5aAaWIazYznVf+2gPAC9cVYGiYAEwGoO45t0DTFng22KUEm1DXfxiGwDE6ATzpx
S+XS1tCsPIBahB8TAzNvotzfs/zulji2spkVep/8crFJYOkkoodlchiMHUwOGQKO6eBsrAvNJneo
bMWFuAprD+zlkIllmvWLNXtrFs3sSCCst/rhsSH3MNJioBmwNJ0/CdX7CP/RGl15Cruso8eUQyhm
wpjbA9d6R1GgCTn1/JWkCh2NjGZ/3R72W3u5y59ni68WIMppHV56E1C+O3NtxO2oKf+SgfqvGTZD
DLTaUg++Kh+j8w5u8B3/bpsXf0eQ+TWbXiL2+rjc05qqJYvN2/JAeRZjcDrbwtU2ZbuEQKfrY5OR
HILUpV3mFv+ddwVZnwVDbmpuwxjhUMcIvW6CXXmpRiyaiLzcJOzgEfDnoVVoqA6pYGrweV8bjC6h
RtzfMvEpgkZLmGFInrz7JD7rL0v/C0u6wkg81gjeKcACooNtN+WtoH0v8OTE4rxlPFxZJnFe9qsY
A7njJZ4aEV9UXyAn7eojjMkk9FkbQj2yn3PdEB5bhpd43pD4VGABY6ZAVqvIgMSlgFztoZSedL6Z
/ajZ9oddLl2/DwEueYu+xyEtaloaKsf1YSIf3kqi8L/RpP6TA4OBZO5JQI+L68+XaKnh2d0Wo/yt
zU1YKjumxHrS8CHxhBfY0z2bkwE4VkMihZibMzAe2ZrQy5E/1LPY+y1b4nWfVbnBq4ILIFEE1Psq
vRigKI+iwBM7FgyqKG7kBjGH9nR9wvvj0WQKlLQM9g8s0Q/9XZPgA6MUf9cyQK88vwcf301NRWVF
h+jaH2WAbSgBUPeLk/Ym81aQnu4qg9AMd07KMOh6aPd4nEs+igpWmvvwg4Tj9hhVtQNmqY/sXuiE
QyYxjJWJCRdvme2/hrpo8lm2eXGmNUVjjL1hMfITtZ+Ztt4teX9edT0jDTHjjOm/mNjap7LdV3P4
on0ZOq0FBY5OA8hRwGQ8Z8lZGd4b1OspClllhWJFOXx72TSE505wFOYojHeY3e/RLNVqSm++pq7s
okTpyxsKJQ+kLvSxUH7y8hdhR0GPe+2Mq4LzL7g8Q3Mo3H8UMN6QRKrsVpNQEUTCuvyZfeVEDset
8urYL8avTg4twZaiRDJcnZvQHlTqYGY/lvxq4S5BBsgP45Xit9fvn4kq51al9SJPpbAQIpW3dcvW
CYH+Njld/u8MzuJRZWBk4HeJkRPx1W3i3aL4cwmMN4DTcDi1HxkxfjsLsmg8fe0xSSXS0bpdTvKz
/AqeDfoCq1bJxT23g8D4/VpB7kx5u/5UsmdbVq2NYpk1alTLYLKd5OyqsuF4fQae4ZDxxrYdOI5n
S3etiUHMoSdv5eOUwinyh6+FPeFbv59d5ZUy9LKtxCHzhdZ49dGEaMDDpiOHO2VeO5i7QspiOw1r
HtryXelii84i3Cnj86aFHNtxSwn/e4146DXn05Aa/yygF9l2gp8YzNHcSlhWFIpGc+sha4s2Zf+1
2tfeb5DOmN2VkQaq6B2S+ItKq1x7Mcpaqa/6QEnBiQXL8jz7VzGnOL7IwvfWDPBCLpi3uMk8Sxrh
X05bzQiof7VEgeoAsX9kXEMC/VRz+/WhoxZYRlwRo9QYOGnU3k3rvTvCCKjZdU/SIayC1/JlXBY8
gwE4A3GE2d2ofbeHIIKq+uywOoP09bgfFK5Kq78tGxLGV4w0P1AdoZuvPcYWvRksp9JbqSt+mVW8
emKTxBWZYCKfNEpAuwvf4gX0bozQJoTVor4i4K2qUcCoen47yP1Rddd8zPhhiJ8hQRxGaE3nArx1
AdwKkN/8dJZpSD5K2phrC39xpTNBa5qN+GFXB8J4JA79Ag4kd1HvIx8YbM1ip8+67Y+28RIr5qnz
YUlhjZJUa47OYxuSutfB8r5QD8jvldZUtN6eLYMlU1Ec30UYivx6cpCrwWbMShZv8hUUxYtYIV7Q
MBq3X629ihsu+xqMT+/Op8GMTxE2Oda5CUS3NTQV1lkDCfHC+RpAxV4z4iOdWSdUjNiGVzjdDzRX
ClCPB++PMdvgqEC/Yuc1M84gRm6nJYtUwesogYSxRoyeLIVNlLEUiFhkq/wCgON19PCmU2XKOEac
58NGsuDdbPAJNgFvvHlKC0VC4srHpQly/MdxiTrDONMU4GUSj8okwlQXIVKvhBi9Izcub2Rojfg3
f0eq6H7WU8kNARRZTfwp3SRSgZYk7J24IkjEqosW8UfbEg4ZFcp5UFYD6MzflNGQQt1Nf+6bdynA
qPU21JcPusiyVz+J87AP+KumcPLiOxxPW3WWxMIXuxN88rerYP+oO/tgM9VAtv9BgO62C8si7Km5
hgtXYRqcEwGExaenD8E5LlAx/piqdciavemMm8M+Ke8/4zq+5bTHiYso3oMG30Cf6+FW+uLx6NZc
jxCcFm2k11JShLNnB2mQEPrERVijDx1BeufFM1crY5f8i6ffXVf97FXKi7eivGpBdUBPEg3kNgAH
CuPcq0WK5Gx3ekX0lxTF/p3X7pQTNrlFrSYpUFfkYUC5QxHwXY85MSuIqeU8MTqC/lOEg4SDZiGg
Fw/AWXe5KwvO0YgYHP+9Drg+hd1xZXbU7TNg5fKZS45R9gpGCq/YrjDvp9PISrrR10e2kIEUNmwV
YHU7CzqROAnMsjXx9ww8ivcfupNTANtwjfklGxgPcc8mcMlKZSqCKLW0FkCemSdYOO4ZuOj3Uv7P
LB8z3FB8qoM3vepnO5ZHNek6MRdPs+opqKDdENV+CMr16v8p3vkxFiThp2yxyXndZIZ6TRk8rBx/
XO7h01ccS/GaY0vWHhvtUzuR9pwLHu0ynES48PMq28GebApEMbIVGxvMiqVszxqe8FgZwFRKBCUg
k9sMI8WbXX12I7muRyeDTO/HkbFINtN0pGywJB7Ph4Kt1MQyS7FuJ3Nq45leo7+SjLn9IgmQ3VrY
p+p+s+vx1ToCWTWQGud5PtOqEo4yXNhPu2KuZbzuWLF/nq18sxO6HnBLvBvtdt+7YhK5g1yzKpbP
nT+43kIcGXt5DeT2jDV7JpUGtTDKHMQ49pjyEGU2qfXl1yeEJdzHQALcO3m762OUeWaDsIXAQi6g
SLLMdmvwpH+Tu2bFFpOjpZSLznOyJsB3x095BpNY2dvszSw1TL3kNmWqUp4UzkEemm8gVakhlVkU
j7H1SSzRihdS31VG3xCOhQPLgmQIdGWUBWTh7G1RtMXbrdyuJ4sOFVDIJ8lkYTwYXQqdijVghtSF
gam/GmuIuNzxmFawPri4ACWqBgXgdwUcPazXWZ/jV/Y5MrLQbroMAztuPUAxQrG9k2LtktFPpbkY
dXTGKJaGUYaRMuWI4KwdXivh7H5lvcyruqycBR7Dsknhh2oDa1oskkDZ1G8RUyUqVIP3HWN6izRq
QhTrQ4iSSotM7r8srmTCbWIvwrfAO7Y3l3j/UrrkwEOjePqbEXWnA0T9S09BXuF3mVoJ/WrV25/i
Zf3/UWGQE05sxrZaUudd1zql5VcjI0UweDFzl/iA2MM/S0hg59l/D+lCalpEHKeCKZSxE6kY8HsK
OLTgglRrW/enqedKiBji8lSwUvlAOLtRiTYB57jR/Ub7+DmB6k8WJE36+Zj7P/9LYQsLTH3V55ve
BbU8PPkvZTRgVa9oG0TTYGisHm5ooRCMPlf6prQKHYrb7a/Vbcr+FqsbhHv4ymni8C9QEXKCHoA2
58DteKHuUR1Szk9eC9L4jQPdwc5rNg2FMf2jJ2jCvgkLB+QX8MRZZTxW/pDUSu7W4azSfj/M3uJS
gKuJgf5kCZepvwsLkxOS1skr6QlicA80Ee3SvapO2neftsAhOlSreKKO3mdoay2WAo7vEyEjmaYt
gKx+c8rj8gS8H4LTxCn9dwdwUYBSrdG/TUekDNh2tgkZAB9LXTl0SfL6Dy09mQkr5p+6k0BFRJZO
N8wGiZM0h5jBjhtGOOkW7bQHlNuWXFMbkLEVyilQtyU0FNP6qGJmrWP7keyQ4BDqTxlrSVUIrMWu
FRTdrnvZnFzvivotUa8+U4V3UQ7j9y0teyhp+NZLj2tXe4EEMRwkd5ipy9f8wV2mVunqbXp2vyPt
1VIJgDbpktdJNHYH3RY4FugWiBqx1kNqzrJlO1Jg36PmMlpfx6oiXiZ1hsnk8xuTPez8M/pBkO9z
xltC9ZU7hB1tNFYArgKuHHi4Hx2MaxkPnRQ1MQFWzZYYM6fvkZL9nqc2p/bdU60lz0EHUlZpKq57
8Vks27yv1hRklfGC8T8GjwT5hae21gT4DRSSXjIZnoZ5yod4TsWOCtRuV1PMqDJh75+rjHwnX8nV
3+/vCwKsanxwD1uK79KYhw3h13qio5Pu5uNV2s9QbvHVdujrVtsArecIVM9ILSNo01cTyqDzSLqR
RToJw7LMp7hAYLp/8NiRgoiv2wOSNcR5b5tvfHuLt+7DQOG1zPawVJZ8JURFfMOD5ytF3rZrv2un
doc5XZHILO3NPCgugG2HuDVyfWUve+q5xYHS953AH9D4v6aVlZCbZNSYnAZTwigXq28L5K+1eheY
Dpid6YbMov9kxTyM/VwUKBOGA+oCBNO+9WjmeAQua6D2rddHN9sy5g1CwVuYwK+RyUE0mm8GRw0J
C959w8zhSiOTh3mHDlEmwvX+oDUFpMTE3NTYJqgSakPiD5WKfsQd6F2IXCoxxQGkMko8fWSLUYe6
+1pGSW6StGWxsF0HLip5Ij185XQ+HjrkSxJvMTHUDb6oQOTR/CqRw6M4Al9EoOqyjdelsv9hABHl
YgksfHFFsGw8rRx63cRWVkPQ7sO/UNkbirRxVNONM2/lQQhQoRcPWzPkYTTp+wTipVZ1bvvwcTTT
nlq2bdqpJcxTml57T/bsIs/KDRUCTQik3+dM7Pu+iynLV0oinYLDiNiVgSDQhRsx+d9LC4birX5O
7r1ceVrfoCStxek64Ka54oRpw7ktGri4YuMvhOcAzRMTEqVDQsvJ0OQ7OLbiojdIhSvqgPO74EPt
cYo2/5WcbwQp866/Il7qJAJT0okzgei78lxz017E6rMWGVnRgpEGVdNC+Z0NHVvyDjzFd/eEJL6I
UJxChj630A2kYIHgvJHtHUkQLC8Rkulqm/HwmntP5miXQOw7bWlDGN3uDAlIhPnWFfBzSQj/Fv4q
uZfdaXmH5bzyKjgMp1b42oeuOeHVf5tdagFmRNIvj7hRqM87FsxZI415IbgbB6tF5OcEQ+LaeD3W
s/zGjODURAOhZwEJ6Qmfqdy06AAJHYrl4F8h26rlLDk2BZ7TCwwqpgt9dhttrciH1b6V7Wz9JZmX
ro/Bm31wrmy4C2C/Vu8cEDOkeaq8A5FaLlpQvesGYBCii6s3CC7np+wyoZ+XsXdmlBIQI+hcEHBm
8pUyT3RWDg0VuQz9YiZ4/7JaEE3raiynVdj5ViGNt7vslsLVk++Ko2wZCQv9hKeyNH+BxfDrSstk
oOA+WWbOjeoLgDDwsS9xM2PPW170cSNYjqMjLjNsjvSaNCa/24HroYPA+PGAFWFHarboHOAIg31E
iQV3WUUrZPeqcDMTjQPzcKA9pLsy24zzQxrhqkBA06Lq12omq0I7zuBFiPLfiA3F6wCeEpU2PDgf
3vGeOZI655opmBefJcttPICHcLOi8/futCq0DLcxq+Vd93ixfN71uj/wGZxawOHx9KB4B5pSKknO
hk5OqcViDYeQc571NFxhv7mGnZefoK6u9QoZK55In4pOWrGZL3Oj/8MG02o4L8qRiUWEL9AdJXef
gd+SzZmm4qlLdWoxRxrn3G7uyBYPuWWzOoZC102zDz03MDzQslVGRlwqfcK+gdNaXdvoxURyTESP
Wzishj+P+3gq9W9Vr357h96MLeXEl9N+idztliLcaCZph/6uIEqGvJNzqKBD9mvYCVzy4E/ZSreu
zBnRlufzfRwtQluuaaDXfMfpbU/B9TZU17MocHyn+SOOwHa6/Vq8ltKxyEHifxaMF+YSAkJZWKBj
fb8k40BNUQArG8kgNM7hWZBPl43QJ5QyQM+yEiViCLqpjS8BQj7NhrxN0d5MrXI//XYcT8yz8lmZ
ZLA5P8SxqUuTj7cFugXr3yP9x9V70I5891fEHa1deCANBz62QGWDXihi5H7Powt0jC7jAkXT0fIc
i+Fuh4nXcTPRW2DU0uzaxQhSGnvmhiG+ynSwvKHtT33cVpVC75Saw3+RL03ZMzXJwTmvseU+ooEJ
TiN0dP15X/yMt/0oVutGZfE+58gY7AZuVTrQgn1S8xQ6X1CdZtW/eoLy2U/sKi4MfNUmPD97orpD
7tiWBWT1lcBuUdX5/rzv0//wSoQMMPdRd12uOiNZrlZvulvtR64+vNwfDjViIovrgZoVFMBfPJfc
j01cf5Su0Mp4d28TjaM3h/KJzHXLBKjBaoKck7hE8fIVuaaxZGIKMl0jvUcE2aotM71deFbghNmU
67BTl5+H8t3cvkbQycA9sd6Hd/f6MOaNOnHKoUSiZTZFgk3yquNcOOmiTnlSt9e5DuZ+lb9CCX2Q
3S2CJ3ZzOW4+ailbul3HhggBEPc+WHCkxH0WZSjkBNod9i2qg7x/WlDOcy4BYhlAVwpVlDnY2WBV
3Eh3QMCPwggRZXW636dX+hHBnCk6O/Mr4HB0zYQ2RPlK+59oGLq0Be/TuGEJhm5Xn+tm1ak60NYc
e2d4tKqGee/3zJvgMnsHbsA7ccugOlw6SdKd6QOw4TVMb3bm/249BVH9WLo5lb3VF+ahNRlfszkr
Zs1gwP3DwbDrQNBLIn6rbBWtv2kHQDh60xGIEs2AnE8wmqo0lMj36Ssgo8FHZlZbNY08kQLxW89n
7oM03e2pvsqBpFTGYdNUcVopMTKcewK8oxnQeau7y04qwAIKHsSF9r0Usrpj4Z6RGeXT75fLtNli
6Ujmyi36fd0VceXQs31xeXOV7CnvnYSILGf9Pd3JEMBPmPLDD7iIMhbpfmhiurarax7Q4y8VSKEw
6pPa+RmO8lCDzMmTfj6BAxPbMB6WdBr94ABfQZn1Cn7EZt8ABriG9fLb/fAbF8yrEZLa0xLtS8wj
0AUikXcBf4StLtZz1cqXKwIk70fOiD8QP8XrifyG7MtFb8SXUsNGECgCmzvnXDza1fZCv8XjTkKA
aIhGgfRF0wE+43xbc2j5l4dkRFx35BHQMT4P6nYz975hJySaFLFqeOWsUI9l0knnCy2xzdFIDvUd
pgIME7Y6GIIs07/60QqXS9KpY78FaAgcTo1zL4XiYblZVHiZRmv4XVe2xuih+hBKttThDCueAm3u
UlaJuJtvMEK4mlXXsufwNIgKDRyuqXeP9R0zUm7HJvu4lBPfS7pEKlJaAU09Oz+P/mm9og0bTaat
/AmUiKU8FLwi0iy5zsuj4roQRZQDC3LvlD4Vk6AJPDBz1yRZfGvqeXZdKOENOGMBppcoFPytxF+f
MNnxDDPU0LkyLJKdRbKCATmDPeD+hPo4kh28LQxpuIgBgpBtXPpL5i5sWOS0H2oufJnDf4An7ffe
gK0mpCGxFKIrvEK75dDhdI0HsApL/zZkL2lNzH37OcQK4n048629e8l36vTQ+w6AGvsqKF4gDxeH
x5psVouS3EHVg9hmb9O/W/o4NiwCPCkkpZRiHF5Qm2/3AUhV1Irx+Z7HzT6zHbWRpdF1+JQUHzeB
l5jELj3QSq8QFXJUGqL8rzOA8EHSI4ym2YjoVRXhXytxRLxgZCwOYgZAhPlkE3z1nqaM7/3wJ7jv
mAltsmgpddJSiLVokYOu5K9IKT8LhMg400iEDlYhv9UiqHBOH+axWN1IpxUkawRNCYo5iE/o0XQS
Pxdg1Qe0Rend2H+joes06g3BqFPFQNQYD2YdksACHC72miI6G0CWCeFyt6M+RIJ0b7k8xl6okzBl
up3YxrWR6v3c4z6lHq+8Ks91eLANnaW+fbvcpe7/5WaQm57IvfPcfeUlzuHdarWDg1GgzLW/a/xV
XAR83ZrBf/x7BpaKJg3ouXFeSuB9qfhzkOPSMWFjYTt4dm8VOFqWlBzMKWfbMSX/esyZTkoz4vp5
kBRdKyZ8dkNtuk7YsO/IklC36voEw5Ez7zSDAojNezX9BNq1L0z8qv6IPwk+NFS9uX7VhcE3SnG3
grB9pFfm8Pi48476s3k4jB9guCUwPOfdewobjap9V5SaYkMOfhDEO0N2t9TgqddGY2TZH0fIbVjZ
b0FMsbDm7Vi+Apmdu+R++ABlZw9+zsU3+1U823qMMWNyBh/s+LoUCrz+ms3Far9INrrLTryj2kM4
/pe6viVhiTE/Jghg0Q7Gbi8sZMPJ4zLCeCHv5DTjDzlqBDEodV1j5TsnltEdHXTcLRo2Q0+x9vpU
Kn0BnVajV8zhBdZhmWHUHE1QZonnJlkkAJehoz/b7G2Mi0hEVqC3U3oDm4npuLDd+rmAUHWqHBC5
o1GWNdqStp5F+EP5s7tyVQ2QY2LiXBoK1ssuJmAJ9lEpL/gNVHYwT4Pq91lb2LSl6hGM4rGw/u5v
CFysZmFLJTaxApq71+hI4J62cfND6ErnM9AzszarsMj3MenRma6+Q6C+NR4sJh2B7k0aB7I6Cxu1
8GbGqSMuXe7VyKkZ+OVe6PEMU62FllzG8uslZY5GZ8e/wxzP86072SnwHZUNJ7HNrly86PPpfIYD
XflDdi+Ce1eSY35hxVCmwKhykfOw5MEGmYBMnrYIjxcsRqmteMIiJEpFSAL1GMSuLdJJjjlIy19K
QXmqz051W4BwC0e7xbQ+LyDPVI7RQyaE5IvR+9s781QU/U5VVR2HrFza0Bv2q+WOnmM2rDRd4/D+
9POGlXEIgMDdWyqXVHYsVWwBLe1ylzpZSPiAjjsrMaoDYMb1hMg/oyJT/SdIkjuHl9/z6K9ZTUYH
mHK1U2xl6Ob8PlzvUfwZjokaX+byHRBqprsLIU25SKvMP2hWx0EGaEVTP/BEPPB6Own2I4UEjDI/
oMAwkx/NIjRXKOLFlsb5K7wmLcKuHgzQbQ5I2a+ZQuscTizeJwllnz6+SWsN8Ib89JQcEiJmMRez
SuGetz9jizKfbAGh+m6BI2tN03GDgfcY5BY0vb0aEokIpskbh3O1aBGNdEDFJ9asYFCQSO516PNe
ndz3yKnhg+NWlfvvnG1wgwItJoGsvWaXMO7wjPnLSdyh/jXFQnlB2q+dK1708A8mDwx2zLNCNPoc
rUpZRpionqydqJ3ySrYAlFZ2FoVrqVPW6EVGAkmf+irl7y0eti4YoX4TNLPeFMPet/NLIPk4XDMz
q3VXCLAH/JUrJaA4uw14P+PRAVFMWFpzEAJZ/RITkFnudFaNtq6qLH8UGXz0FXdwEE2cIfxMqftc
BohPh3XvCFD8JqgIfPxMO3BXPjXHbPN2MIhHAzeJWfGim6H9N9JHdhJPFNj9YSUyzAEBKe43LlPH
yaL1NUyubCi2fFkySO9nHqlrqDGN8OjrzfRUzAycfDXNUyLOxNRi6x1O5yJTgVLorvB+EgdTyklV
xq5RdeT5NcZStybpGqhWV+gQpOdZ7GIrq24Wvl83lHQe623+U7F6MlAdKHtGSf/oRJtr7X56W496
Jze0a60FMc4dPIgx2ucf4hAnF4Dk7BYJJkPpHCaIKbZwABmpLeSDSAO0BAFqTMXrd8N5n9APgxF4
tGwiil6CsFFz54TqeqrRhHQBqMAAVKM8H7wO5yWyAmPit1PkS2/0ItKl8Tj0cert8buDsB6daXja
JX/R+Ii/tmRGO9ASUbXHxTLwog7P4mC/SWdI6CxaGIy1lOshH/1+1PCyoapIvXyC/T3G9FZw3FtM
xySW+MHYL3bqHgqH57GyNVowtHIUHWORFIbBcafZX1NhQmKxg60cyCq+qiefSWGppZ5+jekB0QlE
IN0MoaB9/rOfe6etu1rvKpybEkiTH41uo7zcdIvR/ieaXu4o/rNwbo+iqB4VVOizP5XHuo25Y1yQ
8walw6ipAgQpiW1DTUrSgbz9G5d1cL7HnGvcMkqmT4fXvK0eHduRqOpITmmeTbRDUAvdy/OSrNP8
MoAmTRby+xt8uaFzuhEPRBou47BF+OOMPoHREw2UykwOybm6MVD7kza19rF2o4j9VJlCa9Q/vXow
X5xohjtPtdwblYhYOeNROu30GwMTTfMrvZMzm9R+NtY4m6Cohc2N8NC6m0oigueARQ19kRgd9We4
SkvGsy6iFJLurVtp0Kew2b8MvsyfJo7wkSQDPSgOVbPYAia+N4c2C9u/uDA4Jdqyfl7TpRvE6MZL
Xe/s2r2r7alA4wNOqbrjOTloBk7oY25SvkCkhQfX9K8y+i5c4f2nphpTHJ2UqMXxVaee+ZnkUu58
im6o3Fo3mr+fVh0QVRi0Pjvu7lWE6oE4Wmh3LVEc640GkWEB24MnLJ+cefdQNZyQs0ZlqY8h9kfW
fCmDgKbonrMFLHYvvLqffFOqA2GlwvW4bbNg4ySp5Qo5jrC0jqFz4jpEswK5/shnsx75DnWREQpz
Utx5z/B5lOq8t+bcvmkqKpRNRhakbrpzPQAasU9J2UzPhyZAYutKHhkk/2SMimMFhqszGyPNjE4X
hmHYg5KJzCZ1e+STSCjueHFfbGLcBi/i4l8xyWHNsxOEf/c4YWkWs197B86SCRPjTUGJl/B5Pcqs
QeITBx5Wp/UvfNG7SUk6Ek9tGvgvsT0dnxSJLnb50fcK6RJ4udAsLvHu5JnevdbRfl+rVMtf3h4y
6knchV4ikvX1jK805Vrm/cu8/KU39ezHi+3N0WS5qlLxv3qBVNQGz1YCQzRFqMDyr2ifRz32UZzz
I+qKG2Z8stnpLF8HhHinyJwXYbh4FWd6Bsw+mHVmgDI/8hXWSCNyOHaDFemgQWagBFhwvrW5IMBK
OtC0HQCLbfECopW1zSqNVjv2Ad3cjQbq5WhEsRGhauXTOJXLeMLVUL3Np/5X2QsLZ2VcQ0kpxu3/
Ej25hbM71TRmi7y7rumNNmHu2jgaCbG5zBvK8cP2ThqSA2KsHy+IdIPT3QavKNrX1eOXSY1WdT/D
hUwRUxqGmo6hm5IKOfxeinACsLrMC/QllPWA+DnCZkBc84Aq4EBd8FQO3H4i6PGdked4seDAuyKS
SOqVHTRw+Be2C7P2MSVJ2nWaG/dozkQ6F18+DDDevrLEI6IEoesJ7LfPSeiY2shvDTG93RhZ+zjm
tkM7Q68NJ33ooqzdywf2uemht5PJNb4atq8pH5ncau6qylqgMNsKgay1RhSJWhiV0Zi9ANLT4VWt
z4INdbegn2+CR0zJT+CN0MY7Zx/vCshlNNxiA9ylnYg1+4Q02jwlrGU6Gdj6p1n51LD8Cwf9Fzu0
KcL2/qMaFEChH0zPCLSVd+BA0FtJeTU7rYtFQToJjslymj554k3cktaUBHdifHTAXjwOPNpYJXJi
vnUevZCc98UZ6tr/Y95fAvwrtJ41PkWhHLPqKmNxvD1psfOWZbiV8tlymyOWy7vO5kc79oSXTujA
HvdiEJldnf7bIHqSJJ5cVI3N1UvaG1s36msB+jQ7Zwuc1XpaV16cObP1HXiqynI84mLoTt2ObPN3
Zvu8I6a/a7YTfyIJABu7J37MuHTnZ9HL3p49THbBzve+NGmrPiqhkjNDhJEK4t2+ghH0/Ciut5+7
U6TpUfMINVuOLzTcwBZ6k9Mm6Cp30tqf7ZttPQiClmfL9waRj3Z6BhXJ2UA8MnGF35NwzYNHNnDn
pmWKEQb3SoMnbIuZJsy/Bw5DQpW+0BUfz82YWx1N8QG7iZQwKn0YS6z7pJgCiUckxJz/81z3ZUmZ
+xpPpmdMPAk+bsteHkeADF2t2FsgbkKhSmY9PBQuuLF7DqAi+KYkwC32RZCl6I85wK9ZxANTtEpo
7X1H1u7dvc/Ve6rGBIo//N97JNOcP1GGSG1YB9upQrlNjVEjQaJuntZJBaMOo2+f2CV5egf2qOAs
7f/sHYoagwU4YVrLOYV+LrMIpGSxBCMgg0ff3ORV9Wqg1JUlvKnf8e5D+Jlg5kdPTG4GPmDZWWd5
u1ATiWKZ9t14WDcy+Gp8lss1NQSYKPoGS3n1JXguws5uXIOeR8WAyKcuEV+egNaWzgsb7xM4i/HG
sYqqki3HVrhU+7bJ5BLEA/711+ROL1NcmTIDYdvfIacRtFIRIhwr31gF7qpxgF1byB5+5jAmRXo3
AkyybQNCSNMz3h1YI3M970W+tSxi07nA6yk7wj4XmiIirc3bxU4dtJ1sx4XPl/Za3BTcXAw7ZAXw
StX8zKaMasc3qNqeHMtQLR6U3dNfdSBxVt6EL7aXxhrl97IJhAfw3zNa/t4VUyOyPNWih5JtYbVo
MSk3IvNc8apg6a+o7GGmUSceyBp9T+b1gw1f0iNF+cgJI81zlx7WiAzSVPIiOklHwNyX/Oe9PPyv
jxqRsQRMjSM9W7kwBlwtH/1xnaXksZu1cchvqyXQYrC1G+u7VPTNq/AB8z8OTfsDjwIHqwJUvpUI
mXEt08kkLpcoOak2I6GAASWlS0/oRAI8ZaOCWQ4hTjTf6KJi1ZnVRjzWoTGlW4TTujvoPjZVxDEK
0icpKKgzlP0I92pBzMrHk33WZuUPkBTh+3Bxwqbzn9piUxJovlL2e8fW3VchKazz/1ABaCe8LN9H
US3aGI681hIsNas/a+25Ba0gPB3eEPDhelhDFBJz2OGqSfjHs3bNbBTkCiotv27jIThZVvmzwsNC
xtvQjWVnV+Gn/JLMsf/VQnllTpfVlAfVx4REdQehuB308fjZYsdtUzjw0PnpdN0Jzf3gllY+5a1j
YFmOmxhMtmxlU1lyX82kPQE21hZHSRC7Bu5n3ph/Bayj0QB0y/di77HAlLdcLOPZM84Ief3poQms
chS3U6ZuTJ7UyLsjguMZVpC6PEj7HH/UBSGfIlMOAwedSvlZtmu4lTm4zzd5Y3eRRL2Wlz9QdREv
n+O0wNKsND4Zol6E7oW5s2mR1ThAlPIa7+rcxSoU5Rt4eTKPLeDt2yR9b2uMd6+/GmQW5PN3kKqL
oJ2lw8dPhwk/T2Az1ZtzsaLjK1CJzM8kKcLQIrGKC1G+qaDHkvJpSBbohu1BWes2jwFNtYdhEgI8
yJkO6wzrhb8tFxOjRRz4Jo/ynWk3DjAXYNygBiZv5MSB/JsS+GjlYJ0brD8/upd98udtOJ9WDgxC
Cdm5yJtqi3Y/0GFwRxngiQSIFTXqPLmNqrSQvnJGljWGUUAIIFPOLOoeYd9UpDBnpYRAkcpfYjhQ
1YcVN0XqGtV/PTgTayRHX/N/HTZDUS94A5MPJOB3IHoiCoRN7bDCteNTJRXBq0melWkd/ykOzPZ8
ICndtYPNLtJCRBf66VVfwMgrbkKUnCUIlO0imFtTrUZqq9szaaBdZ31XDPF69T31eaBuXqb6TZf9
8sgdltHrJarzPNRb9BoWmc6mO2jwI+6sqpLjGM56Pu/QjgBo1G0UkerhxD0NF5vi02QPT6xXFr+f
+SdTcSAI6THd4egtCbi53WkL10oXrvY+yDHxCTU5mkQWHioXAPAS0EDY0IAeq65F+Igliqca92+t
kR3frQSCWclMkD8eBb/K/8c+dxr0VMUuIyiZJpAW/6OR3bRQu1Yn4L0E3+nQxHhrW6ntUPvB3vgT
W0jfFX7WyRxSN18AnVr2B78yVCgYcByYUKU0iPOaXTXPJ6rlWg8d61q3edzhs5dyXLCz7aQMgcQk
FleL2S+pdcU2CWmtucGPpqhkcmu1bzLotPv+uJb/9kXdn96tUZENDkQQAZKkbUQ9lVEb+Fp3gp82
j1dW9M6equ+Zw0z9pbMXIyq8RFw/Ypqc4/09zGdqJkY1nSKc2K0PtXPcah0KW1oGc4YLgY2biFbG
tMqswdVyK2vGZt284H856vGTOQbBq4O+sTpqDto1OPW1/v+UxPHIpMVdCXVtxiofr/7+3YcdPmd8
mlIfU8ux6O8rz7YKYlCEbOx68NQGalCGWqvvFI+eY4BCHn2zwMbJxb90+eI3m1yITjSG2AwoQvXX
/FW/XEN83y8wCFFmfXo0Oqxkov6uqTqWoTOyo5nNhIOGDrpFzpdia0MHTFrPzDelFLm6L0GzexYn
nBSsPYau1dX5SwGM3vuPqWz+nGD4PYrZRRXhzWUHTvFgrqjiu/hsjc6M6eEEAScWknJGNNzaudx0
z2pI962ydSDvaoPCo1GcE+vCIl+o5ReXEwlmyY/d9FOqZA29Ef3a4beX8K7I6k51Bbc/5lhzgqrB
uy4adOj6l3zlymWnXtEULgCeyz2W6qkwXmrq7hBU4CxeBTJacQ9nB6pWP2LQHSFyAhOcCIMQNhjf
XIQ6CGqm/MHZaBhbUzBIiM0+3rMnR2KTinoTyHyae65UBzyWRSOEFJVd8M7yzMaAkPn6jleXxREt
B2Q2s6wQJb98NlGuOrtZ699VbQv0Dcu24xbAxCpn1muoMWyCfKLEAdFjTQZ5Zu5CRBNiUjkXSbBF
DUkacOcIe9kjO0clMNQHo10RwCe2L14LjQCGCz6F2bZ+lPkU04HqyuhzXfJ77xIwNtsi3oorWV4T
6Tjycs4Txyd7izAi9uZZIrV6BoZmWSXg3o9shAqAbvmLTOZEDhXBJQEDetk8kkE0zV04GDbt4TwE
JU8niT17o8bmugRIMDAtgL7/q3sOkFbfiZgJba7WANciBN73PnOsfItd1B8kVijud5DChEYeqvO4
1UAWjpxV1ev5M5U8Am8y3EcLOCVrmw9elc7uo9df0fHkHnZjT2ORkK7D3cnorooMXVeqCwLoJRxL
8ZikFGDr+YqQnpBAaQEhfHigvCSfEuc30PrSkh2HYraXTOKayblK3I0GAibegRLpHBDw2y+KPx4f
9H5vKKGjalSf2wk+7Bcoc4+86I72HlgVbbMQJu6YCvjOVO85bX3v4MZ5x2rGagnPCCFJG37Aa+j8
ZMPDfkqeagP/Oj4m9+NajfXbDNuVZCsdBb1+fhtUmYX/uyzl5iAKp8Eh7cxWLQNRej/yGWoXNx29
f9CJo/fSCYnBdZaOZJ5Lzg/PB4rKuTYychaeWBMtCrFdoRc4NcvLDSR87uQPRavJUH4uy+TI8fmk
p+YOlaNzd4+xW/8lK3Df17JkicSDJtLymegk8uPFI1wjbwwyusySH7RjhbhcdgbjrCfSLZauhevx
YPqTvBkkCDJ8EYKduWODyZBdI/nXYtgtom77dSNMEhLT2nSqkyFbzhoCvcMl4d13vjVVvCX37jME
YVwdRxsUOXVqA4uw2q22K+o8OAuix6wBaYOAvWJ3r73kqBe+yJA+THwR6FI6uAZcT5k1xpS5JFMl
19mHqTRAd53wZEr2Yd06wB/pPHx/wGEwbasuGDSGTdClYR6XJeyeXjrVj7RExUWIyOIKLhOkBaDU
tGiE9gYjhABvzB0Q846r8J0MQrIoHz5HYYa3YB26K2bONH57hRxsQoCVTvdBFFKGC7nBojln9VHx
HWMwgQKB3cw5w2HNIp0U+4k/OcXIsmiXA88kJI81GSoITBUDIZSIOnfRkHiJovh/F429FIe3pDYa
z0xSnLT/9rVxh0TZveYGdR305gUHopxcutK40HWMgjUJiUfA/uT/SGhKYiuWzurW+EcdEjfcVdf/
bqYR3V/6Vd8P9XyIpSb0CFeDLsWd/8ub2Sy4Q2EZ7Q71p48I/TOIvA+ymdh0mV0flgXuN7efFXCx
U0z6GPtqxpLE6areDzPnhYDKtQFAkGNk/nU+A8Jq/dSfD66hPWbKNcTFixyQKV2bR/yH2XQroVAk
9PzA6Wr0aW9297Fypv64GMT1Aw1rhZVQJOpZZPHWMEt56vCISxxrkRYrX0MY4gSHjxH3wYnrU/2g
Kasr0EwNdt5yKNCVwEs9uaHqKltA2uPCdxB118SZcgW5AhWZX9+XJB3e4BLLdGnVyymAQqXRhzSQ
72Up/C3bkXuU1cgc/eOCTDmwhtqZfR2hIg6QysEdT4iAbVXDdZPsVo8N5iBSlpFN24OsCuNMCZ6o
c2L+UdSLp+zWxtpy+UjlfvG3MtlDn9P8or0o713kIqWmILnnnCP/UljRNV5GwR3OSsbLWGS/J6QE
8Ka7HClDnINS5r+/jATgkR/sRYSCqbhOqALjXaz6nhYoQMnfG8s8VlTYZ2e7gHSS/OG/HwUtyqCx
eZOkLwMOrZjSeIY66Sj2mo5WNN7q4Wmb+hzJ8oeegPkyGsfFGVNoOQfzYjkZkC01QqP07ibjtUCl
ACmVCiw99cd7hNIInmAYTa4nOVzFtjtaU0x7PHN8y6NsZd3zt5jf5Z4cxzdz419oDjquCaEvfylK
xWygPvJ0bEbN8AG5hI/tzCeXgzZuYDJWJxMluWC6+SN+LHEuyjD2hQlcCTPrOO4j5myA/U4RxjzH
k+Kj9ljHDKE/0EhAo2kVuEs6O9+cT+HJ4vC44p4I82Q+U0EnFVedFQuIIvPrCjfqDvF50HFnzHFR
3yI+7p4LV13hjVZqUJo70EEqX8WA0COjakDbuvNZT76Ef8HZkSn7sEGSG5Fp8PFRVMXPeVtIW/IW
Qd8lcCUr//PT7wrJW15yoJAXPW9CGHkxJNxt8J2rTHXd8JVPEOgAQR6Rn6sWem6wgat9C0sKxnRz
T2R+3kw8TNbkrIPD1WclpMZCxLR+bj8x9orUUIPRn1OGraTmReihaT+zsp9iXMB5RyOCpWpgRE7E
egsoYV+AwrPRN0pybHZEajBIFGbAkjQHC2eZfidIVjCUnU7Ui8QIO3z57920QkWdmNjq6rQbtYwg
F8uQ1BiWotsWXdZRmTkLeyeTHWLnvYhncJ6Mcd5nyf9Y8QOaWdQj9CCL/SNBxkf5nq20skhWvJVw
ljlujuvJH1BJPXmzBKei5sRpMhaM+r3dCJsXbcc0UkJDgS2BKCbGSCPdg5viru+3o9BmGDY9Q5EZ
C8TzXvuzxsK55nOWTnKu4Abb2v/k5sY2LrH8/WM8WKLwo7INQ4OBiZG51vTRGbqivjIRSN9Ye0Im
9lLgnRKa3LKD9AYskG+XvhYVYSvesZ2Qi/rJ/14iePB1A80lfL7THHMJtCZHqcCVxaqsJZXrbbdv
qJO1NlfIOJcB3Ktbm9N+1LjiUYHM0W7TTwJTwyRXfcYrcHA5t3tpMl0J0uLAJmjf6wLisZZsr4Td
5UNHj4ns7eRM+7eNKJ4x+U4OrLAh75VZCP3G6+6as55oiSnvvbJhrrqG2WoeX4UjHgQKZG/g8UEo
IntCIPPmGNfHMbLJ40lroi3WIwC+xQMzM/o/+E8HHVDdl5NBF3LLXSPccGaWRMFsx5H1kXTDej+g
G+QhzWhuPM8ydxmSU1cI4uF8f60ixnMvY/Mhbm6k1/5apbQyoXWjIjtiEEt7ccju/TsNEe/S3tHY
Tc8Pz0G5yyXlI8/1aA9HmUJr+i8uPUZfx4iRhHwhH+m+JfxnohS8Luqafos7ao01zHAUdeAUwPvx
YWei+BhAW3YcXqBBM/XQJUjdaO9WEAPehcbUSIerYKIGd8ZiKQVvc1b6okkWaNs+ZOJQb8onevWo
21K3B4rNI5+G7RdSwkaxZFaZTLbIOjdQd/tTbbxRVrSLxHcv8pj2MKKI+YBiOcKgr4rFmEf3Ahlo
cLbuzMo2P52c3kQkfJgzdHhpCoWntJkeu7os4i6uA0Urd6ksWck2RrRNkcYAb0Bz4Ka8WZ0tVwEj
EsbryGes8izdWiyqhWsc5+mWYv5pQmiXWAvruVM8wx70CIQZ7DyoS7FVCLGHQzJ3A8gIxNJ5+u5U
Y3DglhRX2HaYpllwQhxoFCk6N+VjCYQzlvdD2nTzvn5uFWGVaqqZzvh57EXNI2fiZzHJdnbL4Zj4
mAy5IxC5MqLMRrj6s2MKzCl2mXt4uFG4K8/mdXmydBvsf7sLXTY2/aL7KlPZPIyNmVqUngH/v1OZ
4qTIyaRGqGC5vphCblUMDAh4G4jHEf9hMpjyKm0NcwDBLpdXYfC3xUJJuiIZ9M/YygibbnqbJCQb
bC57RxEkVq4md5mMpqO5LgNtmrewIxb0GdFHNn3WwHS57rgnBS9agkACa+AJHrForksPXQXH7o7J
zExRa+RQUSehm3kqzZfrW8fIrtZ5INUlw8pp+co3znkkCZIM8Rn9qEojcDb2QaEBr7uM8vs67uYk
w/mFLF5lU6l8b7Q/IFdfQ0ZO6N8rJAacOoFV/oyUaLMiIOkKE5XLy56H2jd8QVXfWZCexN95aylS
+ZKGSUGPNuVRLgMmz2R5CzoKxDjE1OQwWrm7/o6D3F2hlIxGqIXrTkf1+yj3XvwxssT45MLUQvxk
zwaLsIusE2b+AetUZl1cUX7rjhcz4WeYoPSme0OTU90p3NMmpOg0TgYFnoQ2YRnec7jNfG7Cvt+M
yOyi7owHmGTjGEeu9KyzqbSmCztwutGmLEXmwbplylSpx54PuaSkusUZBcMKziUi2o8LxkAUoZW4
u53rZszfnWzEFqNF6t1WuPga38TTwgPb/87/Hw81jW0/pOvKqgXTFQf8RYCYKndNyNFPE27fcpd5
xXz2VPR0n3Mo2pI6+mYin8oGuQUiniMiwGIjLGpaAR4pxIekulc3Axq+k50F45HCoV4j99b+T1qj
EjJ8Z93iBg4NeM5JfA14ElBdeDA3UzjCa3Moa5LRXJTcGepSPN+4myOqWjjROpfAygUqwWSZtm0Y
xYNhIdGd/uzj/ICorM7rclJ4joOiCicYpPLHHg/M8/xcJkT86Oo+b82zHLxGZpKcb876C0ggpVTT
4fa+sF0ZDWs/915oDkyBoi1DW1uzo16iYrMNfeuc9IQcvRPWfKb7abqkpvRk1BXG8yb8qmKLVZJL
Gi7F9mAQN11XNyu0/VpZ32g4j29HnTiNl6bgefwJYOR0Q62TeTeolUDeolUVjSwW2Ak60/HMWvcQ
YQNXy3BrFHkXnAt5GqVB89zh8Wo3eV78zoRBuan6YiW38vkZgqmdqQRUx5g8nToYdF3AGL2QlnaT
7bvz1N0esfZSjkO4+g0sSyu0mynE7RVGTlx2Py8ZxIVVNvUA2ZkD6ZHWP3AQKncJm4uV2gh92KlG
gRUAZ/ejKeJgRWlQeZqXrZQunWlxW3SoUstYQNtgEi4n1o8PqbD6B+UniF6jnMTxBDJaAixAjK30
sPX2bDwHXgRnKQ2I1Y1fwoWp9/SIohYlgTjP8p/iabd9bS2V0Dfe0CYtIdDitR2Zbr/GlK5FMRmX
WcOLh4Txrt9Z7CZems4QWp/e5hu3EU1aJ2LbdvSYb9ycWSy/8ZYhLBTlP/u/Wmed1JtdcjzThIls
RJyxsGVLWTxRMaBUcGGw02Rceqv2cYghQy0LgULyaJmj+AK9OiHFwKX0gEBViNRsoPDasdLszujQ
7q25XGijJkz2/rDstQPbhzuSsHj3WvtTP8MePNhEqelZQVA6UoTi5dGnvO3s3USNaKV0Co8FGjlA
4Zx0gVxAcyd5DiV14+L2WmKRFz1jjkTR/NmrxU9BRHwMfuzbUwPMEbcXOPnK4RVWAcjO7V1/RU6g
xTWWQDoOGDqszpclWDGaeExcw1ptMIi+7wV1F8aFhqHfeGJOw4ULKI6b4a0SNAPJ/KbP5LX10dUA
AtZiNLw0b8Sskdk5yM6eSGwRqr85dPr1Qt8s91OWH7WQSVkVcfTVLo+A0TqIUmTLErBVb9ouGXpz
Dbk+BYWh8a8bhiWF8QqvxR49UaqeOp9rpIylCS8XGZ02yQutMPAwzItGyBEGWJumPZ92/DMhbquU
3NR/8ACiuGApIXaf8chf10SxySyE+VNx4kk1BL/DKw50tAmBcpng4jgnkjxKK8y/qkdX6cBNQ4U4
iykNUv/oGIDumXK0LG6NwrC4X55xil94ZJBvrZrd/MkOfDPD4J+pogqxxbBixhJ8khpetHJJ56XE
IHRABOzPFbzUSNe4VLG5nE83EajrGCl3x4qNdPKjcDg773VM6EeGkLWyFCi1EpDv4H6LqGn+k/F7
k+MteIAny2acUrTPHhlxId3VPD5ni6xzIuUFvTHj3RogR+8CHoj1WKKAgMuxw/zifY6ljEQ3LoY/
6T60J5BevmleChYtFcZw5urkk765s/CooEnFVeHwd2g1KZfYuezYQWzTnynX7+rFY24IE6D2ii3L
nfmQpv//2Mg8fuBfSs11i3XdDYzGeEE/w0b70JYnOcjlKBf9a4Fzf7dnkM2QSgRpTrf3NpqhExvJ
+4VN3N+dYBBMg4QLZq/aa2I6gKQtK3Z990M8Oeti6eF4VVl8PibHs4hvnBdxktMd4dGFwTxMNl/C
wybY8u1/QSB00YIsYMhvjRZ6MO6KcMXFqa+W+9TQlhTyIpgT95qIfvmEgqyygfed8WvrbTt2kjxI
cgnfZVYj7YQYVknweyZanNT/WZM6hDm446CnkeYsRh+tiszfyUXv3uF31J27g6TBkfmCT9UgzFop
SfPPMqU+9zraBbv4U2YriEcqWaDS71lb2OVKOI9ATiCGPFphydp+SxbP+nDT9tiUXf26NNAYG43U
msC9Bt/2hfYfTLgMc0Y5F/7t/361ldex8LvkT3C9r1vkHqAfusR/zVrBnReCw1BdTI/2lBhUkZVl
lyCZFKq+MH5B89G5zElaA9KJ/DTM3lnLTG5LMt3JkZJTHRQIMKemP104SbOSpHuHrIFtLkliHMHl
HWvlk+bcNuO7aW9JiqGVR4zctoGdE9gcd1Tld40WwxSMEbuZqW32sDkrj76vsAk+iB8L3I0+b1ZP
9MtgihNDp0nzPAK1AQ0/PmVyFF3UJX3f7s96C+GmbH8SmtB5hnVFfT8EpqyIiwEzw0JL2km5VtbY
8o8bMMRo3/G4Xkz5g9FOcnMqY84mz2zUV9jB8BWXPqSHhxmpOLwHJDxpLkwieZgrnw9AJO/gyOhh
DetjrwZxCbzVwBB2vcaz2a7riK+dZ89ndbLLbsQT3ViZ7UF2y33m/PVecrWYufNZLIpt7Jxs2CLs
qY+fYz6WAAVtAri66sBSewZaYxhP6dYfXs6FPaSSp39BqLSLZiQ+mXBsygqRIPXO1Bj7uSY7f0Bz
h3SoNUGEvgDdiDeN+8xU9Q5aZCw4MM74yqxgwZ8XS5h2tQI/QSI8QzyizcXKyTd2Gw+adGHSl/Hz
ZGAPdKdkAejyhHIc+dS5kGNfijl6+JvE+WYGum5miMh9lR3AgaVvlqQ5BjMqRF+wrFycv83o3dL1
bLtzRIbR2JD2CX54E4D7oi8s/gl8K6bRkbuclV3eaUXpo2OLm4/lojsLH7Kr9P+hQh70IpD49njZ
8TOGnarKJNakm6iBrxXIDLMZx4d3vM9wrOHO32oJpVcb+nA75VDRn+iq0d/MhLbHdoP1RMTZjPVV
4oWZFZizD/yG+II663JlpnYF0lTsNOoBGy20jj8OZtw8/15DCTDx/6hyb+IGCyPOryoJvVSDuVY+
1jxwgg8NW8csANEQOJAXJY/g0KKKarF9gS+Kb3696FC7FgPADCpu8B56Am2av1112+ilLhv2JPrB
ARQ85ZIa7hL14TzZQFDwde0dxHdVf19/6BkWwt4g7DaLK/XUH+TxqLrvWGt48mSOw/yJ3DWE9wlg
757VrM4L+BuTw96hgtOvwMxRv8kWyiEUjUy1PEk+iA7VJ/MevZD5bkujGp4T6O/xkPzoTzNQv3Is
a5AL/iy4W2udMDsWr/xpvdHyGPyegqS1jMKtY/UI41mr9Mpr2jyi00tX1gM0V56ctweNqsaHy+Iu
qGg4pW5IDfM6ykvql8dcVhugfxgbjFcrIPSzKGNlaBMw8TrF2sCLY23XVJQHSOQ19l2RkTK74Zy/
TIO3j0EmUjmGdgEbylzzDU2G3HB3LfymRihhbCYk07pk+dOnoLTVR0wcGjvpzzv1mD8f8AvckbP0
aXQKBUjsNZxiS/vCzT6dlrBPteX+OGcLZAonTKiXt+KdD5WAaEiNVDpQ7q04QKJYiEfk9QdWJp0R
kdbuilYLKf5fBUNxkrw0uBZ13/qxKQXbec8399w/rLTYgtgFcqMN6vFEjsbGbJe2xkPrL4Bi0AHU
Jg4wHUsofQGbo2ccluUchxK1vdS+i4mB8Cb/LZL/1qs0H03K6Nu9WVMpDXt0rOysH6Zbrfd2Sdvx
ZiqK3O8jJ5s54LrRB1BPFIB1d7YlzoU1yoO8HHrS7NMtX5UB4KFuPuiXKytO3QA8EHgz73fXZJv/
1NojWWeDp8QBjKpFtMb1qUk+3GpHE1HwbzC0pQcT6xrMax8gNSvz5Ry4Rdqcfyeq+5dffZaXAUWu
HyX3qGOXJ0grVW1KtT0DAnxNJDz8ch+Y9mCmnUIx9vxOjUVwRKo2eT3yAAv+sOeQw1MBta4H5mT7
9wNeAl5mxkKg1iAf8PdqlCE2Urq2s57WskzXXesM4nxB6ft0pRcptRRqtM5EplQcx6gnGCS9DwLg
ubkuAnSK/bhjutNySdBsvQZnNTEjTzaYcDNpBn07D/VZ4qtt3O/a50fLcmFQ+MeMkF+MomIu3B42
TUkyuExTInOZoskhtgfJ07rwjuuBP2KoQyFJN5RDahL57iCy1VT8f15gRA2I2ZCW3u4BY/cpg770
L6G2vqnAhkQLZlJK10bcTTYFFn+t/j3yKjLS2t+jdZm6ZnfpKF1MRLo+72FSOuau8X5WWvat19rV
MfeBqEmXumJxqT71//AmbIW6iU6unkdcHrO6u7+mDV9eN5qRtikOgeo8+ACKmRz+OlSs+kW/ksPR
gIUhX4s+JRyNu363pn1UdxWEbB5kbaWQKIlPgoojXS6K+SMjqVXDuNEe/0YUBViMUKnxf/ln9B8U
2MUR0iacT4MLsIBLSUdSxulJSgp6IC53ete7hZdxL10Yj772HS8u+dUmeNLbYJ5/UphIbH6/n7AJ
cznQeJYpwiTm3+PCi9bGMdpit0Vr8yqLJIm4D+Al/yYWC+zQvGzhCbMnnEI+A60krqYsKltFBfru
VEGu43Uhwb1jA0WmjrXi8qw6ho4bnFuuKrZwcMX6fNeGjHzWPZow8gz/sZ0LGVS9ydQkGnpCj6He
xYmACQHCJca60O5pwAyTyiddSNiZweQANmd9huJhDN5N8XnwLVzrpJo2z6G4WxFqTpQRR4ixcKto
Wyz419s8rBBfgbicoNsHK/Db1JsRkln8EaJ/k+ls9wzEpGXooW2DSYpDX9skU67lYatQwoJdAQu2
5KC1VxFQ2WzXSXKCEfDSLXaJWmvFTcWXfxgN5FNk+D9kqqUD/HfWCVRqctkXuAbZ08VrSaLyPTHY
mRbnxrQEG+QlxpW+n71j6YF07ZElQinnl12unKz4oPQOFFqI3fXGhi5gSoCOULqSQuG2LnnSYVwS
1rdo6NdIheutbHVvmrxspM7gnyPnNokY9OO9UJmMA3GIPypftwHnbToL5e3mFFxvXGwKV9p4Pgt3
7EwrqJ1UXx6JlMJdIQjWzpboS4Jzm4rYF69KS07gO4VocV46vvZjYSpCThb3LI5LmlosOmq6j5Hd
cX++qLz121Eqbt+IUInzgJvJj+OLlpegyHAgC9SoxBkRLD/3vOQnVVsUdbTr1aQsuWJHykPzRfKw
exoYvaYrPZ8PfHLdNOVeR218pTFmV/kohKjZd609Chxp3U7MBLgrTEXmMkSA26on6vFnvWuQlQkv
hrwgd6NE9HrUbMXbMJbD7bstxxHjTR10KsoK0YO8Gzh1uGrsNR80SG2FHYZFDdevZH+FpL4Lk4aK
h/qMmR2b5R3ps3k/g+nRG1uQW/kCcvfY+oW58byrqcy98TtdfOhapuQftxy67cPUogpeG49L49Ya
JAgLn+OCVZHTBMMyAKmtEJonQhDQ9wTPhIxJ1M1JBy1XDr0RclAmdSfjNuGWfqVjfihvsxedOVOv
DO1UmwZdEsQMWml1NmUh+8My3ybgZxMQKEtPnUANTGc0VW4HXSpvoptsng5IULEnJRnkuQcWHeoI
hFOEvuzcrsCcW0Y7V19qtGeb1U1jVN3RV9PpA9oWBTr4Ne60FovBxBE+cmZtmzsra+/29MCjcNvd
x6JdveVOuZnY+3mrMQHRPRBIZnA+g12gnw5Taz9F3HZPfmt6FfTzbOQNPdTaDiRurKDcnTMLXk2e
T8UyQJMzJ3KaxlGov2AcXlDSu2p6xaaseROqxyArWm1Usy1ALqW+dRHkZgdtMyEq0V+qG+LhdJHD
t3DaNE+fOwZ+VAUIq4gxVV3R+ZLzpY7fZE3E+nNSLnnqGqU/zD+B1jENTq1MOLgRJoSH99T428SE
JOnlN7qfqkvInri0jDrFy2bYDz+u2l08CLrVQVy/N6a7gS3Q0L9lkx5eU/vM96Ml+h+KnM74QcyD
rNYShE0FpcUBlz7r19v43cleyw+3eEApmnNVZzJuAXow1+L39FjK/xrRVJz+MYfnFRydbG5ckvbH
rbeJWJV8cMyMr/yjhsa3zZghTtDZ/jenpRGKTh5ncu22WxWq2TyErg/cm7q3PFutn3hxv5Mv+Oyg
c5m23jy+rZSgKn1XtqLe0Sduofgb7FbnoY1GZKKZMntYKybu+dEKuRC6pgBg8prulu81t/kXhp3+
JLxBVYlcbdwVNHUsad2IJB9/CRHAI1y0KsZ+NNCFKWfotKPadzNBNAC6KxXLrN0Akkl0hK9OSV5G
0Xmjwx0fTFxx2wU8U3SErykCgHH+lddBZ5wkoaDNyGUycRb4r+OM/WSQ3WnooBRAWR0BnNnAMO66
6QNKGtahS1g9f79C+SL6mT2t+6BhEqgdyiq0mtVncbJ+R4c7ZfVhXhGYxpSbBjhsTMWgs1H18Km5
3jh2A6NitTgf+CKWX5+aDI/rkVngF5wQ21aC09vJk5aL2punJpsi8O5NPcXkQfW9XByee+eUjRtp
kgug5EOuNg29QnhdmcRwIN2TeS4B3yChWQqF2q2PLkNvVlTTXIqorm6VZCoWbKYdqm3z85SFCcYY
aOw7J5D+5NdoTiDnn/0/Osb1RZaja1Ye0tpz7p+pL1mFrGdAT5pj9UUVfI2mdIi7oXCPgu8xVoii
KYTU9aSYnXb7iI5r9EgnLoJ4JtlmthOeWITNCpoE2PGEiadeL3N6Y6jXmlx9l6B0WLvJaoXAucuk
sjIZH9we241TzAIpHKTtEEGm6JPRfft6cV/7bJo17X9uReRnFZ055vvgdqmfDci2n1oRih8ShrfT
/f41iVBSLNij37Tlm4gTpT2EGEuAFqUyq4M8zx0PHy5lmDyU9UMNmzmK9R27EcuNywywCuYL+k/q
vvg1WdAPegD6LNCY/wtpweKRKa7Ll6y+xPLoD65KCVfBplDfNrYsrIBDyndFJMXZQ1YptxeNGUHu
1ce3C+qm+5PZ+PIbl8jsi7ABLUVLEUj8KYZOAHMn4YYYfGeu7purXiKWpPcSPnJX4izxvrayCctV
6j5UD7STJtWq/J6fOsVTnbaZULQbYRXMxNnDG9IRw0afDyNmSK6s4XA5SORgrcwdeFZQwzDdONvn
0Suiuvayr5RcybhnWAE6jlnS9H09s9FyraB1H0UEipjucH+2zWmI4zEAude7bBCciY5nDKmOQvpg
e7RAtjDvFhZm7C8+IpoPWfwzUIUHsw2QgWqrhF+Vc92jHmAVRnwB6PJejfgmLe+gNiNEFs+z0MDt
ddDABULEP3l/XqASEGtnDDA9OBW02Dg9UG89UXEle8d1CglfiP6EcSF2e/7gIFgS6n4kyxO2PCcD
EVuTMoslJD4ELYveUwBVt+tJRCEzExQOaSczvQ2H+fjeqtNG6ROIsmk0cZAa1dhs+1qxWGAW5t5F
RQyRffIwBvSAt95TqbT+B9qEJR24N+hqDeahxOsE/AHCn08EjjO1qJJUS6WQs63iZ/htdJNjcGU1
Kn4d4g+02ILQdIPtYXL0N/OXL/R94cuDf6kPTw/KZuK+Xakd8kUyaq9KuPA66QSn5A6Ru3efJIpr
jnxvE2O9MJwpFkNtvyEfmTdhrqpJZNQBOBfE/0c3RLjtA9TaWZZvAn7c9pKjuOAR+8nPJ8pZhegv
8evt0fQjp7k0Ee6O1hv8yUlinJflcwWFtVkw6NvOJXVbADde/XJ+3ARiVtxCp74+R4U5mgEgq+Li
iurWDAoMYVu9vlrVzQ8YoPGXvwR9K9v5/bmAVcotBC1QmEUNkoDGp5xlVCAEWPi7Skf1LinCyQ80
WWFQRREUi8t1N5Rkq6gdL3UHmedejtwsuPHw/4/Me9FoOJRWsxihxbgjKdQMWuUMuxC4gycWRDVC
SrE3qXkM1akt9qarKEEeVFHY4G/VksQYgLsLFsb0TeudJvRqRRGvf/JLfgQkLIoT89Jx5ycwmgpZ
5IEoMHo5SKRfW4IkyDSg7YqDGW/Q9RvXfJuQkU1E4OJKXh7/Gf1z9EMI8n8Dr5xnXmdfK4DPY2rb
RrWuMAVHSw6ek7uK3Kt1wfiODHqjzqk1T8HFz01rpm6xImowf9dp/X71YrAoUD2Ep69R0rW/JgQc
pFaqAD26velrM8pAGWGLWNS5ot8Y8T0LEDC4gWh5KNsw33xY0Icz6Fm1WckdJa9yc4JznYm9yI8t
pjQeDYmbmU+cklUD8nOfCl0Wj1pCD0hK4Z9imiK0TDtKG1oLTQOXRd4q+N4Uip1nuMqi4OGbSfi1
rwa+crI6g+cBABh6DbPIAw+1qJuN4dnr8yU6vu1zsVbbIaaVMHZ3SRBjS/sshCu6lW4r1AZw2i4M
HIaC5ohFnftvPy3HBZ1ID4JsxAp/KgWpVYW7ZCETNTHp+CI6o7b6ouWLa5mALo4sl8ELtQG5+XPs
kN8L8/oPwLTGtCXKO4GwQFrVoaVvlUM5xTJ95kN19ccWBvZEDcFz8q4WokErBXdq2cdj/X6INTl5
qODZLCB8fcm12C2wT2A83VhLqDohaSaUmpcNzfdlbj97kEOdfnptOzGsMEaa3aoVXurXC0FVoD4v
7bAF1Go5CBhzEvC8lbVGUnDT5s/1Us4nS2Ji6qAyeeO3aB4pjyC/2GMalX5TtTaczhqNJp30+TS3
lRywGimaBmqGr2fo382F3kH0JuUOu/78M/QJBfU8AfXcY5Elv3vpdu5JkQQz7jOlchiNKT13H39p
eFbotVvWSOnOvgDAeVrKGHi95K65iNokLP0fqudVipPhD1UG2aKhv3HWs/ppIyDiMRWNcHN4OghU
9HXM1ttDlUjfJVusng8nFISsGH/TH21BpviMhRZoNDYxOBWKm6r+LSE4nDXJQyFQD0yGoiuKjWmp
oK8hR4tU12xs2nvC3dcDkSKMiIB8O1RpaJBWdih33rSXMtlkzEuLk8lq1hHuTi1u4Ys8hLOyQWA+
Zhc8YUDshBGOWgnPMH7kgt2k0k/Iz3d6UbUBqQxaQl/OqhLPZyB5xNdfNi+zZvBBO9MirwavD5+l
CrhOM8Y83mjKjJ4e0a7k/XZWRpXPN/TsBTacZS7Am5g0Lqr2C0JuTaswaEFAjoy1HTvV4kSEvt8K
AxI1SjC71qHTQsWfsqZxmq6YnR045VZFJelYQ1cppE5H1fjirugWuI+2p6oygdhI9zpFOjsG2AZG
wJkVjI0mh/oHGNFOBJjx738jScsgith6c61J7/ifhiVFJ5rCiu0PPr7kyacTolOlNsfCnnVkQVWg
VBOmDRtenDIz91zLh2FKfE2d4Epggn5IloUwQUhp9CSd/x3+H0Xj+24gk9iwwzreklAyRTLR2lei
PvNzSNohgEUoOj03L7TbofC2W6o/V2ApmelNWmi+zHdU0PtIOUIlmk6wLQpUp2fG3LeUAFQ8Cjnw
B1fHOgKSnoeOR2f2N5HfGQTqNsyLxssvUPZDjxPQG0QEVx8Xf/BeVUkC2zyZetX4QwjV7igcII+l
7Wb+SmbGeU6lpOO7qtDmNdj1l1xURjYrflxG7B7L5RuAo0b7cBcrw8srO5zWprcYZFePd7ZIM7vT
J21sNRpH9MMeMYhva7XDJNYprDdAXOfS2mMCs59lDmcJJ0P9J4tI170HYrJkcSafcXQElYzHjGPY
jDiL0QodnDa3WmEyCTY2VHFttG4JG+EloDMwQRspkuRwRP80v8oygmDze+b+WdMmHsmrXiWl816P
5m7WQhqEH3Ye18hnKxn6x7uOXh2LfN70ILmeOMR1R+HCr6QCvAO5F0jbSpL5dKnmoxdE4OAALOlh
ROaPWnUJ+ruTJQEEiIVJhiajuh42KpUPAjhA0uOi0n2rd2LTFmJZxGtvJeMHq+3r6uoM83wJPvN8
lYgY7QQNyo6ve4UZULSP6aiHW0YGHMX/rZSVE5cuFTOhF9aRk7O8evNVTkBUINAHrmzD311bW9+v
2qJhhZT9dOcNewfxS6Nl2xGyioafLgtNKXQ2JcmGXHVjQ9JdPiCLNwXTwVKflkpIsVGFfk/s5CRq
GfKCaZZdXohqjIbcITyyFdSTwnrPCyaf8zaTh8/gPkp80ugJKJJiRB4aa1Qrx9yKtrWqE8U22Bc4
zkDNXiD1QOmm/XKPLLsflvORnH4V3bsJFVlN9EfirpMMVx/edRPxzyeMJXPeahWijibsDTczNeoK
ZeZtaJN1EKUsT6+fwOKmU4q9XYKriUkZzO1tm0ovwidpsusSGbK6S8UjZcZdRqZmNk0m+IR0Yoj3
K7JYxxiTmuLpR5XJvsCUgPcC5JtgFZc6EqNpmwfRcam+brKbBKJ3qCQ8NBKHLL8S0i1zhiEJ8BWi
51t8lRoAKWylb9/f+tQRp7LyID66zUnxPC69YHM+gFMYSzYCxwyDsx+3g6ApB+07S0tozlZn2T4O
VQG6pBKxrRRKfwfkU8v3+PjeCQuVyBJWVE4ZrET6vRDluvWxbWt52qAMtm5TdMsnvYaVAnjIjNPl
MXC61YDFviObyXIad+oi5F3mUONqHddJu3Yb3VTw1rYNs/x4TqotIyA/AHgy1gh2jTPHFWvnY402
Di/g/FwPAzsE/pdLQVG384834H74wXBV3PQSSAaXoHJ9IjRW1UV2hC55EwnpM/munV0ZMBrEB18m
GqnwCMp8ADSE2Sdf0K3wi4Z3zMGrZ4pJ4EcbThFu//bZKVpL0C598GYqCGoJohvbdr+er+H0LGWY
ptAs61y6e7dhSCxsGZm22knBjkDrbGd2v62FIWvB71l48ug/Mk5JtySZkrQg+jcRph0qVHKTTFCF
dwtW1IW5+pVymknqJXIqTJIsR2gyl4ofWhdFS472tf8M57ETLGWGEy3Ljvt2HIUENHZORcUSJtp7
Kj2Y+cB5/jyznfGlhLsDfRYB8VCvZZnJiKk5gX+KsN2D7p3UcP3uvjvxx3i16fyNaJtAGRhQKqbO
H/gmvLfX1Fi9zzacrR0nZcRcV6EEfx+ORkOiIlfnwwAZXeBtrZ3PB3ljZ0+sjhX+JcwFxjodb5hZ
lvxvHRWDBBvvnC2Ai2IxswtVIjTtln3jvILP44c91WuOj2bSRNCENpfhYIwkVR/KZxLvBP8G+IZE
8yQwD1t+lfEaGElRN14kSY/K48CAC1pfLFZkslUvVmPa1bdNflWnydPAewi6szx+U1O5fEg5CVDZ
ABhp51BzGb+htLUIrHLeqFWTfzR7rXr0T+0z6HA2xegykZYwKdvsi2VKv8Z4hXuYVNzu5iFE5lI0
l8be3CS1ArFdYbjZrRonqWJsQQ/hGlDjcW0O5ul2yNczUbuRmWWdYybN0l7SgQBAEaHjCAy1l///
NtFQd5Yjm9qyD31CGvaR0vICJovGp7f9qNmM0/YdEj8Qg22IZISfWcd0jJ0C4Zyauhqo/yD+SQm4
qe8Iw6Gxd7RBYvc6dO6dMbCFw8csKPHp1UbYTN6IURSEJRghEdC9gI+F6238ELI57WAyAwe/Jhxe
UmwYHEw744gNyzSQXGCKkvAU3Um09RdPmLjYkGW1a2ddyX1Gc+YYHfm1H1SA0UxidLwp1B7eEHmD
2V4s+A2gVtGDIRCmJx8h41mROKqxqU+FrjHr8OQop9BN2f7On8P/hCZrlkw2EO8hNQP3BE7sufbB
IP1d+R3K91W+tc6NPwEDU1F+xBBdYTmnyr+6Pd+N4XGeDOw3cad8OJQQQ2EOYcP/dtN0D3F8HS+l
q2w0bU/RXCmuVseE0bS2Hnpk/fyK2u+maoV+1Pmtlj/09A1vtynIOURPe3CcYYSze9A8ZIL7vM4b
QkuJCq6sIZ2p2DUGs367n6FNQFyBr026r5COW8WbfWgkKDmbSNZKlyUqK9Xw87mfZLkk+ZY50wLv
cl1MN1vKeR6wYEfKbkTJa7ox93tHE7XmfIje0t6+J2kR8KXcijTGawkg7kdeDS6dF6eRknYROA+N
yRISCJqC8kqW76+8y7Oy/dUzH74DLgGBUYYfBENjni5btMI9g7NQ5Hc9qF2LAwX7ooHVtdYHiZgE
S5qsTKVk/uyNx3UcE0zLLh8If19iyU+ztzPB+nRhlT+csZP8vgd+cFo3XNUGt9ezT/CmyKhYEIfT
86RKYI0/9SP35Znz4KD4gStfnPNSsLssAOeZE1T1FhK3Ayapub+J2zueDpyae6+qdRgOZShFMi8R
vI5G2Ji/nL5wxB0t/7+XCxS5xT9Od2GlOBWNfqvMNQzVImm1+2naeuOm2RL6q7UU+wGeBYw4Z6pM
kBRzR6RU6ef5RM1TfAv2QQnRbErd+/sRh5TUnfIKnO8YrRzYzlQl/WD64GBlo2jgVTV1oqpXUFEB
iqae7436GDNjSnm9IAylvr9F0uF6oEmZfGmH3765GbxmCFEQGDsDDxic+V9nWf2iLZK9+NfT63gJ
lxChTtQGIXj1cv1w/+fxzbrDLX1UvtOfbQnNLqy2Y8X2Pt4tuiZE47WQA+I9mP05AG81YHCAKpVj
LmaU3prSjnGyhsDB8e9/RSc+pjGteayEQWEhXYUWhi1b4/VEmudIM1lnlMi4cCO3iPr44LbuBNQx
pcREt7ZJJwczBNAivxZM9+6EPKL16GL3mz+kOoh1PnAeUxKBZNnvGRyb8XkRablgMBn/lw0c6I79
p5v5+0AS/z8EQiLszqkjb795rkLos2uYGYyiONfxQfUzw+aFyy2uNUk3zEXHnhu8TyI0e3o2Dbxi
aoWUIlJRgNRnwCW9EYPz+Y48xMbztDHAJN8c2mV675I+d8Xng578qbAtInlC62ZA3SwOjKh4xoII
kr8jFeuhwVUhc8aYkUVLcwG8xuW3EqqcQVPejW3SEGkAuC+S3PkdFjoDF0yAeCWyinZK2umJp3in
/BzHj2lYW1PDDsgFKnU8/+jPSXrS2cLAh/c7duk1k6raoqNPlVRfApzmJ/rKPgKxYTl16GB6vSxY
VLjvxq8L8ANt8cnEZUWNfDYExyPI+wC6cgWH0fQ3U4I/Lgk0e/rRZh3n8zCvo48SSSpUOdt6EyOP
uW8p+uKvUUeuCObhVATDQa/3u8n7KFL217aNP+Rx8ObjTthIUsuQCtDwkglkMNuNT49ugeD95hgW
h8WoGSSWwWs+A3fC17wcrBImU9uh41S39WZeOdCnkMsBXYEaAl6x/Gq+JogAtGwXJJU/RWGZnUIn
5DgqO0F2qB2fFDj3F/6bDBp7wa92rmbzNBg07LaAYAZJZ/n06KR1I3ErPwLX4ESOQ+l7VQXdzhth
qRfmomEFsN+4Awumok5PfuZ5CkribWO7hdrJnqsgpUbZr/vf9XPsLW4sZPdoJla5fETWN2mUxyDV
P4u62lTRZ15oV2zvv7IUrUp9kia/1wgjkENK03+ZQiQo8V3sRjdTMo7EEsfuw/vDo8I+GPB80oJj
79FiLn+bJkLnw9XD7ZCadLyxKSOIA+xqCRhJYHQyZ48+k/n9ejUrX3/Rp+xdZAFOsaUYB4g8CcvZ
bJIn8KPBqSfK/uk9rkm4zgAdAKnlZ5pvDyb/GKyFQUZlvahNSHo1AFLzjdU6brGMBiavh5Uuv2Xn
GswJpuKkYQf4DwS/Xp1TpM2xUX8h+R1Y3t1ZXoWVKVil76/Vpp++ZWTFi3jXqtXh/tlSGVK0xWI0
g+dB7CsDfwGMyMPlxLqGbcXMf+SaQyD3fhsizq0CMDOeRpFUxi147mGhgIc/tQ4nhrH9YBeNPE/0
ZhIxI4dGhdJ/EgBbXVEDZbPEw3CqwDhLvgxY0m0/aPgAyjKYWEPAJ7T0KCD2YptEUrqQUUqSpyTF
Bzggf+GSR491MbiY1siPIoFszOgvY0zjcqO7n4oQqba6lC6MFeDFrRlZUKszqqHeqmdzefo1/nqj
pSq5ATe5kMOcA+Way21aOcFJT69kgew37fXJAzgMEMmYua8PBDWt4jnepuKR/e9C0dA8AA08ITdS
DDboHwO0ertLywoFLKoeuFaWFzofsLbQUjlVTBvOn7t00KjElYmMzsMa9xS0B/KLQB9LHmfsNuPu
W56J9epUtYw8vU9vmdUB0hO4JIkMgFtyFBAKd8gW1drjEF3b96amrJ+5BvF7zc4rI/wy7MrtpAZ9
ESP3xDKnmPLnQkzzH2164qzCw7gwJYBPQgs7qOvjRGmNLJzcSGN19PYhBr4qcTrdGyZbfPJppvsL
i2qBVk5dFqBsPhuBn3v6d/5O7xJP0UXkIX9L41axB1cyGDrUJPZU2heKqSnbxKtg+o6KChEsQ+ya
EJjtJUxsa9yaEY+Qar1NzwG3y0HYx6pDqlTzMN4B0q5/TTbGIyZRY2+Ut8eeRvLb8muRsEObhdgB
sG7Yr8oHeleYDtRS8oF73FGREkI0AhEd1NuXvnzNG4CYpTuQ/DKkjwtIgzZwhrv9TtgTp+zl5Yjj
8rUOEPnbW3blolXADD3eFg5/SqyPmzNmqF+yOpCCRHvYH7gxN29eVulxoFUzCl/SoJf6MYPJmdXc
cwBk/GiKI4V4N4FzjPROvd/8lcDPhrFzqJfa0nds0zdwr4BrIVRLLvLNFUg6WMK88b6RzkjrzPQ5
ebo4Of3dsPlnHjVF3oKgeB0+oovt8Z5Vua6V2byyM3R4aKT1HtFvBO79nZUbbBE0LC13Mxo3IZ/3
GKK3Nm3RGxZOmityRFH3XeDTi2i5v3NIb3HxMpZH8z9Q5Gt1dNsa7LUhc5J41l+8ArR48/xK9ccQ
Wpg6EkLeqyx60QlCDw2CJLt1v4qxft1f0lyrtOvYUjYYC5HegIVkqzePvxRBCPs/WX9xpD0jTyVt
/slRrc4Sc7h5Ll8zfiziW5HqMISC6gQIMEBxT5lrMytGqk9wRZyNXEIqERr/CY8ttoq/m0LOG2sx
0INZHnMNoXi8frfsbEFPqkgPMIlGfB+ZiAMD+frq2+ztHUy+6fqk+f3jc3nLnNBKOr1QV1AaaJcl
q0Dcpnvw16d1CfmTbgt6VbYewBasQWn5VsBikMC28D48IVYjPBxnxqNZANMBVbrp88WE0nBdD5ag
WLsujFENofnuI2H/cykuu7UqtIorxgCnvKkqyJNW/5DUCzAoM8wMd5dwr/RshiBzEmLmqt3XCoO5
1zSuYt31C055U7SNcWM2Vu/radl74VeDi9V8oxHzS9A8nm4NiyiEwe+nldwl+DtUx0NlAvbN+hIu
BBG4N+ym8mwHObCCVqrTwu6vCrMgcZXiwoBUtCGqLQWPpuUfoTU1SQLK2ssckFkvFXvsTLIQF12h
VOoGcTzsKMynCmyA4reY6laJ7jsoXfVz3QQ/e0sG5g/Obwo3Gwc/eDBnZlnMOswU9fmmyQJP+ADI
6Rf2BmzfCNkvU9gdY192WVMURbFdbi75Fu8RWWjXLip5Hwl5cu9vJmpeKdZDyJsgxDUfek5Rf7bD
85e5sxuhWJ6itOQUIpdOFaT95vO8LaEXvqfONDmk1zGh0zNXrbwWhEvEhR2mhGF5Mv1mwMm6ou7s
LvzAgyfhmOO8r3c2jPMXwuXf8IPt3V/6EsMQ77OtirAqn5OQk2wJoUaK5qJF465vR5Eg2vLWxsGF
+4owtTSSdkV3kZlBbuu3JN6wPx5/cemIV08HBsukn3IsMFHeQeAG2jUZTHgo/2pYKrr9nX5cBuDV
hPF2FqeTH3G7sGsUWt0hhDLYPSnNfPOqUXmd6egAbbv2UiBrQVfKPXHkclhA35Gdy+RQZuzC3Zaj
s5ifcbWglZspLQ0qZpWcwqZ1jJ/a3VyIp+BUqZmOmD1vWMkQx6zD3aBHodmNA5MSTq8gQxRo21/n
1VCY0JHwIBmRBC9/O4puOsqw3WLwYAkhB5F2vGFejCqdpxEcGhtHYHu+Dsj/U4jP+A0pEThn0rd0
mslMQkkv5VBjG5VOrbGNixv+m7YEoMf2jpZ64rofZEhR4p4JWtUrKsNSr1bx4wvMaNy1Ch/AxTkQ
OY72H5upqDk/bdRjJhtkZGk4571CNbDut8k5Gb35XjU88id3hOGeG7+4FYzZ14jTjCjHiQuSKmZ6
573/opbCxenF6ohoUWC1qBEUkwrF/p7gytfDB6MU6M9v77odFh6DmIDAFVAoABDenxQgDKThuts3
wlYoo7AJyC2ZXN1JNTGANy9QgLn2sJdquMQUqlzKOtsPMH9k0D8OOiXjE+1HQtg0gbe6wSwTEkYA
SamHBrKSQNdW6IPlvoIAPuwy21f0R8rszFm6kUjektfDbnwDNFtsl60nUR9MU8AGvtkJcZKO16A2
CKnGNOmhOuCShbusA4aVBFCVMX3XAJcbY2CUeMbEugsut8aGEf4HaVU1AqQ9UyMYFvNOyVlscEzB
+r2ZPwhObWSATqywLtfxW6GyIRp5QDR+pYrcpRbb3+Tlkp74rMkgmdiTHXoNppVzYhFHUXNlTtpt
7AwgXUzXD1O4HbYr0O6hl8IFY35zrx4OKscUdpplu2wWeXlI80GXxMVf1SMJEnKGxgUg6f4bn5ex
Aue5mTDAAjnVWKyqtAs2jkkNTqTvRDMKJRf0XRMQd/5d9KT5FLFcD+/e7dv5XNNmJHIOuGgAO14T
l+uYBCipXtR2ylldJsgHQ0JYrtVfYdSqgd6wf/9rgkNBEzp/OuK+D78xUn8jsApIGTuls9LLs4+D
GbLBvL3qZsq8uVVpT0qzjPPLAJWTEh3i7xHEi5B7OnlYvXUoN5JN1268Sqr02XndfIQY+j9e85qF
XrPACUQwcSaP2CQgGIpuOBx2NT+JYswr/KvTm6Cpkw/fptcKAuMo1DKekV3JzrO9NamSSSrrUIbR
Y/BwafFcXJdPnSJyd0p7Q40ednyO2+fVSfQ9zLUsVIXkdOMLmG6OqUhZri/fFxd8cai0qZHUP1tO
EiIq1lxXme6fTI9R0ieyhWpom2+tQQc5C1lw7hAT+5MWOS9nvfd7ZdBQ5QF9K3YIP2OTG52VA4cf
MnBzQv4i48xnJjOgnXtwoLBPXzpYoBOVXKogw3cY2FJorExGgQzHSe3R7mC/9sbiO8nPHTyZzqqu
9spZ/S3XLoV8Vq4KNXdmU5/gbUU1EmW5auJca6wFl/uHAN/yc8hqp7XE7G8/sFRV6B/HyD/rTTP+
1+i0W0ftRIqz3R6RS8C/UNXb4vrcBVs7cmyUwj390XHh4//V5cU/tUOXuhM0bJWjFnMUtLHqaaaL
WFVBQKFxKtjs3MMvbVSFxURiSsvheSRX1n6qtmuxsxHLmu1ZwuZf6HaafgvEcub5v8jzfdM7NMz8
+cdNYYjZwqPZ/RgcOdGhQgA+GeyE7pNPmkV1TmjnV+HGyEU3zW78Uaoo5+6ZHmmf0vIekAHDVY1Z
pv9g4v/9Qtanzj75MedGJ7NLpBl6/zszOQlddIGss58qb5XBDfV8kSJv7gKa0Zr7ai2Cr0yzccdj
WnNmsD6NVjJ6WzHKpdDhBR4K/g8/M4WD72OUE0Rzl+PXbkrtn0KXmhWYLYGIMvKlVzFTPcSxQiGW
cdxnjrRYTCJGgPOTHr4/zrkgexV1cACef4PsBcs+4YDKQE5KiKkZOjAdf71jS5u1dA4J+j+NQXzC
FPeGTy7ZjPnJMg7J51e5JXp1XNayJVw/i0x5qqWfC+He6dSHERYJqdbFDlfbaNGwMfl9tSQW7rst
uxWkEn0wEp/D/cqcw6EvJ9c6RYc+DBoW4/rKHla0ZeEwiw4BOHpGIiXRcvl6aAJf7rJghTEMlYqq
Yl5FilBDRKJ4B+1D4aonDzcIDsfWl0/NfjQyCLTt4i/6iXbSJncic8QWuS7QS5hwb3Z/L7JZqhZh
ZyDH/DjON2RfbBMawPr9TfGsj6/fXk0t6KcdZsnWeSsJAjeT++2yYmr30WdE+Srr1sHQvrbOL3Ir
Ov9oqTMEa/lMuKqV8jwwFczg9l2pEO3CxhwmKEMPsuXRmMvqxSghq6Vy+1dTpeJ7JR/MT/CUoA2p
rIpnNArt84TJRGDn8LGG6hl4RgxARuy964Ef52bPQzaHvOiABnf4XqJ1fuyW7yt3zuXWjGvnfFv8
E6qs0rvhB1zImzB6ZP2iRaWdqQSjwasHYY0li5PWBUCSDPhKU+YwZO2XvTc7mXU21jiDOjrJyyk4
mAvLcSVP7JlohKK4P6Z9wdPuLSOAtqlfjSl3xDfFwENXi/9YXdyna2E+I63pcgdJXX7ldOG6Msw5
NeQveAwX2oyXvWMuT4f38vKYkdtEv0o1F2dLhIs4SetsAved2MtVNPTlDxYDWSOOmU2ohTZy/Vrw
qp54Z59YNg4Bd0LCNX6TppYOHpvhCrXv2ueB72GEWOBV0MUx89BIEDy8gBRbQrFmb4d3MDPVkfLf
u55CoQSeVVA0O1EaOnr92spPsvMcZ8RdKzg5Ck1R9f9fEnrVHBqGugjB7I88OahXi9BiXPOgm9/5
2dfO2HFayy1sMYUJN0OO4y7i9Q7tQ5bYvEO1DxeFqzcQt/ycVNjEQ7b2K0OJMbuHNO9yBAglss8u
cy/2KO2hhA3FBnvzSmnTC7m1c/ivODRmB+XWY0aU8eDmbFQTGMwcCt3gVf2QNzyeLGOiuxfI+cWU
pYwJ+umSGdUauGV8Sbj3GzTzumgCnpqzAI75+Zn0muttPtpWJE/Im3RhRp3MRevNcNbLO2Ntd7q4
LSxrE22elb2hzWY/eth+BHk1+rauFYJqpSPZ5VIbN5pza1m7ncTLIDhh5wC+8qFs2ZiDXifTuqRx
j9XlT6TD/idgDWvSuFwA6Wcvzg9aZD3+Ch5W3fujeh3+Hlq8KjRp697WxH6rGljtXlc21Tb33vll
Fh5CdrVE/chJYlBwTfrUNlXEaGR0QOTDUTFOeIPSIIvj/0R9UtK1Gih1rxKPMfYJIvLVUXSVWFBB
KwWmkTRKaviaZwfblDmanfqlt3L8BP4mTZnCLvpqU+K4rQmx7Iw8NqZxTrKgcJdMlrvjbdnYSKJE
TNNDIqd5fLJj4pDjhlChaO+bmFAHhoHf03H0IhChW5w4C8LsmxfOrR8bDUzTjiTejMqWxjE5xoux
jx+tLjYTRtva2RQLkStGA/BsuTb6Bp/MODucS+R9mrNYHD4QXZvBZnrVAI5xOLUNf3ZPhnJ6sSVl
6nH7s1Hq6ayeOiG0Zk9b5BRT+5OkgufN9tMndU/JKc+IcxCgWpY6RYUIs4ZKGSlIieGjvpMaZhh6
ca1InXT/eJ9k0VkQRJ3GG8qbT9ht6vaZDyDwmKEtupKpiPrfTE7tC12Hfzmz2CFhU+vsDatZF4t3
Sch4gU/VV/YHQjup6q/XVhFF/0eS0SU3wlouYyn2dXIAxG7/IxnGdis2DbPodtEna+406cfbh1eA
hjCTG/640awNUi79WXVQUksFIBA+6HM7NQZfOuUvpT7FUCyhHRxi+QJgiMNkXCghQd7pjZqy+FTH
2cAohtMPeuBwEYzLe5MWRorTPCdTKWAlCJP0ztpRVADS3IWfyCdhDOQKuWTEDhMzEoVIBIEs7KOm
mvpZy05PiZHuEjJpkzhBqDxDWx7IyAcHdozzVqO0SD8NDj/jUQhdKNG6PVnCKhNYBHUA25GMFPa7
fnMrFBMTazO8GBRleCpgOSc15zuUjwu2EHsZv7TuXicvy7+j44WxM1+wk+LkEcgC59yNKi6OoZzg
tHR45WqI+kgIoL8lrmRqXfZ8J2P2fjZBmIjcb7s91ueqQNhh6xt0klfenfsxE4HG4dbKGee/omPs
x8NmjIGrgB5yhPtpVtUbWcncyiQaJ4FDkjfh1jxDlOqe7pb5mM4K1q+MAPYyLrvt7S+XNoG6IU0T
FasSdfL+jvn6aGVhuMeO3MsRzTIBhLiyrZw13Dyk0d+0WzIrQmbMmQD8dElqhrRHU8/LFIJgxS9v
vEBcQcDG1Y2LZPjQrLoxlCMYT0cZfpBV9rYGrfqlTMNiYKnCL/zdZwen6n9GeTkrQFn+oiroOcjE
9PD2xUxcCm7/qXWRC8DqK26+ynwweoelZJdZ8LDZzRAuDlZxYEQKMYnHE6WQQMgLSgOsp8bqqxiQ
5Ee3XzliX1tiLPc6mJWhkfmIoJrt4E4nC+rK8ROILHoaiX2gYwi5KDY7vKqjx7tkjyy3dXCvK9fI
7fBObvi9HoLbuqATJEAOk6i0PZY9q9G3xjEorANKTr5WvSfl2RXeqkv8CZf3J7Kp0i5cdMmlOPyH
Y102rK2hnJPkgWZR1KV9zt6uWjjysquWnYG3eqVkOH4yATPYqKcd9V4OcO5hRH0ZiMN0rxJMtgtf
xE6kpFh7bhKe/WAR61Y1TLfiLtM29gb9dRswHo0bkddPSpVE03FsExhhf8GQK1HRmK+uyaEza6m5
/NBeedCSNbnUADAnWegabHqnpeAAywqK8Nn8/PsMj0zpfitvllbtfKiO7IIv5cNSG3TcR1QFdmmV
P/TU6AxmCXumd3J363LhDL/U2YZS7M40YLKcBEMnMaMY6mMPKTD6KWF4LdOfzCRwrJJU2KYk71Ea
NBsON3qXMYuB85GKYpgUTS4Aj4d0cVVYqduPXn1YrTaqfTkxR30a02jQYOAJi+U1yBYyHnu4edq1
y/jliLx6m2zhSHbtoIYyCwtXJa/dlPy7LQvSY2H9fdydDxpXZio0+j2GsH6fLq1hRQobQeu4IQdr
gbtsrlUFFe9lyK1iPu6mZJR+nE8jWBzVTmiR3Zc9rvP2WsCQJZHfk4LFgw7PO0Ds0TpcKwSUzBow
DXjOfNDzuSvy4WmNxolAQ7DgLz9yBsant4IC7f+pl3z/oHv2lcPBJ3yLsqNDRhnVujT4441Nrx6H
WQFV/gGPhSctcuqFSH/qxwqJwp7N/+2xjqAD/+NqAS9Y4DfQ/aiZezzP0lGHREIXhkQL6wU/i1up
WIfUuPcPX050B27h9u13cEhs1lmcNPRm4jKclltHRkiz0ZALOC+eo+MjiAuEXMqYUEIkXPDK1uS1
abiDZx+2fScOlw2C4LXI1H/bTpwAyu6a/s+q5lXQVE3rUQAx4oAbFkOTiaPeG0FrPtq3vs/P0isR
rh+S1Py84ZLRWlt1fVIsZJR78A0iuYBPEN0Bb/vsMK5qlY6x5C24qelMi+r78rLknNJH3qkk0OxG
XNQ8jKn0sDFquo3yEPJ/ABs2w+7j/EqN5FJamqjbwdz0F4x98DDQpV6fzKDXdUIiiBLarNEiwAZj
QoESqmYpqwmDjNPJyTC/5aaKTnRh6GDLMXn2qWF87ydHsipWkTeEYbpcDox/HJSeLxQcUzNm2MNZ
962CaRZarI2QHcccKlmeGvyWVvYKN1pEP07JqIL8hNEMKhbfYIlLkbiH4f23KdvPA2sL6iMHWxGg
pOYdNe3ytpY+o4/uh4nQYJ7E/bg4gU49hcRh7Rz5QDl2pNzFC5yUQ8b+4mlnNeEDg/rpzkSOuCSg
6aW+11Mx8jP7G5Qj6Hu0eUvbSsh5z91dhP4DpnxYq7JlNt9RuarZSCmtmb2Yjral0vPdggtul9Hn
vZD5Em8Ip5wRb8UUIq0kZQih03UUKNJhAEOkatoI3atWpnMOOGljXII8H7+5T7yN0IJg12iM1/op
XtNxHaFulcWQ2FoWKIJeGSmPEVkIK0G9cxjPDfWgY6lgQqNiipEN7CCTZVQCIcYVTH5XQcfPJkPP
t0l+LR8aTfvMf8EGJq04Q6f6tJEFlqAT5MKxsQl1fzmlDPR2MOXaFD50luwg1jSX37gydbOTZFxg
A9BFKAJkjAJ4R33eLpZRB+jGhDHaZXHC/fJaO/YqtKSbVcKFGiQ5fUxlN5nIiAaSoy7jhsmh7ep5
KPqeKQiqCDHnO89dGwBN0jRKKGalmVUJn2U0emry1I9cNpvKzNvpZKc//lLhy3JJBvjbQzHglQIH
x1ns1kGDptVsM/9dBlJ5ffuL2KAUHlLFjYc0CNEqiVLDjCVLgkB1TDgFYBJwX5+WDEGEXZhhnuhi
FJkviJek1zbw1aToQfU7hEYhwkeEHZmvX4sZUDRVeTvKlr0VJcT28znI+5z11PqKDuGlnKVElsUl
IqyDtenYKPzKggXe6I9AvWRRtPycg0Xhww4AG07K5fsQMiVZGxjRhWU3W/e3zXfyfTNRWl7xkWDn
trpDPefQN9N2B9vXnidEpqSpjWEO/PtuF8nuJgApsN+623FJfnmkMiFCWpwNVZTMzvi7W5uDS1Bs
rJifn8YFbLyJEvAixWSjiUln3l6GDjZpahBzLPYuTwfS/wWMJkUlpM41ljCdgIWJQBvEjOiLXp6G
fD9QdiJgPsUw0aXQR8bT1pFIfM9tdqtqli4XnmeIng9jnT4nay3HpAFjAnPgYFzDg1J4INK2Uwlq
/KUWLnuTR78pyiRM9Cg7UqPPOiz+wtopYDdcVOYjZLqmjN8Dlcbi0ruQMKz88Q7cWpJuM3F6JJMd
fF9BfFFL/UGanxEVAn/18+OwtogCHeLyuUuJhuvTlwIKGCAyyzqJYWa5RhaZp8ycZxAE75tnkMKZ
htNzuFZqTbY3Itg+Hvqijc+4wjzrbtFHLxYOKPGmF5noN3HtGyX6TWsTgz5wuscMlArhAMH/tZnI
hY8z3ahm2zZU74/cUFqipO+Z6WOV+HUyNbsGB7QPPp5dC/qwTdm5wGr8gnCfGTw0CFHwSDGp6uAb
D8TdAyCbMxhYt5ajHFl7QxwR1IMFa0OapYt0wswz6TNBQwi/bE0Y6kCV1Nbh7wUPaiabzlPZTdy0
ZYIUdA+9Y3yFfGY/9RPbZRc2hcnUg0B1rDA8My7JnCr6babhPt/1uTGnlXQpH6kbYsygwmyLuA2p
EpOAj2apPeRRWFN7QeCDLwTfvCJKhIxjErcrziVlC++W7CqNmTQzHygzPUarmOEx/C84wqNFjU78
tQIeAQumhetMzp7I/4KWZLGwFUs5Y2TMtNBox74GE/hqjG22WVl0QYVQKpN0o/w9oY5vr+C4uzvQ
MrdGs0J0o2WLtqfBEPV5CMt/w6hHkZSVVYLphcDZWAeMxza/6kx58cA6F3TH/Dzzv3ekb+UUS74W
+FN7ckTygyWXJ6VRkldLcjVkM8qwMKRQaYqE47QEQLa3idF2/XCTQT9BTidTYosqr4Xl3bphcg7C
c1LW5RtKWZl4b+Jnum8jIlF+/t5ku8YPV3UOTDZ+O7nqUUQn3adI7Radtt3QBAZxCzl+9E61FR4J
1dklJNQ8wELw0fRXGZHoUP+hO155ISpBKjiq/+rn8iLpPHLxYWDI2DIK2rm/Y/gIp5O7yRQOp9pd
SbTL8wntUcGm1J+2FoEbGW1rXfAHE3vHxv6S0nnuBJeAJjfJKYDizkWFfLRRdc51Y9U1Cu5iH+S3
cmqpL/5bCYULWfRUTIYwM580+pbB4AAmI/Ir7HLFHyvpsM3Q7mTzJe/YKtkZUN1oJ2FcKcsnJ6bv
xH7ucOkM06rRsATQoayBCPD1ICkXZbGEyAGbGf4qvwD5Sqd+0u2mFXTmi9IFNDIBFQKhYb1y0nTU
b6LxsSgrkopDdJYX6gm/Z29nOs9ZhcRIzsmAjJ/Ng01YBQTWy7/HoL9Xnw+XNs/GoeIkI2hdLOGs
JytSgYF18j5OMoPTcKaOexV4WSlcNshOC952eGc1ieX+/7yboVsiJbEWksIbyF3eLy6TWnuk0nom
3CpJwsGSRpC3xqDFZZcVnzNtR1PGUVjap0fJDLuj+oCkAgQBzkp3RUvxWW+kkhVdftagXIAsoPWC
HmfMkLgipO+SdYKMglH3UthOH3zQqATFJbdOcYVDTKenfL7zlKy+nCLn9a77My5plW8ttCrVL98S
LxuQVhfwokfetNSI5yF3kqmngRPUA4RpRF/BY5e6lXu+IWbpBZovfDfqPcnJdQfmNVf1Sm1hGVbc
iAgqxjh30/NZtGmL351Nlg+R3QfSOSgI7AHKuFj3swdGbIC5Nrmb+gidjnBeuJvk66v1lFoZR1KY
SC6vFfms1X4ugjBTMuX0fieQkYcpliZykonj8zaJv7PUzQNl7sJfHhe0MA1P+nQzqGoUzDgZNE3n
KUor5XoYnpCHvYln2D2SN6pU8+2SFLb942jh6VGM8vd1gb7rnJ+d+mgETE9EYFO7O+XIdcwk53AX
0kjoqTxDfsevwAEWQrj/AJST10o1dMpLuEznVAKSt6Xqgh1jYB76bbjH8wrpe1UIG7hX349R42GB
AaCxlTvBddWGAcZc+Sg2KKlGkxlDx7F5tDo401aMpau606O3r55DjxosjsTviRqZI1N3+cHFQo3U
W/1Flksi77ghm/uRYRPn7V79/sXT8P6GT1T12qJQh+GJGcIZ+PXW7C4wUViinu+3PQhexWUCTE4X
Ue7va3M+868iMZGoQpfAw6lZ4aUhFAweoxoCyK1EZVukDTgYv1kzjJTsyrinpnbHb2hid5Ju5CsR
GhJ4CSZE2sLFKo8fdHvUz3gKeG9Du+QLYPS/8cfV4RflyTctkOOdQ07JS3R3/kGN5IvTWDm4CHNE
5xv3N53F2aMrPOI24uaPt1C6t3phDOCt2jj3f6tBr2aC6MGgZtNbhtDdQDIr5IUWER6yG2B0SlYA
LO9vACZhgxZ0z1Q2n6NHdbjrtf37QaB/lE2UfKXH+syiPmpCq76DF6uNUAFqm2gBmhchm+4cOxR9
0M+BvlHHcMDKc4HuF38cZhtk1OY4cuHgUBTQGQ+O6TZYxaL/HfuXEisqdhKbQ3QrnirXg2xXbvbE
j7RF51UlljB7r8/6UYcH4oEqP/nHej3xmmfOiFMA2lGMgMumx2Tq+Hqjuyni0Tz66LE4JIiRbP3U
yorTWQSE0TeHH1NLJkIjxK0OiDCfIi//jOrOPBOsA87gd4xQdbr9PBEgNMybrxYEv+xH5b4N7jOr
cnMPvA8VYZSlUGQmoYWiTmn+vJB3UBCOo0V3ox/HE//WBpRrttdEtrmnVOrts640iXfIhM/yb3Xa
tL5XVpwBCXs08wVRzrtw0dP5rNv4NpU4MNjGryRVUFiFtoDvUG5M4/7U0ZMC70Th9b8Tdy7j3/dt
XeDo0qTOFnjDHGfGBhpZEExrB5MqcbUcGYrYdyxQo45V15Tk3Vj0teIw2rDZSMt3Ul+WU7A5MWrz
fkzd/XBk8pvNnuoDGllSL67R1U9pGSyLkIaMfINKPwqR+080fOUVm6jNA8Ji/DagsfvhTG6ymgcP
uaxuCp+mPyg19ZVODPeulZSOszgAHZTTo89cau+71/mLCeaX3rqQ6/oqzuWFTDvm+rKKPBkuBWTC
nBmy/AcFpxJx4oGAiHJa2Wx0A2rlzDh1Pn1KfUl2q28pPU3TO3u8gtLYTUskC8cEAwcIacVOeBt+
JVzvLTv5FLwFlBYwVD/FsXvRUSxNATla7NCc5XsMLGcIK+7QrIUFgjU2JQr+gEHCeWhmQGlcdWqk
kx8eSljAmeuF+7DFGUKNVE2OjGxnTNMcky/rPdPV7LqevKAXPoN9RhmZXLmV+Q2JXgO+Fz9kyTSR
vrbb1yi/ZU0kifbssbA9472BfFStqgy1xUcZclgPtKt8BF4zglmYRHCTS6izo62NhsAPJdWPEXJ9
NBF25KVkw/8WrGfImNs4kAqvajHi2eZ40xRm8p33Yey0odQ0qDml1Yx3RkCIxSXWbSQbSuG5wRBG
8BSqfLyZBSI4pWGIrZLhnSkwcZJQcec0Y1VrWrln1tMaGPMUvAZWfy3MY8tqLToDcPrb0LUA37++
tcRNYmN8V6Pk5gEcnipZoNeSvsFL0wwC4DlQT7pNTVffcy5fP3AHNUZlwRZ/8z+XLLWSfmG3c80V
yvK8mqhyyfusT3L4CjlaxYqW9mFVpNa3HxwwnCW/WhBGmxYXA8Tx6dZ3DwHxf9ODn/bPj83LvE90
CfJA/VHjDavlS4GWWHtHuY/MpjuR+Cwi224fntizwQiahQ2kCac38A2EUqNqqDgnVro7rEolkOq3
FwRWMZVCdjLCw+ncBFopUjfEBuQN+JodufvKBCQoKYzhhWJdtCnlyxmljkFlT5yn2W1CJ0TD8VZu
FIGLc47f1gDZoRdCwmNFLnb3m+oc6nqOmhYggBL/iEQzZWwW8LQhXfFFLPPTT+wzPCDZy0czC9M4
HjnvG7F2myV55xfJGB9MidJsOHtungMRLxulxA2IUROGsVdPbwoSiP1zqtGc01wNIMbxYYqFdYaE
/LLB102nhK1/6fzFHA+4FcSNvRaorA9Pu2gU7hmGYDO58NZQzxZOy0H4+0wfhBFUsj9WKc6POv1p
vLge9hPhripJrDh0qv6WGsPYO6vnY5ns9whop5i2EpAW4B2DosuD6XUw62L4xR8o2cO+d+gbdKKx
HEWvDoaRnGgRdKTxvBBVy77snL04auHmoAY1lz92UWbc1kxgN89HLay7VrWzyos324lRxVGi2yk5
L31mUtWq5IO4jwdxu9MC7ad0Q0nvl4LJkQ+0pGb+QWaGJ0q6qp8tlBbCciJX1293ifFh+A2AT6nS
t+g8C+3D972QUjkWBLAhzxWMVdvS8EtjIWlmpfjPzK6eTStPqYuz9lVPVb0dGWR2AOillKfHMofw
alh8QkwSsJ7qcWAQwAWKRg6pbYcEivMnx4Cw1NwSZVCzXAJ7/hQbYh6wf1hZ+F8j7KLbKfUNeyWh
YdX9aWwk+8ezx0q1MhZxk+81B0m7JhJK+4yEr0t235O6C6/s08Odm2baG/XEf3GgZAZYU8Y11Onm
5PuCfDQhQcVOzbUS7NWp7NZlUsergA0SkR1ZfX09Owphp5W0MyUxMUDBXFiXSw+PeZLH4AnqvdId
2oop/sN5eFqGLPx4P7SvDTeWffYkFcN/v1MkcFvmrIt5vb+Pg6BpRMKfGfKyvuFtP+XYPjI9y0C5
b76pHKGX5rnkZ0H2f9mQaxADYxcBhGm1Fo32f6k42Oe4854Nyj3uXhiXm4d3rmj4NWiTLSaDEdR4
WXflrY/XE38aLOlPUJuwBI6JczuEtGExVHN4qJwXqW389YzrZtalk6/8cAJoDwkpAAvkyJxnKKvy
m0j3MS2prAO6cOmZ3khYn/E1xnMBr1KeoI4qffPRoYf/dm5pAXmRN/4LDAr48yEzckdgzoI4bL74
Bzzr2rDa94IFWm6yLK7NHa7c4t/EovSPBx3W5NKzIEfS7N0eNu/7VqzmTDjS1GX44SM+QYdSV5bS
bcLcjz6mZSuDGG11noteTIp6LqYIx88DkMr5Fpv24LogBvsMkiO4dZdZoKMJH2ru21PdQak+v48s
nmFPO24/WpVBgmIBW6fJ9NnlfpBhxsH6Sz+4FcD18kpl/cFYcEIKCL9U6GX8RWygSG5kiQJeMiw+
Sr2FQ3/9YyaCjVTZICmv79oeIy34Jc/6rx0RwSrdiygQTUHyuNv12VV/yrQglIQP5CZLvmO86j+j
Afl5PbmRNdDgN/TG4dIFahpAnM2NzCc5ck8ZpZhmppBnkmAWsNJIrpQSB7cSm1nXQUzpSYUA24Da
yijEF3SQZ+UEejiAtrv/E3lSJDEszROVMhb3bVVMq3h/0sO3qaZRneYoVUzLTh7TxkQcqJj2vz5C
qWZO7Wh77Sm4hoQHa0HJgyib4NyqgtNRXGhyNyNR0c/+sSWMveyHoLR2XY6t6Ev/WPoMfNvsSsne
6oXzG1Z+3DVyDvG6TEEn0Kwx+7qchRGIniro8A8eeTpwCitMoySRTer4TWHTWbvmX2WJ9f/2exSe
YqSBAt8SJvKNtiHIrSUaE5wL+Y09bXxuDkDZTd/eMMWDLWxTCYbCfwulSYSWnLtYHAyboKsLv7nL
cFlC4J9ElRALr1Q7awkdxb3ngd7IJnC2IHyfLoljvWuW73wS/YlX0Rt90OllEH7jqBRRG6+zYL0T
8Mmh32koUQKeyIghSAMBLNZToH+jeb9YRrWkzfoMEOVuny/Cyam07fOCbBKovs0mAKwBbDkEoTNM
TtI2D0deQb3X6b65qfeQUWi07PIGPHOabQOlZ0S+UYW3wPShO3MwiqdWlZU5KmEZsTEcdLYcir2N
msmsjO0YUHvQkWDAdjjXik8o1IcUy13r30e+zbF/s1jIx85Fz48np8i/FzswzCIOKxrAqhsMK7Ar
u27w8yLHeE69LvS4OYXlG9l0xlWdKt/V7DIQS3BDVHioUjixXktUZZafZTbC36v4AF9aOJU+8h41
Gu6krmQTXrHwxjhGYdvKjrq6C/7F5LDX8CHOUdmA9thcniImUi3GHJOd/fo6BkFIXS5xfu70XBjb
xo5Oj9I14ft/aderO2+tdibBbid9Nu4gjYowVj2n5V538MaRnig6evOmlK6pqh139L5wEkah+3mH
LH8kJZ40XhY+KzfW7OPpelrc5XcLvDTQI+v7zRYNe9EMab8SqQOwqpq6c/XntPgghxrW9tkJY79W
rPEpfTElHZ7XxUwZtqo5+jkLyKa0S4Kjtfcs1SMcSs4UWyt9da0jqs8wsWRMG+0UpClZe81bRgdm
B7DkY6Vb2pWEcaO9b/6GPQ49Y77QE/A4hXAGaTaGi0OVBzYA45Tt8hFjCD1G4mvJFZ5C8E43wQZy
B0DyktdZB5skSaleVdK5zhBu7JozvFQIs4kP2OhgXnQbATBJf6fna2tR1g15yRAtm3SY9aig0CKa
NoFRysC9b7+O67aatGDss8G0GIkyOMsOSu3Yr3VwkvOrDgKSFK9LOSNDdli+nV+yx/PLw1O9d12i
yVjRStWF/rjpTdGYVSL32xaIEeFo9KcpxoqnDSZ2N9rpegozCAISWVpBHMapI66pQK58maQqeN+x
u0RzknhUoPKMNQiOlxdQKMYmGKcnCeg7B0kx/v9HCtf9CuAWYdeRcnvV4O9m/dWfGiXp6hx3MerV
d5TNetsGppzH02lAyew1mhLWSmguepdRsZSZpM3f+wrfHOBmLtUG0fXHJ+kW+pIVWEQ/EVdxWyHw
txlvXpifz4KUYNDAf6QKRXzVfvLpqhSeHTeFYCuf1agXLXHQFdcfnusZcIpmhEOx8AT3qzXvWeYD
SRbGDvvhGizWr2YC/KQcEgKZuQtnSoZJYP3ou8Va3rOC0V87VTg3HFL8DouoCd1LFPhmgs7ElB57
97F9ygYpQdfPNHQFf8Oed9Qo7Nu9cOjDJIx4xmqTyb8eDIk2hjMyz+PlG3nUK0eKJqyFpHEKkVI7
5XQyWcYHha7yN65Z9zdrGMRYPmpQxc9yRptotbSYuhhDZ2x4Qsmz+2OdvJTQobbKdC4IGdi37zry
uD8fT8GOP+mCzD3QekAaqQ9rlyOv7TBEWZbNu9CfTgQ1PDAYMHfmRTuszsNWyJ97Mvyoi3IRX9Nl
xIJH8eqq/uVZPYgiT0LchG/D59yTt2G5v2DyoVN85bjlXbR3J0OEg00+RfGjchryd5j7b3wOjTtT
tqnpDgeUgwkdlJ8mRmwAXVT95fDGYM1t5phklLUEcyFYWuppw1jMOhHP/Zu/FO3xyoDzHUoxMxKP
YCFFp1OcutO0qRx0qipaRFCDEcBIgmr0QImjdCpiKqCAwp2lY9X8ZJy9U2kGnBtF85rhRQK5Udv8
wHhKD6UbIwXlLGbk5Y07OMf1+izglBhcMIv7VyBuwY1znu+iCEzKmOlwbVTyjohofAXUPErydzOp
Wsztopgo5l5QYZNmHgjqpu8V4PxIiBP3IC62ZsshlqbodIKCgqouXoQL+ofYwWyeF/jiIVWoYz32
Enn4WvDgYHnxZeAdalP/ZW3he36sMy8StYyhUyFHZ4H3nxuEpq4VqYkbHsTPMPKizRKkiF14vTAi
X1Hpw1+8xCWupMb9nvqXQFTfeiF/u02c/b+VMB98nRs9DvpIDI5gx7WRSF5Wl+p90yo0rfFfKtio
pzzzhLeGqpaR+cJ+Jv5Bjyji74nvJGD1XeZudKy8jvP9/xsPKv+rLxcLAFq9utwl+Awyu34+J8zL
lcEuW7/Cpqi+IufDiSY5vgTJHTnZxIeNXaLQOlSJo32Mre7L3/54AVswpy0gc+TV82W5a5x7sEhv
22JA/72KKqUTKgalajhWSThUaWagFWeQovWFi14sup2Dzq4DwOXZjL2yDcrk5Mg2RwfiX+z8NZXp
ZjidMdJl4lkwYlD7ASpKAm3YhadF5otZt6yhGDhX/ODiFOC6auezg+QQk+MXzyFP7Nxdgp1Wm+hJ
AQkYgmgQVF0e0BKKCQby/f4jMxG/cExupcZ1I6JuNfNjr7H8gaxzFvpFYlprgPnjRXOYhh3O7qVX
TJDvBfEn5iHOKtFeD3CDMS1IT/jFYeMXV5rf5fex3KYeUGgLfAt1qDxrsCLOc6JLQhUdd+mBURYA
IZ2tqDh0pF41upyFXPD5ZoYlvrhhb0W4B5v3w6h+6W1J+0N/r66LK1Oy8t2YUOjpMstqv5LTI4xo
abqqjTXfulkT5ws/ZJ6l0bppgv56mDjx5RP18PHKjnRFkzn6WYK9Q1y9HuqrOOPwvbbWCKrrETd3
6ClV1sHWxjAClSW5S2SiwnS+MQlIjOWwezTdtER5zbQROBHba/z+u0tGXEzug4KLD2KU+AG7c5Cg
CWjpumxrsxabQ+GD6MBpBDZXjG0raqHheSSdY60mH8C561z1AGa0jVLVYA+1f2qptPjttjFEK1GX
+eW7LsVakMPVw0PkP/tuCFVdaeoAK8rg/pftSx4BzEzgsDqGb2mS5gw2Irfs4zPI/a1iqE8IdVuL
zHHSLvWihajU30tkmh2u37D8DeOIB2/eXb8P9NyaVvJO7KYZlvxuvGo4N+K/Hq+NRSx4EyI+z44c
dBK7RakyUUbutTNMzEi2FhGvohrY27175TfCU4gc4orc718X6bImjPRjLLRkcZRCx2E0mOa4r0Xi
mVuUowGO4U8x2Vzby1WaKPb5lWZRznwKBwhmrede37qk/f5hnGEmR7IfHQ3frTwQlEhGYmy5rL22
m4y7YqyeZiyUrrb/4KXwYK2nmGFQQMRYtAgC4zNrZ5vs+MPTlCHU1UI8tVcUe+S5W3X/MEsWUJpk
2htCBKl4Dk3Vo//vRp1AoTiF7LsDcTXM0SytxWB6yJG0hkEQZZD6/n66PONyvvro0TsZrg0sQHqu
YKCVmUfT/JbT73Om2WVimKvPy3dvHl0rmdECcZZbBYCnXoSw6VdHk2dj26OL8kr5YI/YeoPUYFj9
Cb9v9lq7y05VoJz2EQIEqQKaXqQczpb7Gtx0ko9nnBMUuAqzG3t30JTk3J4W8rakFoIMGcG6zCxk
Ril/bu8Ud5y/FapjujHOXK9gaQFPDZmhqDt3uae0gbsZu+9I8dVVWAy8XLNfVQMaCj54opfClh7t
uMitKbH8MrS5tnBPNNLlrzcOcp3UxvNZKhPKCCIltxf4pb0qGcduZf3W4D4EpTsUKHAjs2Y2ACXB
FyRwn97RxlqqHXXKWYQnbnq3DapBWp3nYEMSe2xf/++QEUF8dQcFqS5hA2G2l2sHmS2yZAr/Kg4D
fzXWuX14JK+/Wu0uCRu0r6QmcPDESSKOFQ4tlD2RWPz3oz4vmMEAcFwwR7EVGIIuiCmXSl//2n08
pycEtXhqXfeQnCUdndFwCIfRWMup8mLfCJHLYTaa/J2ix7IihZXaokIth59zJn179LmgLa6i+oEU
k6b0yaoZpJljSQcZn3wIXmo3cd/y01rx8NNuYcmI7xjVI8igKSZQzPLBOqKCdvXlUWGxATVBeUlR
VpKgpjautEUn2HgSxv2Bld2HWfAFHBKgIt/GlFGmJ2sEg3WUmWbmYfjsAAX+IYsoa2nVaVKoGstS
APXl0Q+oekp778BTzumhwGXnF7fThNM1bh+bSybZeZGSlQj6fbMBwoH52tmR4Q92yR1JRcYKjHQd
csSwkmdZcVYKLBwPULc134RFXAxpPWGFum5mABJZqvgpHTo4Xw3nx3GcQ/5lega1Z7Fbtxtdew8f
NCAEp8EorgU7aUFU0H9gQNjl+QcPCRq8gjuaxrOgbpXAtY7vkTm28cPjsbAUcqjsZHztAMIoLnKz
i72bkMzc8PJbtKYZR9VKDBGTxYdaNK+7N7S8NOqYMCxvDtMqkDJjNxyVdrqHwJFO/dTvH7Ul6XYW
LiR+i9vDnzF65PRLzTvW3C24H/nVp5fPl/3oBwpkUCl4PgFCVgywkRgHrR74RbRs8PUIAmuynQpj
gsNRVx8xhKy3+lcD9860EUBH8s9dK9w0hjhMam/f+RoRs8wxqrD3puIo2V/7RrfWmu6eR/t/eyCZ
CqjK4dn6+01W4xhCzZQeHX9V2gVrE0eaKdS2H6i3uo2b6wR5DujuwI1jo6wDAHkC/xOG6uuuDlyu
fBI77WJB6lcLWRqhOwPJAL1g6OeDsT/KRqxRpTAisx+s9DM09fFpcXffWXSq1HC5BMatdpHxIXcP
rlPt59e2tgEPp+THhsZ/YZ9PxLHEv5z+iKUNs3jjpbyb+2HjLFpiOG1cnXzQBX6a2bnh+/e0r3Bd
JLwHKyz6amFiMqh8NnfOj5Gh2Wymk7R+QHKgNyqH1cfCFmuezTYXKfSVDanOuIEGv4IHzdOkQTjb
hVVib48Dz+8rDchQcEbNMmavJCfqyvWPZI5WXJ/ZMcsGq5ulZ1SdnsCG/VZSXJscAZyI71gLfehO
BgzHxihsaur0AByyb+VVU2PMBKqwkSS55qBg0R/t3L62CsjBMZaRyOYo7FxKPkrI3ZZdWcgi1S1P
XtnqCSZIYQVBOM5BzLwlokZrqm3DS/o2KeGWBpXrwsAJdjTrex68/f8JD6cE7R3dGDWYOEjGgn2j
iJ1CegTQMHwmaLUeefVlRu0HfcquUxB3BIDiXoSps0QalmFo3hgsFmwKocCQOkTCO5E525Z4cKXS
k5eA7g/gQcJe0zUuCiVqqSgqM5MLFrLKz0qHmA+neQyfH+daWro7xHretPilGFzPOPILHeUZs6It
WW0wocZWQK0c8F65vjzML4Y5N5oyHluTyjO52WWnz7PX5lMQEqporJl3g+W4Lhbex+++Ui015I17
2BDFkefxrkvNF1YMIYFSXBzArj1Ap7Oou48BkVCqiNukrg+MkpzG0vm4uHJ6M9pcGpCrC1HTYl+q
5zQux64mPjJfe60B0/QsrojrO++1OOjOMyby6eCaX3Wlv610Yz+G1UWCXcaqVyLgt3AtRa44w5dJ
AKKt2r8LleJtI32Rg8pWIQyYMxFlw2PUeGyk78GSVDG40pzNpQhpG4WQJKcjjaSHYKfLCpOq8Ods
ADR3P+xJnRKZAgOIYo8XOHK0+hnVi/r6v1tNTeaY9q1QZfS7X6Of6CS/yDhwxYGxJE1O+C0xmU2a
vf/ZsZcEcXXUw/InaSra+iLr0tHKeACSE2p2Jk3WyMea7nl/I0aKm1Gt1JGZ6V9/99mIkSqszThg
yTYrbdQh95L8nATMLo7tiXmYLNOREzjzKVLD3Bys8tdvs9TnazrcmZxmwAtIAmtsvcwlkxWfKakV
nIY8Dz+IZ1s8XOO5HV+mweQaDihpxjx0APnJ1je36bgBY+uRsyMV8zphuoYN3QH55AOzutd9Kjq7
Wi5FajI69pXjadYN2kNfy0bk92JbT8/JtFF/3YJPvoLVBTaDFyRD2CDsbhiOVmd8uu9uKDG5GKwS
yZJs+EnhdXmowPpdW4UgcxdI6RdiVZrBkEY6GBWIZQ3WxnlAAsfQluLZXkHF88jxgUG4MoDVLaE8
e5BhUqtWRsc17GTfbKjMk82giszke/aIEvFE9ueyanDlhmIbHoo9AUtT7iNuSNflIBFXpMA//NRZ
YSebOIgO15pchiEbhZFWkCjgjaS8tH1zudjP5toqhFgdRxaMxCXdK5BWFuxiZuHaMBIr1xcpYRu4
vGdqleJzpXq2F4LHNPkEaZ0VrqUscBze7K83f/ST72pg/XzsIrr/SYTObdWwLrD62R1CvBkgK4tg
EcgnfMZGDrOCa6d9IC+cIvTQZIkI+mo0CMY9m2xyl5YQALsJuV2c7tiJbhWeZnA3N+w2YKzosFxO
z2I+leA/UmKWPnPKRbFrcWdtgGVIwQArG0e2W1Uz6ssGttCYWxCvUzZHWQ8tmY6CgJmIbFjoR9sJ
c/QjslfRN2GgG3rpxwuGql7frb/JesdBCFvbreu9oHzDbAqUdCUgJ1NFvuZ3VqtRAw54iKMTfk5s
tMGb7zyk6T+0TFhRHfQCHQ4CUbRKkivNsWEuezA7nXViiKe2mp43uCvl4f+Orln3wvG4SkzH4Rbd
cwjRvCtz/bXPJul7H1TJpYqUKR2AdXShsoXC95Ico9H5O8fP2dtFfxPLB5dBCeHEBqoqSNFhBI5e
PQmXqBFOH8gESP6oyYSjs/ksrM8ghyTk3uALukNXLzapLq5vnnlBc7TxJ2EQgJzVd42VHXuvYE5Q
qtIX4iowz6iMAgAz1yoTuNiiV/hFnlxRazAuneCTCDYx3Vzpkmovfx/jxgaAEcfTx8YQntM57tt+
9gycwxn7JnGWUbmggHYRGvoDDC9FkJ/6aXZTEhHWuR0l+GZzds27UUSO3yIA0F/dV6XEFvMpTgJ+
9DR4B0BMz11UZdpE90cAPkArQBQs+mKKy7JCSeouGwTe808Wf3+s3E+sRAb3ODUyGZZ2SqHsncIt
vFV3bamQzv9iAnKvwL44PrmvpTtwgCTpur/q+1CcI9edCfTATPDMrLw+84i1Y35rdLTl48kbMLAa
NGHbJZt+XIj7LosEGHxfHXMZ8qSpymp3i48/1A7sx9hUlZFN2VV+UMOxLImN4d4xonyycWyHXq67
yJhXyd81lbaE71+a8cdDg64kk5J61lzWtUYJHL3YLmurcPvLoxvGS4/I4eJ9iz/69zSRqenk8mMm
5vvV3gI2tspd6jb7RBzhLkupbmpWgYtyiUXBFvqv4xffMSuXEFOvGuH1ZcBoHJ1JNbndgv4dgWZS
5IGKedVRGXw4QRqg2cjeS2woeM/dS7ZLX0UEHDL8yFtqQjO4jghIpPt8VeX/SyP8yheGei9TOmWW
zwaUIkzw9Uv/Go/DqZXggHA+fi3pAGPQYzmFr8+G0zqgvHs+xHlKkFZTlAVQRKXb5Seb8yqGD9k/
il11aaq2htZKEw1ioEvBBDywe+E++jAYtR+5U/7deaKBJpBI0ufY+0+CpLQI04YB+caJBThaSA4Z
U54LLQdeaBEFclhJ8HbFKYrV0YfrRMbmbPFJ6bawkOjFYa8dHUdVFwXLAlweCztUF8kz5RzPZjA4
n10J7fx899QRZ9uP397lUhoURAzlknyd+yEbkxrf8rp9SHtsnPPhhjUYXibGi/9D15hhVGXJ1JJL
WyOkj7TBH/fkPeV2PWVotSm9B0NB/Bg7mOStUHcIlqShL4IizKTeSXKpyRRucSGpshN6PAKbsDWY
vV/LamYSX3NXHE2snmyS0ZxBgFFmx0f9BimVgJ3W5a7ucACWpZgO5+hVrQMOPjYfygxmz5ym3BzO
hZJbss9q6G9AsbCRMlWy13WsGWBEEgH1JNXd+fGuVVQ28VZIPu8t3m8ExAitK32MAyuZQiR7oHgI
/JJm42L4IsG0g8ioqDuY+DQ+KQ7MbuVIEfqHHM68IklPvc2J2ArlUwdpKbPYgCKBl2pLrn0B+Z2X
0aJQ2WMfdkKE4iZdZp0Qg7arfew6ewpgxTS7aRio4M8pE3Yu8lpw8B1dRwjMUaeZQBCALMeIHlgF
CTzOhAWVVcPpStFl07kCWrvxPULl2vbpGSfJ5Jh+rqvNFeDNR8J07T/z5ERVu14pbGRUvqktF9Cg
BclRbayWnDZFOV2Sm5+z2XEXHrjWhycbDpUE8uTz6RAVUJXCBA2t6QO4f13SDgg6MGioVf1rGo2u
CM1GTF955GSfslw/eggiuC3X8ql5+Gn38iJgc5kHBlJi5fvAiCjsVYPdGdtM+Yw4Eh5rmzHns+01
t8ZA1pg0d0tVyBxxznC3vXqxon9cf1ico8zEa222Sxuci0nl3TQpHg1XX80RbphoUNt/hL5qEkvq
FBj9Qw9U07DxXEz9ABxC3NBzyUwBER9G6lkghaOU9QZqZMXTo01bx/ywP+wt9tKinq2I7/juKcbR
iubBb397JhSVh6pJ++ILx44mF59EtTEDV05LCvQm68pruSav2359kIMzGrcZdmH66MnQYqsL7maP
Llsk25wUuZaVzXS++6WYAb5F2b/uoin45YkaU+eyY+p8ToxTnYDTqU1ZGTJd6BOhAmjeGLv1ihUl
l//zxZbYq5Z4a/2Jv/VRgxIz8IzlY3kYRfRONz1soi3poo/JV73AEdvSef0VkifRrUiMX/jy04wM
nsqLuN2M0TgJ2hMSpDJTJiSVjPF1QN36gccfEdWZWllDnbtPfoehxYl1dahYpPKW6osYMbc0RFRx
Fg6zs+AcPgCQ/JhU+Rnw1WHaAyblen489l7txv5gUy8TGMBTBTxiSIY0MsbgyTHpcElYDID/HrVJ
vEXruhWNqHTSVy16qj4876+hOleGSO/nFcotZ/zFxPrfpWA5XrV/FRUxjmrnOdvFh0r+OpunIPqF
lMGN5Xa94/GcTI2dWNyvM5a/EufV6e1xalnZYRbhcKDf5qbE/2LjaxFEWFXvGVE+HKRGlApsPIwa
u4lOeUumCmQ1HyQWAP73rKy4uu8aMB03GDMO09X8IYlRi2NuJ4NQhna1X+h0b+Tdm6cS43DzBfN8
Em1VwdXbC5RnwJ2xD7FGMnV6YKGwTFQo9JOzfzjAjSbVK78uVTX7quk1mRILYmG95kbx0v+UCGL9
mZC3/DnSrcV2tDeIBkuYI8/jHgIU3/QcEMzxpl2JKBPiOKNeS5HAogD8sAgFe04XbnuNN9c6va2V
saql4b/Oz2uzJPqRQnH2ENmGUlvuPjZ3nNbOHxh82pYRGLR0pc5dX0SZdxcTENFYe5xiSYD/hVM/
fU+FXfkhkW3pb2+9ouNOAGe7Omo/o0gPVD9HTp3wXvG7wwrrAhQ15NxFInktslu4BmKSh+R/gWQN
jsXlQQYwkUHPkR4z4f8iCPU2XCdwyIzBCgzw27St5wPiyVKC0LFwAGj3sMz1YIUKPTwv6eOetqBO
Kp26YbvC/tHo1hxdmYsl7bWTpy3ZnHQ/fB2CjPDrDudlejswP22T0k12nJRDHUT/cPSGZA0jzMlJ
qH2D6747XHDhKO2j7EFBqMOednpxRx+FFZ87FJazNwSrasxfzU4l3V274bUOf5VIeeGy9PmExQrZ
LPOLzEG2ZKAdYd3JGvzoXI6SEDGn1lu0EdUvUx9Sf69os7gUXNJZK9j82/YKKJk2BBfnWL9RX2gL
j0J8kG5ydNPByDs2pwkiDeCEwZrrgbg7m0lfLy+QsM0sxhRF2mmcMKq7e5gpSxwLXrpCQKsdGl8R
ZwlBn97vDWO5v/eQi5lkrACa8Wqt7ckF2yCoWbizeb2XY55JarnY7mXxrOYPL91mY/ECxFem9j4x
0mbGlMsQhJvKoSaL7C7pNzaohPc9exGowPN4rrLsOTRgiD1JR1oJhKXgPnHQa94+oN4GtwRCInB3
EepwH9Ob/qiqDI9KgxAYc+mqX3tv93iZrULluKriObzcQ1rahabDiNBFEQm5664mpcYNojvDAfW0
ZVLU/U/UuWZ/B+GaGU+OhrPbiXZkrAou4B/ndQ0Hshk/j/D5Vh4NYQ3enXF99A6VhNRehBxByhnF
VxkmnQTz2hOOxPJpmt59Tlu8ObJXX4ZuY/hO5B9F2XDEU82yq+3E2CPU96eAksduUjk6UwFlb27O
dDOFRyGaUt9SwxM25nrj7/sZEHWfL303dInEjDZo+nkAlmj834gadhDtOyscbblngrgC5hUvWHAF
zGRNnmReHwu8U147uLfHBVmDG1AdvZyrhpGXOeYfFGm4NqO7lOEXbhF2CMkTNfh8rxkqrgNB3KJ9
y5SgVvptiDeU2F0CHCgvB4ck75syLjMUi5yj7z10t+rwS6w7GoxmCe9qf4+KtYE47nCVpHVPCfN4
Bpz6yVrRQerC12rDu8UOwkKkb6+QDjjvhZ89V1cUr2S5B6wmDyPuq77MjY9XNiL8VKZB4YC6EdZy
/F/wP+BwxDpPoW2WQCW+7IuhwQOcK2/asNs4aPKRrZ87oOK3NHghTYN7/ZmPODGloCkMOuTbFEO6
CHy0rLsd/9OQ+ATz8B1CFx4BMrdY4jInPw4PF3wKV/y/bTQlSgAe7lPTCBsZz63elT4G6gk+rs41
rcUmLm8hSYcn//6cJs8nmitLrtxGdrBmmh7K/rQ2lyRNK86k9mFAp83l4v/raoaEFOT6nG65jaCF
ZPnK27/WB3B2Gu0A2zKubVEpbqnHuT+F5gp8mkX+0xmHIXKa7Zwp2u+rhqNnU/K8cPscz49jm9i3
B+mIfFWrwzQJqXI74GXNMdTOTnx+N51m2P+TaP9RDJBmNOVn5cfrQXA7rSV8jvZIimipBhXPywxx
NdrbWEfosWBgwKznMiciGNZr/pJvHCM3jd4YdX1tLwQUeK+km0GSa4X0xsz/XxrQzWA7uqJjaJK9
3aF532vO8xaO1JmIE5oa9hzseyAn4lrsYIK7l1/xee5sGmsx6oEFDTbDibVsh9ntOMI1J0Z2MxkY
yLGSIw3Lscljds0Puu7p0/gaW1TSKwzZpe7BW0oesvN5glcLuF+NwbCxnGgzrAjQtxhJL/UJ6KXl
CD68wbvVdvDQ+BuF8m+PqX3iStRtqklJmxtpsUB5Fd+KwSNuDxFLXrZPD+OkdbPKFHDcC2qJw1EU
MBPYV55gI2f/fherDkELhnnsmXScLmcz7vETuU4aChPkDqe5LNbniNo+T2wMqK+kdC3ywFTr41sV
pwn0Irb1FQspBBQZszT76UctwVBWYJLChs7cXcjUPL6Z2enbpBTgAhnUFWdi29cEG9j3hWpmgUxo
XoHnYGttWTQpSNANldjbaRp9N4+AVSlCBX53oisNcuKHXvwEkKa9AyXc5N7be9WyqguFdYCxeeJA
9td6F/TeeAsCGCzDsP2f6jv+x1FVCeHqozEq83b9lc283pYEIoTBlslvrZFQTwfgi8vFP4x3NN1p
K3wvSb1sk9TE/BiBlvx9YwQQTdzaoFBWRF2buzb3GeAWa0egf4z91ECFtQURVFPTIt5ZcRQO8USw
Gn+DNq6YhC4y3BmW8yJXXG2JO9x0cur4xvm8Uyr3SiXUhQI6RVZSGpkgwT8pQydrtFwsjXY5h5eb
7gKmSU4x1u8mo36cRJuiUowWxYZyDJvkG+mmwMu4wwpVklmOtYLWPig4rnegcdlNKmXDOt+XfC6g
udZZ6pDEQDuMWOdivHAH3csUh5vVVqBnbHL/aP1So06/4lfBdamLjUDHDRjxXXbCGt+50lNQKtL5
wbkzZaQ1a9yOWUDyTBq5kN0eeh9twv1sSykY0dPlz6uatRxfXtZvrFYeBFZLpM4T1QfaphVHDhSA
ii7BCbg/g4ubiyhOi06Q49ACYmkqgNu7qyLrBRC53rQjdWRYRAjnvGsPCD8p8+2r/85J6cniXN28
ysT645FXRczjrd5BrzMoU91B4J24J/gCwzIWkaJRSHPYy41vKOnLrGHrxnLQnYPfpkLCN/Tcwxk+
BZawXNmeQIYFutdiZqBK6uAWTxlCkM4oO1wt16pPUEN6cdWt67N1j60HgXtZ3t84cJQQOXfD4nyg
12HLJNUg13SrJ19On0+XzkszDxTHCZ5159gYh1klS7vKAwM1EvTFUqdpiJiVeUQ+awLPHET7ieId
uL2tOaUw9sSbcmar2Sg6ci51L9gxtbKGL5PWi2g2I1OLhqx4IO67dpW/HDrV48aWIpI9TZz3pVRG
KCf+PzMNIxW8n88cs7WA9wnbGulDc/OSWN/nS/mnUyuz+ngjt8I8xap7pmIPr4NjjbCZrAQo8GNz
niZwgMSlwjT2xTc0L6kcyliiehBiVJ+JqO7xoZoym9gIKmCMdz7wooOzTcgrIk59WiAGKazbp57i
zLEgvEWY3NDv2mk+D4rCIZmGc2kRVhVDDo0PtjgrckY6le35EKOHy22fZLB32KbbLC1OPlgz+kj1
h62rBPfAK4elCsCZTVjx+Yd30BNUan1/X6LXKvkRTOL2IZDcXsiDQgAPLTQH5sDzz8TMH5xfamZg
6HL3CZLdg+qyU7sOpSsj1zHNjEDohKPYDuyMRgXCUubUTGgsU/HZ2Gwfsphl9KJcbh8imHMHjtum
RhOLrcmQCDfMgrIHLdTpp2KbBs9mUCdKbF/Mcm38Xq+QQkzNQM7Q/TtZoSHsm01czUmY74c/WnJ4
2cuPTCK1pX2NufhCVmuF/zlxfLGex7RsXoiWhCZhOQRRafps933eJvmikFSX56zS8AbMIHcyD6LL
Eet5mVu3nRa6xgpxMBjgEBpMP9KQqh8IVuzDPsC7mMnZTDEnVxL+aSzKA49QuLDrFAYIPcthqNjq
65t9iBVOKEd7AJ+VxHOR4v9XdjCbOkaQiIRfv+70c6qK5WRNjHHBlf802b0DQ8zFA8tM3Q801RdC
Jkol4+KyvWCEPHxdb/+0YyMfftmn5QW2fp09gjCRA3xC0Te/TI5rhg0oBEkG7o46wyeCNArxAftu
2cTjLLA6Uju/+S/f3ha58pTnuyBi9ioqM7yMb986v5fVGhKPPaHETbZeL7/P+sic7NAhnxjpz5kZ
KhArcZWwniuVMyvUURXHVcPud0LKMfDiSdJrh6uzcY5rCo7q+aXtlTuLwmwuKlrunt1fdCb77Ryh
dpR4fBFSYi8xbXHyofJQzwRKkaqq34kIVrM1VnV33D/V/82ueK+NLBGCL08OdCNuvPEwnDz4wWBP
qXHtpu1JR4hW0Lqo+hUHXX73YA43HyKg3Gesg6uNB00hQKcux8w2tGKYs8pjetvlYMLhNmKCJTzH
4UBw1HTpqfaqDifLHSUcCxviRVoHaeOJftmPmmL5rgqrB/7wYLam/XBUjBJ4v3t4taG0QYgISvBl
Awl+s3n3/C0FT47IGP7z4b0Bk3ccHJRQzCGCfnWO5gqWzIleHbCXaWseGRFvT/Vo7CQ9kfLnLtyB
BI9QVb0fwrEepyTuQrxk1EZtSU7s9jsAQ4qO8XpAztlTMcNZO+UQV09PhywYM+sFYJ0TNsHzHJBB
7Eq2DC0uEO5bIw+JAjt0COeBSfuHP04KE9qVMk/cx4b1633u/QrrROpIydzD52LHxPR1iisFKUIK
T1qO3FeH5DNWKz1xXlWhrU1tXXod+wMFu1H4oIgTyBmEDSAnquRlVIhgUODgM/3mFYDIvktUMfi3
flA8LeMfjcTjdn2D/hPqkJiGVPUbB+C4BWCXXLmkH+OF7u53gdoO6dKsKGNAfSnPskdTtRhSDB6X
ZnRXl7i/+3F7EaV9SMMbpqe/5YaxjHxjms8bGEipo5jfj1ITzNpWU+tK72lHppMDA5oPxWpYL++9
58ovQNxjUdPOPbZdFG779Dkjn77yagywrlAfmFWnlraEbmlMWZ8D9vRXRmulQh4qJH8foFV9mRr9
DsOf99xmaS7sjmHLrgM+gg98Tt1+Kt5131U1GEGtLKe20bL8PUCO305rvElGZu0E71+VIm1tGTrG
DxA6VBRAn1CJttC1UXEz4zTvLjAPXD7FmDo4n8dstQzZYUdij5B3J0qphGYh5eqhzGt+tBHjYjNs
8aeFRex7RrjOG/CUUwE3aSBIDJbFf8EJ7Qh0xWtd5fDFKLpcAMC08eHcb7eTAwY8jFDgKRNaBxHT
kzKjBrUhtCh9oXUMOUj/5oe1FBzn8oQv3kPFKTv5g+LZYcK/eyHAK1g2OkBye8yehvSDCMSPXsDw
G6ulz3Ti87QPZZEAh8pGsL09mi5uzcAphc/9lxxR8EdrUcnla2vrVRy633M0+brHQwHtMypEY/fH
Hy27Fu7cR7buhDUqMyUdxVb0VXvEwSg5Rh3HCk8CSy0fibtK9K55Lhr2XLR3QKrP3sugR/KOW5+I
JjM65fXL6XFIe2K38eM4Ztmrp36Twl2UvJ/17mlHeD+IZEsrDvuAUa5HW1ZoPv4VUmLYDlFI3HxW
njRx65siUKsoTDA7Wsljn4jgDESHAeY+lctmyH8Mkg0WnxB9WGlKq6mzQsM4YExW5L/5YhZocJgE
BDevRfMFR3k7aBxjj1qr5NatqRwz4twnIwM7e40/ZzwdGurdDTIQIhuYx3CcAW85G8a3hIx8dXWL
PVLG6Al4kva1KpJXfxpUHRtTPsOx8MS1sAHgEIwPTezLY+1nKvdAy+BFMm3o7tXfavZ65856BERk
PUNsxkQlmz+g7pv7LC9DFt9xWVKq0f2kV9iZfslEFG/FwnSzjeK9vKw5PcCJwRK/vRpi17oYDZfv
KCGidayVVN3tNipr3uPOZG00IfZrifAhKNXxzyb4x+sCFMpyW5+T8gaCOMTlsWpGUuRn2ZJp/mFL
JfV33aFEwkqAoMidYyuBMRMDijLAJvNoO7L2YQzbdDO+TT7cI+wz/I7dHccqAFIaTATOwBVkqJ6b
isMyaa7ijCbeA4SZKImwTwTkXXp4rNqk7AhYfzmVaZfQrGAcAgx4oAxXa9p5JQhIf5mT/CDNX8/O
SQUFXf9TRUoUYCy508dgAJ/LlFJK1oQSfOZ+6VNuR+Usi/TUjnSM3E8d1eaYOrLYPTNQ9DCOkSsH
H1ipYrbJML04i6uv5VtJsX1193AONs6wcpqck3uLF34ro0eRQgaOlAQPFk2OXqjU4TEnjlVnGLtU
RkteMKxPNMztOSP2EYQQ/7+KoarPiP9N4+3L8kQ4CQdwud8jjmMLgQKeMRKX5v8saMbSVfa64QRZ
hUokgqga/o7yIbFb9vaYrkIg5VH3ryYpPIPZ7qt543+Yyc3B1Lso11KOu95JkehXVAx1pU+XI5Nx
FVLda3EM5SKRipJvXB4pzp8cC97/Jm7WuZN9veJecjEjtP3NeWvrfHupB1xNC22VrZFW6jGXxUDb
RqGHOzS58FYmOIqztWrdJvUAEeg6GiriRAMDoyadpmsfMDte/F8/TjyPhkzGTgcCFosFl5v0N7Qk
NdGNqJe1qF922gTXtwj9QI8AelDLrWL1ojMwwDj2Lbh17VW5aoXCNWaIlk/nRG4z9vBZlVd1gQdM
JOE1avEeIhXLc3q7QysCP2psePK/OsvKFpseUVYKLN6ylFrpnSSpx4LGK/y1KYFVaC2cHVyixELY
gXFbs7Wc3Eu4ioZ7oRrwdUehoWNthUq4JVENFyQa3gdKODu6n+iVEflU6Rz5l+VhEEG2LXBZcxKQ
jIlYQsWM4kJouUdGKF6OAD6rWbZKKhTxPk4BxkZ0I0E1H4EeNlAV6GEeVyBIDwGLAAEo1+XNXiuZ
k3J9lQJwsDU0P84nKOfW6a4NkhpTlyf2c4EiM9khLNMFTdrX1AV5WiO/5xynV/sr1HsX0BcysSe2
muuHMg0y6zjik3B4SG7WzRFqjZlJGgfExEFemd9aK5pDplVj5bPtFUOTNb46Q1724vJczJoq4Xs9
AjQrqWqul+I/26oOmjr7bXKMmWuyguWrNwGj+usRjrBg8TcD2voevm44xa03sm5O03Jk+ZQSoqkj
t6u3sDe/PP9IKu+su2+wXw4c/NYmLAbjv0htQtnwCJ2f4hEetmzdxd0jwhnWGrGNUcObeqIhb292
GYae/dZUefX67OjLIy3Axw8EhsMiV4o6XGIn+uyd8J/opVomrav5CbsSuwVKCURYvJo7brF1ntR8
Zcx3JPOXnzWLHlfuj602giPE8CA83/2j9L0wbkjH8anuhzhmPp9M9Vzx7XbHZqRrpulCGDzwrBzD
g0/BdgfmE0T2QMYjBc5EB9imYQP2z/E7P1L8LwLIBceRq2W62/xQUx6WwRRFPOjzTVCVQ7a0Pex+
nFifi27aHFCVSiKPavFYj+Kq3PHXggOIX0o368Z8Lo/RrOLrfloINkIsRGgD6iMfNMufDXH+jwMz
0hQcOvPpO2gznUuQo9l71mAnF1eqKo6xygY9lkthg1QazFZjcdJFc4UKZKDqj/CwMv9H2t4/BhtU
VQ4jMKGfDhO4i9ZhD+/kp+XMmkesYwdvLUqeDtCKvJSe70FvYuVJPZxxsYGuMVm5zWlbhbNC4J+r
QKhE1nNGqffgVv6LdlG44Ma8biVYWFmnwVuq+VFgHYxJxd9CZsqaxpuQhrNRZlb0GpXC01kblFmC
usfbuE/SvcufFIANRPNvyVDxkl5tvWXTbMn2+6uozclHiwGO8ua8jIPHBSC9k/QF2lCLMZ3Zqu0o
vfTuACXl6elWbjobIB8UO3pfAhP+9mDT3qh5StcuMr9Hyl9nDg3kaQKJcgNaT40uKEK7UTUSFgmK
NGB3eWlTHY4pYyrOteqvmbxiwC0J98e6m6vs/xnKWMyWKixJwXWnq/KRPX7kjyB829oUWqG8W3+X
B8rsMBlzHeJ9dMyqeLXaDtAqiH2mjQRkkiQzKznKCw8vgdr8dlgWQXGrkXgyFKRK0qg7xKOemCw9
bUBKHYO3QzZguQfYgp6LkdUBbcmSpJYogjnrxEHdjzhY4npRVPq4D4eq+apGdcgTTXMuQH7dnd2h
i6qw4rnsRnVzcxoQLGfefwJMzdUQ9Dify5pgRUukbgnCvc6vLU1R6/nHvwrYB7nlwoPruAzDTmS5
IgAuCrBKsx+DcVLxRxbqR5I/8qKIdNfDPt3/uQt2c9VcCuZJ57e7wV3eoUvnQ5t0w0IBAa+upeFA
oyLWzerz8tkTeMG7yabxBs/S3brKMm9ps2T0aRvekRKI2ppH6AJkELS8S/iqbn714q6rXqT5dXdq
qGgC4v5xOZ3l9pWYBXn2cQK1GBiRWSsaFbyGbS/AA2TW43c+NoTI3qO/X8QrCfINIzC6GUs5X46L
/yRjsfLT/wvSHuXHQZbd5vtqKwJzzjAwkYr9ze0ObTHN0PtqGN//rlpJlF1wKaczhj64w1nmRA8Q
q9Hx0FsWQJdPOpXSxytjzTQ0WGpmiCXNvPzbMhACMTDIgWqeuoUinyp8z81088xaN9JCuF0t9wOm
KvDjzgpKqRPg/0gvBb6uveTgxoh9pCF4A6OQElxqwS1ifH1NTQiVL+Qig2M86fPX93ocg2/mP5oG
sF6TvgzdOGSeXQZXo+KX/8Arw++DzkixsUs+lagAakDG+aKhdLnqlE7x/xhacLIleCQnc6UfqMX3
b5nApfUysMaoAU2n1Te9X+dRh6y0WeO4/zWhZR381VTdEgM2f3ija8hrPa2XfrZt+NYkQ7WdDsiR
fjIoXxXJ5czxlF7nx7QJRiy5QZBviF9Ss78ljFKz2HO+iBXQttujujQfWZKfDNgi/+fKUDOLsNir
QaHjEqN6kHXfE/EAcrG983/NfF06Wm1/2Jn1wrd4WLETVdxc00hjn6cFrVH80PRpwOgz/9+l/Oel
c6f3axvhRMwT8p2R5BjE9h2aawtVsLyBGLl3hfJoaKr9czyCTTK5jLYNWHzpjpRhwQ/aV0nKMHQ4
2kJhWtBZyR8yRfhCq1HvYBL2NIJaVzz7PJ88zAQZYk7Dwga1fvoP+xQ9GqgmkvwttznY0Zuw/bIE
z0mLI6XgwU05QtAYlIAp83YwKlg5IXbUPL1yQ2Rtbs9it4cPFa17uyXMSMcycpRVkPvTEZEMED75
w9kkeI9+vFyR351LLOafU8XRgY8kAtseRZIuKtUmkK3olrAIz+V+zmZAuinnh54EfVrHcmq5BKwP
N6zhAMavcEe4HzeaF6FHYEr7YqMrL9f0uiC8amyPkcXmI+nJY9LPGFALOTW8uLfz1CbFrwGyYPSG
VG90Sp3PwYWFjQ+89HR/TSH47XNrPA8WO5ff6C6Dt19tjYnzrFxBFYzMQQ9X9Zhfxfo5AQXb3SY4
MF6Ydwb/hUZy9aMex8cvOgkCMDUbnqsMu7TzRsicAtgGat/Xz//t0y7NzUyBJIuCXwizisqm31MX
Yqjfz7750D9zCYAE49EHD/8rBZE3jLd6cZVhcSXuWza6Co+bXLqhAiMFtN40M0TAsQVOWLXcc2HY
Jjb/UIlqCFaXQn8a/gYx5L6zwmz48OrqOQfViVSzIQadWlR+VBtjXXFrvYYlXp1xtLFcCfp1NY5L
QwfKzUipu3F3M5dpu8vrqXoUeqFL50bFRS8b8AAdth/Q1ODRbQnzzGrouykZkbPTDuKsl3NxfyPK
pGtxWkguUMnZ8Aw5pOQmGW7TNEk6daIKbc66qFs7Kxtx/lPWgwz69yhHxRRWU8HwzYtiDeerLnFj
EP81U7RmizU5LU8yc4JB3RvyQkwDQrbPGcVUbyDQsx0TmW+eMAoCas5KY5VIGJnyFd92rZMOgMNV
/KvduNvfKx8bp3M4rESPTtHqtp3AQdb1w30PAQML+3pPjIKxihfZsRVeSM3RpqyN2sdIRsg0rWzu
AlQnKidFlWAyP0obOmsQDmL4Dygibquusf/xizS9tRhZ/xM+hhA9h0kJg1yxKazGViJWneaL5ZCy
xIOVQsnyPOGJXvNHgZVGP5v7AvjsxSp3qHfBxIJZ1GomyPFrO8uCGYpWh1d+awwd0m9PrA/d4BTj
Ka9E4E8AUwzyLMI5LanKASQZI+SPacxI0SH1DQTPNuB7tG78YELacLgadrIk8nxKa0szdmAlZImE
bkG8EXyv3ytQLj5i03ywArG+IdOlRNvJyBK/7kFveUjYlBNxtVPrR34LcOAhBsZAhwfXoOHBxUUD
4MFhr+RXOEElgTOBHJPKXQ5MUTOInBAFcRMGlROM/CjMHMxKi/qnit5Ah4TnyeiRM+rRjeQuM2NK
OmNgjpkyLIqWqSs61CTv5nEu8jh41gP36HM0k1d+Y0/4j9PDLyHgABmjJVQ0NNGo5O2uMh1lL1+p
VUf14FnvqIkWFEzobbx4vLnB+0NTa67vYtUbyaEipPifw42ZPpb8mMjVbF4VfOdxWmEtTJJlJCiA
vc5Lgqmq1HEzB6lUAXFVMgyTXTFd7AXMR/u4pP6XqX9AttcAePwg3E7Ot955DAT2OIBTa2GUU++D
hJBYYEoL97AqacXKVOyoeEb6OfWMAF+tgguWn+qSipD+ptoL4Acgc7PCmYqaJFax/vjrlg1xc6Xu
MFM849iVBHdDKUU3xsRkYZ56hgicwaAr9lPSzRaYJRO3sAkojHLSSlDheImSu27NxQL/zwtF0Vp2
s9O5h+F1q0yqNIbE0eJ5z9psyjgEYWlElzHgPTd8aybo65bVldC89j7PPIv9As3iZYIrDi0bhhRv
IAbhaVUXaWKsWACLgKjxpVcDLXdGMdqxN7RUPKP6P30CbBt8DYlwEITYSxFzJhUpRsi4CtnouR+7
uOb4Ot2GSqzSk1i9rdnWfLKMWdWyTpM6jjC596Z37dJBv+bmnCuaVUnwTMxQQ/E/G83e0XEIU3AS
/vFMLVpZ61Sn8cFg4sSG8pQmSwohZrNwkNTx4/B074LgY3/3wXC4GeJftSlLkDHjqV/DzljMOfEQ
WPeiyscsU6Z9BgX/7dfnn1yeaVvZQVQpFQVE8XI+l/QSEGuAgUMeGuz/brRoYKPBTEPAngR+Qq9m
ETiWIJuPFzfrghiBZRb4ncp6IYBSufvUDmXRVPYvAQR8VK4lz8qbi5MaMnGh3rrMU5P4F9o1V7R7
kKwsEXXt+k9XV+uuW7nMevqXF+ZeJzYLt1h19RXrqhuNeZC/CKNEF0LK7VVL/OcM7FZV0Rxvy+we
fZ9dLnzed0aPzu/LtpfozLpg/4zdbLAdOvQur+wcTuOINy3pDafWyxwzCZEy/zHbbFJ6Pg3GgGAz
ROGDrNx/f9YMwFGfPnqgUsUMedgNTLcHqx4EkVAp7NpLVD/h+OVNlJuljMOZgrpbe6vqRE+kpqZj
xOP/oY2xt7KQZNVoRGuZ/50cQ3dddZp8k5UHQ+eMCtTmhJ487zRPjj78tRnkchtcL5NcXHiH1wNM
GJNrn/AbR9nwfMI/s/YIbzPEHDHNfuC+OkXR2NVUxmJvgmdUDEIHytJb1b0hR5uiqhVboITKVMa7
pwskdL3tSgjhNfW6j+JOHMJzVECp16PWQpCgweTz6mB8IT/7zk9ZcJWgZoLj7D0KEkslB8K/dyrp
1+JYKulZHi/8fqBwT7uv61E2BxHQ4sdQkycyjEjaTC18dFPDg/MzKr1xifgrX3g6LR4ig0GmkLC/
qfXheuL5aptt1fU3ar1MlzN/3wB+gPvQp+JOzeaywbIlRgsuQTXIJUN74L5HD6CLXuot20y+5anM
Zrs1+U6PWiGQTZbjdhEElhHvz5/6i4YCeF8jtGHdvLi6vuoE+N6j1aKwiN664vkQ+DonGhIqnZLO
jCnLitHkO6fuOyv9+ztxCcFU0Cjn6VsMyUDtx6BFsDWlxIZdUWOFoGBl1w5eFamXcadhZHBon7uu
6xwxheuEB664K8n139kpkomiFbTohYTN19TReJfIZWr9FP/OimmZWvw9vxHTUJEzHj8Me1G6dYCv
YQKyVU4B/vaWECyjDE0O61ev6q2w4DlOKijzmtGC22M9iw7aQw2zOzEDvsBtha/cLZhqzb7s/z2m
Xx2UNidWfA9VPxrOhe49mWVRhv6rljpRL260RGGhIWCKmJVmPuCTrSYt8/EepHyN8lBWqGmq1KpL
3yyDHZWdD1ohEPm/dXwbt1omvTmXaf6T9jAsQtXTYtSUeq9S8aICFMoxOORHPDkqQvSayFZwsqtX
+IheR7wTpE+u/FSxQNmW68SqACMz1oOIG5ttMs4ytntL5AONwr+qphd19zw1t2ePZ0hieCVKU6Ku
zKUyNoAT2eiL71mjn/HxH3QJkRJuta/Lw3knuAyY5bkK/LktCcS8yhSq+t2Z+NOkjFqlJpvgCkVE
sq4UKXK+tDJzzcFSwlb8t1TS5FwmRdVB5xDR+C64Bx+aMzROFDBHm4ipHeENEXXkBEOMffB4QgYZ
kL96y9kTjR1GTi6ZZJ0szQesCUfWQgP4bUup6R/ObYeFboTUYHCU9rzmN1oJW335173Cw5u1VsqP
K7bywxsc704l6159MtVY/aH97bVSFll7Z0blGa0fb6kwaQjLcJE9ntdr8b3WnXsRcDMH2HPflutP
XYOVsorboPWBtcKrDFXQOfdOACx2P4eUp+5bF4l3tMvvuoLqzwwUPiOm1C7I/4EZnHL7Hxjlhkmb
ay/lRmqa3ieyQAdPhEA/6rtWIZha+BOoBUi/uzlWMI8azckvlhA/ohHncOBU9ZKDAK4rPJqSDfUR
iykts7w7BscvNBapXo74i/2uqF9aTC1OHINRFimRN8IjYt412yb1uutroLeMSQpGOvg110oFMSXo
PMCmosKsKZsJpWcUDjXD5kFCMWei4AzbMZiWGOuH1xwCRmA3f1zHbfz71wrRZMeL8+VzeqBYBaIL
nNSSXQ5OqMwpGO7YLfaEFqqb/Z9fWHmDM+5O989PxEhfL0MdcRne8moS40ATZpzGABUncJpm1WGW
y5olbm8hphotPxJM4pgjtHpMBMiToFq84mzzYtGTPftJ9WEMdjGZIIf7Y1kY7lE8iADqChkEtbAh
pE4lVA2bgEs75Ub+JDivjYZLHZuihgQtX4skFGaSrGlFazjQXtbSntX04Ld2/UxXiSWeQhcRNlyy
3Yk4Nfy/DfVn0OUREzdJtcQh4S1SFcPHym6w0sPcKtOo2UXpyUKn/NlO6MhH/PY1oO8mMGEZ52K0
/7ViigZMiK6YUMSpTNRBaKACddakHVi7UQZTbY+2vmENsfoD6TrTX/9R8C5W/IZXIbqxR2sIhHQo
NhwXEy2ESGY47HswgJnTuTlVuuhSBMc3Io2SD1wsFYYghhsByzu/JD32Ffxi4DZtp/UPoaOGsyYv
sus62H5tiIYlezxnER0vuBWw6f2Ux4IUgqncJ6zinL+4ia3rjbSdVJTsCYmgtFCYcnj1cSgOuvrA
AdapYGkMCjVdKlD+DZn1HfJIBOWZata9vzcHcrRoqsR0IjrwtswiSe21Piv84BJ39i9Q87DnWH/L
X3kGYwzr2PzsBgquh3lOeU8b2CykoPJJ8kaJaWyxcFBY8dNKGgcf1SgIkXEhEqpCDtnaVAqdAr6T
EtyR9OOmEN0kbGEkWWVnxBEy8ehg7niPyNH0UTCZ/FSveEIEHcXme81dAkevP1SgxxJJi/yUVTbF
RNKYslIlN/xzg2rzWTSvsdayDjifBVQY+8dkBB+hiIt71D8iIDFP6R6vZT5Z4o7pYLOJDcNhghmh
2IgUPoeP4vbeNjk966vsLfFs/Phaq9S6bengRTxxWxDsZIjQjctne3x1yP1iPacgb7EGHD+H3I47
LDf7X9N+n9Rrk1+lCyBQsBJ9BUeJhYgX12ojiOaAavQXblbKMt3XF6WAg1NUnTGPjqCmQmtnww+V
0iokzgxCYIIJ75mRqCAgBHASC7Jn6UmkiNH/ASI8+EtLsgtZmg+/XeqRblaSRkjGHEglhiakst3m
qfxLUOYVPwVO9ny4GuVdIOFuUqx4j8BLN4kAMSVArV4pPVq/AWuY6AX/o232kfT6M57fI4iV8cm6
2WA9nbh8unjHGr1COzo2IF3E8ji9USGyTqD56C/rDgW3f4bAzzJk+D2Shq0NhpIYhZYAcXUwzD/S
Fxtw3H0rLcDceJ3YLxu0dcYMw8GuYBNzNxkkCU4NprWX5CJEr2eJv4SESMBu1V3s10KifdYkrrXp
x+CJRFfUlDnMe/W2z2Mw7UNwRfAkiKrCIucpNuzLsMzp6VsaSgBEPOjJHS0SfFWsIOQsj4ZoEA1Y
wcj+ooBDybIpu0dqeQLj7CtObVdT3eoCftTlUl5MbYfLRvhET8TK69XIOymvxKMoHhTws2xyIggr
/co27i9dOvw0YUqrs8PB7zlQd68Hf/Fa/bdoVSweQW3AGghxVYxeZAyOG4GZZSaf112/q2C+bqLp
z3sR9L91ABmR+vA5uCDfCQzOa2OcQ69f2HlWz/jAskh0FqXizsDQ5uqogaCKRn4JlCyjkBxEY0Mb
EQYdJAJZQPQfgrWCytQf2JPSxuA0pWtgGmAABQqtdv7rg4wWGoza1HLCYJA/NJRg+XcPYxmOhXs/
f6pQD79dp9bO3wi9po05jlxBK8zlsKpwhQe6rlPP29Rf+1ha/QjLWFe2ud9zIJPYZCzWeTDLe+n/
CgmRq2+b5G2qrtu9Jc7D+BG0QASOgKA2RFI14gRMS0jeOoB75z8YCkvBzgWj+tMEZCLUh88ld9fh
fwiKYZMUS5Cpyi3sn0PlGBptUzKDIFl5BxJL8D7CIHFG6x7h99tMvOHCD1f/VEcJuj7nz4gN1dEQ
VvAwPM2e8Y3kkDPvSKdoZE2w5HA7GLgZy8Pl+oz4K+iFpBvrN7HhbwDP4ehxzR3dYLpV0IaKoEK4
+eVvD4NXYwEZjwaiNydBseISEtxs17pcd0hllZAIAY3u2S2tiOXSVbp8/SwmW26JRnCBmEw7fvU3
HTwC97xilgIbIiNsmV20SII45Aq388mhhjvqW3PIAjTg2fUN0lDVuOC9Pf/z0/QA3V0W7xhXGImJ
WS4cNv+dmSSXPghLbBZsdFlEDbQ+aQ1RQUr2kLSf+9QCijnmhkITN7KZD7wfb7SZUKJelNNgEewM
haFk4qRWaJ5CNWLtgr8QPs6XbUhiko6s119X+R8Lou+5lhZBcpbzTlbO9mxdYHB3VsvsfOXEZ2ev
ZqZn5No1iqvEB+/H/AKSWNa29O2vPluwknJxQhHKMY3t8Q6834uuySwm9g52rxPDy4gTCXEQ2Gmw
UTN9a5p00LxnCoqdMVALQgM9Md5xVwaKFYK6JQwihrpTIVVdoNTicepUm0MgmxHl+IvYDj7faEyO
dXJPXqt0RhQ8ULTlc+/lXCqk4G7L62assNCJzHBVBGRgMEdDSZNDuQrKPcgaH0j8vEVG2HPo4bMH
TvOH23xfalYHOlQHVzWzuU1BXEpWgRgTAEfItK+Wj75wQRSZ0C6r6/kg72mQoR9rBr6X9HJPh+sj
JrU9XNgXyKKf/IWrrPc9OglBMb02Mul5QZIK3n80QaV5DEFSwBE4uBVClB/v6ReQWenkTXZsk2O5
Sje9l+6z7J/Cv6yTEC1MfXVGYed8nBnqAcp+dqDoLYdgq4QsTJ9qfO9hNKmCuyK13k/Fm1gpIhKD
ndBk3EjZBnwMkc8I/uB4bwxiFGEGCb3mlaBGpOe36g+ueGBTcC6LHDievNPRCQUz7RJfssLk+ACn
sfsWHwSDjnv6INFMVhxDxNix7j70TqS4i18zTuyOi8Rd6PZc2Az75Fqr8q2lD8dv2rEf3kc15sLu
Btmkzmbk9IxQMacIEfAP9ytlZcChhcFwxctteezNP/G98yNUFnJgMDikqRgIcnqTR2lBIk3fi1sO
1p5KTA0u1aONlMG86PznoSdwr2HABgdayX8kUgk0bAJRn/O+mDqqoPDJMZZeEetobZaFW8XU08hC
C3H/G9wS9Mf4gA21GDaboBv+adZK77F24yq25so2iVVPQMfCi/Z6t1YPOVi1j6H7bxQx8RehLIW6
aboO2johneZQYFKQ01PR1VQNvEHHiA7d5DKmWKOwQLgkWRCtqvAHaBZLvU7x0HwEIZY7KocN5O7p
6jRBFuq03kZ4jVDKx22128mqXSaArL9oo3TO/byU5i39e5NCGaIVobXTioCteE27SnHZQ/B0RRwD
eX4915ogIXVS77ud6L9mhLL/hTpXsdZWBiYm93pqIbC7Y6lpH50vIwSoLngW3TyRlXTwf6cBxDsE
9cxxwFjsVhe/h8wb4954MNOMEsgrbJRMLSwsxd1SP1kkuhB3Ds3g+pANZFG8KzGpnw/wwYY/sqnb
cpiyO/YqFgH1e3STUh9btrLBbsAwQNujZCwB0mkDgve/40l6wAOpCgv7tjOvIHPT6IBIiXWNzr4s
475u3+1jazEEQBsP2E4SzJxcp6JC1PpeyITEB6E3UIb6rpscWnhdaFIlsbNuoxz0ZK+Zpi/K1bY6
JqUBW0pUporFu/IZ8B9jd9N4NhNnU3EC90oznmRIpY5qXdcPMErOtUL+espqiio1JAWG4Vcl/vv9
Jf2ZdleN/Mu+n0ve78VJidMqYaSnpSSkQVMjYWQD2lpEUOLZozrf/bjkA5vFliQ4tFGGIhEGwhh1
UzKqxQNne0QIRrlc9W229JfOHGJ6ULKbQ4qN8tCyTF+5RClTTU+rIlYp9RnZJOx1i2qPTZSelIGm
0P0ycFsXO1TzOoA7/W8MWh2RN6TxCuzO7aiSzuY0qDMuYkuX8H/+83wclxYyDCw/0Bk2VqhiOWjE
0K43MQaG/RJdcWAs1DDhgwpZVDpSDZncUFqe6Jo8UrT4PtwPimh35xKnEGzRpLLISvHx3BJHkCrd
LcSN9BadZ8UNE1gAixlBK9pDkZZLRp3xFwO7kPcc0q4KNoVm6zps67mgrwPI56P6I6NW3vJx6Rni
VI8G+cFGgz6dA0NgHEu/7OveMdosstw81J0b4hZMB6QieUljkc5D6geETQZujWw6sahOZfOPh+Z9
UfszCBNoBOPC3opAemFxOoRoVxc8tdAn+jWn/Ywesdr4ncslaaTqKu1WSaHX+i7FXyOaqBVZhd4z
a/WusIenYu4LdA0c4qbXHIqFFktOthu0kcj66GQzdyRjtfeavUddUJ9qaFiD/nwGvbmNLQ6QIFrz
VW4KD8Q5fv8BDqdog/JB9emnUdt2GaoJxp4r9eLuvTbnevsklbf86X3tag0On55/slhq6MwveV9D
yzSTd4+PwgZ2lyLpSREzmxzIPPdvkvWShmLfhItGSQw/CKxlhwicZREwqSy8bczCKVvgjlkQi+Ow
eu7fn47O282k/hFuJTCXt9T+OE+WbccwmY3V/IvQVSqvrjQbvltR3GBIQdZW8rkF7+LoYlBY6K4e
r3jly0J45ab2SZQIXsYBCsMfO87/FwXvUnJoDSn1r0VPmXEj4gDz+hQwnBz/7zkOZX3F4E+eReO6
loTNN012+Kr5Yj2I2NZ3PrHlOGX60MUU95NkKBDBGwoPJpvlrk9u2y94grE4KDNBF4caRBQZFwZh
X5/+pvD7y9hmo0LZsFascrC8QNOp8NOb3AXuaeE0uBNRWoxkez8jOQ6anD+IKgbKVG9NyozlYb2E
sXobReLje5nK2BmWbLgPauxxTbByYZ4UPnG/PZjYc2CU4vY9QqzuNo/HvpNiLyUvONpK3qs2CdwL
yWvwaGDhCgQXHK93v+RDWi5H9DaMxR19/o4PBRIoifPhNl89V3zn3AsY1XvITXteSX2LBOx0i1SA
CsKVGGSjwGUIwP9fIHrJYO+55iInTCdxsy3qLs6/iGJC89ThAUA8AzpV6t65w/f822o0odEfT1ZN
koXBdMWkXM2cdcLEx9OYHksmcvOkwo0mMLfXaV+854FkWKW9KAUYmDcxMIMBfr1qFLqJeMo1YyCy
RKfBf6Ti4ckcJL3+VYr3NUVSHiq/mCisNvqUsxIpXHLDiWdN2CrOhHDHQU1ITrhMa2iA/1giL/Bb
ddgfGha6bHpRm75BKlsgzEA8NoQwIqmz4bfr1N9JMXbFQTHiqonvIPRNZATTyHwGvhHRiB54QB82
Q3MsmOyasizg/J+y6knVOIEWYGO0VesT+J7cqTIPm7vhW42xwvjmYbmqhi1Ppp82kzC62+cMhRDB
ZR/uvDeoACu0EnNnuLc80qFl0r9mWLqSjGEpZFKil4G1A0A4r0VgO18nINMnzBysaV35h5WNmtwc
hTtYs0qz6vFAEnGYzULxuk/xv6CCQ2UVeWjNFKv2MWzR0LTE0NDmSyUqB9Oa2uE5XdlgDumyNQ5u
0lx0CuFgMbsU3FMToBndRfYf2TOywhfiMGt3bHi/pdq81Hv9Hpu8Gsrrpg1Ng9JzZJ5KZr5dEF28
oLHLZ9YoZ36QxSjrvZTSvfIooRAeTCBvkpDgQGknWBdvkYMW49EAV9YC6mSRTxukymamYGHA6Le4
x+3pLz+6oGBY6nAgGYbvKRb1dsqo57ty+3cYgIEQQbhtSrscYpyk/crj+rqq7bTPPHi68p4MbCpn
wDRNd42i3l4F89QQOV+tUOEorBRmrKPMwKiGl+VQcETi8UfOxQxxqE2+Gjq2YZTSCOWRHvpvNbpQ
+cx8/YIwlIO6I0KZR/PvfcTvdCDyu7kV5Yp0lIGQMTPisxz61VWbEotp92q9UJ8BzmCrLz6KqiV8
pTGrvTxpls18soJWQnh5agYktrpfXtnNYweR+s5tW/DB5/tOvJb18uziWk6XR8pyi/+cCtdsY/ia
OUYMD6i4TAvRWqtjUD9pJwSyc1zX6opQvitnRmhjjLWsSDqBxwvZi5wXDNeZL1JGFn+cO/vsf701
lk0E4I1PV2L8fxE1l0fUU7rjtDyrEl90Ff+n46ahhkoK0oD0Gfw9kg9ihMVvVbhb0Sg+GD+GxEIb
AyWRESizjl4QWKwGkE8WHhAzonEeKbjs91276TedbXeTqlmFBc02hSfr/9ogD4Ngnu7H0V+HDd5w
mD18a3WNcHdcDBL/iMY++q/ueXIt4YMtghVexdZP7Nm3pxi5WjcVQ5PLM93opHkZm8EersOEutFo
ejRr4t1O3sbmsebUbEiigld8enb1zA/TgB+VXL6cxz8poBZOEMzenTJubmNOYKnD4Qrq0ns1Zqin
am86SV+gGW6KqaAo81YjS3UGKq6pbSynIEv4JnLWg1cswElOSPPIciQqA2MOTDglP9Pw3b1m4isJ
+wVsV6VNDauir4EQNbAURTFBiXX1YRkHFRnEwICq26YVcvimw6tLRki/1FxZh2YEhggiNUvZc2fZ
eusO3SRq/SPryDT0K742nOCIg7BzDQizLuntQomfmRDFggx10WKrWia8jiCezxGKCE8PEfJF1lnN
JtpWnOqDLWUQhTNQsq/MYjEdejaASp1XtDCuyGwXoEbzTgJo7tY4qQeoWw1D4CVDlRw5S8iFcjwH
Wbo3NwIRmID+k5OwV8/MqDLP46/0blnf/sn5fsDI2e1DicGSvlnQVlpiOkXh7yyXBvygaMGJRMVw
Qt54byXF+zHHo7W7RNGZrAT5Jk60OTFAe0k+OoxeG6oxSYyhmjL/V+tbnG+hmPD6L32o95b9uRN3
TlEL6B8OibZ7ur5xzXZ2lxq+0qFY4lSEJX9DE49pM91fNcBB1cv/PATSx6PbsDahgmgmqNDtMCcg
lB7lwJGNDI31BKkGLOW7+M3y2ouExvtskKoLGKNBuFE8h0LgwCWB0dyBArTNMB8Wp6qj5uPja/Ee
itu0XwFhNsjRvN2SjBFl6e6s5n+xSjeFjiuNA0PuO5qqpwizaj+6vEAgbHiX5582Aqo/by0kk+GI
tyArvTuGl0iZhsGNBrGehVgcdgXXybcEfbo4rUEGX+pAjyv6Sb+VQIH19PG5fDx2m5j0nyvWqFea
AHfummgI1+gAo1HBkJuIECa5+JH9Rtukly8uen35gO133vJLN7UbmtQkMYAmYToDIrvVhH/lR5yV
4YyjiyXlLKHIfRSSnUFPPIOa7c0DpCnQUU/D0rtlk/bnbJxBhXO5eZD0w8dT9bxK288EFeIxSfnk
zAR+iGQd/FcQecHO31skbXHuaLFd111S+N+WQWodDBiLkZljowrXyXzG3BHo20bct1ypiNBmV4um
2C1e4UeueJDFiNAybfwvOUhwfBc3C+gVYJSH7WSg4bSDB6/A3r+QcBNtrFS5LiwzshL5mTsfXYB8
sVdeLKffrQ6ms/kk4PPwL8ZYEGU6unUfr2BtX0yXBzX5s8BEjMwsfKzGJQCIUC9eOS92QjreMMo6
DuWSkf41a4KHl84I+G+N9DQ2p4dx+WX2bZ7+xKt/98/j9LZXwmdbZ/FzuEk1wiD5mAeF/9BrwUhn
OZV9Wh/S8/5c/oNFSKSshTZC1QKC/cIRykt4I2zZEBTk077LkxQlBIBX+I5Kis7vutQrz12Ta/CD
pq6RpPtu10toCEczDwIA3UKK8NlNmazJ6H2q4FSuGSKpAGLws3DCWg4JWn45jNGWNcKgDk58CeVP
kVeHHg2QM2WG1DIQzAJpxvRI4PX2buCZ3syKs6XwOwL0sAhoD8jJWgDqXCuqN3NaYYL3MXB3rlsk
K2cMLOKaJv2DQIw4/4uA911BAB3y3Po4HkaCX0EcZ5ZuupKkfjDdmojArGbotdewq7ctjj4EBSyW
ZVKBwz/ssABGehDdjY68GDd2P3fG5ppDpuwl7hYlwztgejshCkodticxRY2xMY+grLUhdAlnyUHB
O3AQJ6FaSsASXr96LGoiJ+YTlsVu5R7bivElbzanag7NyVcDmaZk0W60BTCW+up55Aqt1FKbDjAg
nM5Mq54I7vRAgI94bagVIcMvm/TwinWS0ZiOJWZKzeMw1yyKaVeedBcM6jWKG1Fx+NLMSq52wkVd
a42u+dl/r9llP86H6rP10wZltepbbkml05SmnTrxFAD8Ya/fN262UJ2A2NOf0T70z2FrkoKvaJj2
7Tl12ATNuqUKNwC+itGkkRVZxdEj/kurZhNuBxOP3wc0WVqwFyyK0F64Ckk5Fa1Rq0RrV1BEuSwy
N2Guph0lFNhahGN+JephNWzCwFUdXtWCA+2D5whcKkwOKRwN6uhLZJHok5T0YNFExKxRkOu8HKJ+
6lVzD5iZN0i7t6iGUUcawWa2aD8hCnCFQtmWNXq7KDg1kc8MbpKmAhAimkGEVhhZ1laFAH28DGW2
44eduxqwOLTkLWkNqeZMMjBFpw429m6/2NpQ7U3WndQsWrNSFDyqVF6tJ03phsbmrHhCBbPLC41G
y0TToJC5yOC+Z9jdrHmz8ypu95bmF/I/ljDrkTz9clvJazRiNj8INP3DPQHjOUfCASMaCJtRUVTi
L/mwE1W7avz5acDiNOoPt+Uh4QqBx67jnErvcFNx3RQkrKdDTNTRGO4boDnpV4Gt5SYuLVLU/l3e
ejSppUOmJg4tr3lX8jY0IQ9vUgWxJWDrEOaOLmF+1sOOuVz0XQTabb+yZ3GNjPeAyEQijJZaSG8P
5bPYBbMVO8tDDRjOrMTxokveuiVYEkRcJkqQ2XtVZQ4x/TO2fCAFL1aLkYk4KCjvp8pBvecGsjBX
3N6fw0CZWbQhYcWK3INaXuAyONrBqa1djHhHeMDgwRCuLVJf3eEE/6pJW+++Dc8AuJAEANgpMest
rIMYUMnPnQPrvNafDv4HzCCZ9SgMhdaPHFo2/GSdhp1UMUXZG0mTRikW9Y9fhUinHMqxDpoK9JsY
Cf1mhoIels1skABHx4ey57G+5Nk1A/XAtqarnBaoZrP5Nok1cRqz1EarraxE4dk07R4kqBwLaqur
FNVdlN79D1oO1IJ1fG7WOzKt90KEGyoy97K2TwjHt4bsT3uRhqqVE2GCuSszmePcseP7ESdMNt4g
fHUaUPlqAI21Dq0cGpLOhPpvBj1+lSG4nySooCtgL7dkKzAHT0HSneN5TjcpeZNb5V5CZKPuzt7r
QzZR9Tqh2NPi8/okqNdR/HfYMTAKzKgH9G3WkJ1RqdEZonH0jW54z8X5T/qyqqL+4lW33GQgH7ll
gRZwFPGefM7gpcdeq6NPtudCoC0ZSQalLEGFxeHvkUOImX1iOHYJpFqng/fBpcunlSFuvUV0v8UN
8xSmUkDxVBVTsRi8D3OCKo6ThQz1H/B6pmYZzcsthilQT7UwZdRTlXZFjSXHgmJivtm66/j7bYxD
WgpDUfi6uU2kRgIX9y2kQ0nECKKGTGGlDzk1RRoX9Faqx4Qc0haS5IbfvhmmAWVJh99vhE1fGMHD
5Pv/1aFk8HppQLwGCIUJua3Udf27j6VfS3tXywxElM5aMWkQI/msenYvgV/1MtI88X60OQ0IKGRN
fwC1JNC20UZAeJBOw0qBAP7vmE/9FnpVyW9PNZX166ZOkEyFaDb+Ig9JnZKj3AUoVZxePn7/9GOw
J4fRcbH5O7yQYcOLHNv5+FBRERx2rD9QfeYL0ywcoALXeGMOSUd7Pkj6b/Kj0oJAMTu38UkitU+2
4AV6Q12N5rexZyRbL28SrEcY9XOQILMaQiDJmro8sAp9zq6lmvw3rl8Ph9a5syAFIiNIJBFTpLx9
h5E+4XToB/cDHvGItzGXQHmpTS/ohW6QZuw6KZgEkaD7fY+lynlRe26w8dFzyb/IBT+ULCOoFqvR
GouWrGmPYq/+tkIyRyigLPMYqpKH/VGTjWsguF1Lw9CgwG9khIQkw6NfAB3m+gSrM5Di+N4IosgJ
0GMw8IBsCWSSsNU3/NKc0NxyGJIoZ8LozRtuKzsh+CK6RdE81GahBn8IHFNMUwfZw5cbIufeDUt+
aZsU1L4C0sazkIw2PKepLcOecXjDQA9nQOEgNxgBwDFfMGJTFoj0kUGN3DIuGNDUD1SUNI3Zwb0L
vkKdUMMmWfO3UgmJPh0umxQ2JIH0kZbfvlDjvkGXCpocZM1bm9bg2PpcjkQCnpNqbrmeoCRqk9sw
lb+4Dowx4W9KsPIA8qsvRHbqeEtvz6dnH+fUIDOpjqESzH2CNjqxmpm3NpeH4s6jWaLH5J0CeqZS
8YrMIKOZptDbXK9c+OrICXXZJ81pzKjzLG+2Wr+VsskOMCuLG+5K0aTZjnCfIDEjb8/2d9rDv7+b
uO0rwgbmfBLxkOQwNnGTslnIx96Xdoo7iWN6kqWP876iPcU1B8Ofi+dWVjXWflTaRfuLFugR9xWI
WcYcegRWDfEotjkfnvmeD/bYY3LwVs4Sv+0jIUFTZvXibZFNKIpSP5Bp+9atYphTHYTMSeG+MDkr
6fPHYMDD/TE3kpLsp9PiLoQLLKgJB+9YOY22aLaEhE/CxQrk7fQ0NZ3mxXwAOFYkATEGsCkaVng0
oU85qnnXCGBJFBc2A2zeuD+Y2ghIHb2vE7IiYDegwqU7kh8zDb5YMutUn+iL6L9yugch7HVEWi7z
fXALukaYSDug/9GdqZ5L+Z0YPtIdmhlvYsocH2wxLFdK8sCh05NGk53unfaiwq1p3LjsRPEYyfwZ
tNqGv3N2ofW/Ep8TMGux5Gl1gWebASAWiqPw8xAK1AianRixw0ps6Co0vfxii9nIQrCECyZTx+Td
rz/AtKELgP4+FYDGsGHdZs3WaeSLwPWakP8TtcQrHA1jI916DvD1BcidYnVTEU09CySjgMSvEjIG
BpIEqkw1HHb/G4EjJrLx1Qz+6e+8YUq/LaAGxtToEhRcf73kgcFV7qlOplUyop2PH+xPzDvIeDiA
yKSoWmLL1ccYC0uqcUNGppvR8sIjrer8tcNgGw1tXPP4NQ3ro7X93bMp2e2Chy/mtWANVAyuICtM
ELmzXE0r6vd46dmSmuK1uq0Yg6QKuK7NJ/V6um4NyTJ2zZZoEef1lCZbvuWWXiSKm7A3D0U9EmNj
kjeOoCshvrtwEhLZlmGjnqBL1/mjhPar5wYIkScYZCetpk12pO1eKeLHmF/rkL2ArgCOq8fvc4R/
2gzfkPWlknUGZqwu+vSacCJVVi4UPLRY/PpnbF6ZgXHA8btPBJnVx4y1wt52HUQcpzC8ME88lbEh
GF8WOVEUnCE4OpMeCI2yT4+mzUFcauNAY18+Vk9Wn/TWM7Pt2zSpdcMzAQXDH3oddQQ9pnWN2l4V
l2E/AsKfJ0h8r2qBx8ZVospXQ0L5vNsublFfpjp6dx2m9ofvj7yvk3iZRt+8WT9UOGJ7afyQalXA
eQAniguFKh1Akyt0RfXVJkC9AqHaHELMLWZIQoZ60Hi3c0I9m90V+l531ATE8oxt05+9wGIJDyo3
ZoJDXzO+ldTxWGCE26lPBi+JaxxXhticlUF/dwvF02XNFWdkQTiEel7IkAHaMyT09MuWWkSFzKhk
aC8R/+fzXmhM7Xtssw3ZjXJC8CGNfSmIhhkTPOQGe5kzbx1arbJIays+hZXpu8udADafLZGWBC3m
zXxSY+LJJvYx29zQp6EO3kzucknpp5x0yIk1cLpc9sFBJKooHjDX9911WpnhdOS4pHO0TnZbKIb+
/s5593t9lPVLvokkHZ/mIHLAx2km/6a3IpHhdmXmCAhwivDwCRrwwwvm6geGj0CNt5CkklIp32ET
vfKbg5E5TBix3krG7gW4LgzXLO5+YozbmMEyS35koectpDgriscqkj1AyHIIr8QABrArettYmptS
Afn9TPXCd2lqMrJib2zuk101KlFTawIAa4xp9HUIPFUINPL4LkeNHHTHfbUJBEH7rQrg0Rxpfv0X
iAXgSIu+TZmrXvLu16o9xDOwyoMZ/EnBZk5PKzYmhZA0mI8128iXp499fw/wDGc0z8sqpQtTLhRY
dWymlpnL1IH1Z3QZyZleHa8h/gaGsJ8EsZWOTs68OiNoEAezYJGxrJOUDhDs9OvBxaSPJy0gmYFh
R5/Rz8y39tnbGbkqs/eiaUFmdEgzBRclhDpQfdo7j7R8ZbxdCigx4SL7j4S2yczTWSPhXoZHxSiB
YkaiWrOYvG3PUmB8jA2Z2NoPMosW9D8Iq8NiVqtUP6MGyMY4ezYWHM1BEiM5gYrP0SFyVQbapvgO
2a/soSdEGNPD2APUrqfZpmkBfglpUfjFGsBLr3Hv8YtqpuFoDPGKZbYWTG7B3NqAUy6NlS+IAeh1
pql6mj+zBbUF2lBTVK7SdYOpQ3n7yCwLarYmruriQN7QG5JR2IHam/et8E9sLxRCia+SCtpLgjxG
bFL0H/11QBcJ4SA61sWiCnvmhnEv0GkijjfyAqmXqh7/sPdKON7s5/HwBjuBcueTra41mmWWAO+I
qK5CNWzWNUt4BM4dyJUTcxuEYyM02025GjqOu2+jGJKZFx8TbKHVZl+O4Y1fj5Uuz7uphJ4prm7R
xO75lHDqp3PFsC5QtyEjWB5xHD6mLsmTKT0xa0SaGDLc3ZonPu3OjH0N7tkS1TG5fzloOKIhGWUu
1QJqd5QhUvggutSuc4uMp6PeSyJZIzYFABUtqbJVWw0zZbt87GM/mro1evg0aTHOv+L7wp/xhknF
Ti9/h9qNwaRqqIRT+xLvgaJPxxtOBfwu0/AC50BXa+i7c4N/VvKDP9zXU+CmO1qAL21fHIdM1ik4
vNFZwFDIWSxXtTt51gpIhy5Mf5CSAfx/awoDIp1JjoBJiPjANS9VPZ3VrRY/hczf6CZhc0PbPkxH
zLH32ECMJxpckOPZy/abrhtWRDW4FqJpwCHWUMXEtma7DtKdl4pzF5726Sfy/7sGIwCVQwvVoVhf
Yd9MZBQom9iliJNzI9womsOJb2fLnFBMxcv96np5soVHmW+jK65yOtA1QIw6Vk1qIt3N+ZMmnwRX
QNQUE7uldu0DWexPxleCXjYUt+rRBfRf3lJqaRvMDHywKESeTc6jDtRqP1cL0R5XbbRqlWBOLA+q
uw4p8eGpunUTr6gtk42b4YwezzXkzcsHNgB8HHbkbICyo1Wiv614kpPDltGCX7Q4aPYcCrp4YvHU
FgIksLqGdNgiaSzRozVnne3GOuXepuX5fwhm5DtEdsexRwvqPODPE/H8islEgPkLprkQRG8P2mL5
3ksSE+YPwW+Nv6SZ0KS6xkxWAAPKyeecU0BqOV3HTvo8GP80y2PdvadfXSHpfI9UZuZN+oZY9VCX
3k3kYFdJ16ZptaTTXMptJ77dMXQl7ltM3eVKzev7ROYdC4ICWtpRnNw8InzMeHL0eKlaYRc3RCoN
tt3Qu9VvnKUlezyfIjhajGUG1cTEs+0SGTYjyl3K3y7jGBSP33LPE54Obu0CaHrXMtXSswoV3dIs
Z/FVu3U20/8oZcQCIoq1QBnE4CyL7Xg0biPzrFN/0FFSS6O8zv6zjjgN0Hk63cStzVekIOxNh81A
KS05wLqW+RYImYYPgHCB3nDcXRC2+9BBYHpK6vwObztsQLN/+fGdv5vHzneHoE8LdgB0ic6LQqkb
SNtWZUnLzbQOvhZCA/uGnB05CqMpEjhbyl0c6WjrwXHovNNjSg86EBvvY9jniQgqZ255nXRRObTv
TIadQzlgxdOl39KfijgIMnk0n0tqE2UCll0d//k3pIblxFwpsZK0VKnV9v/HN074S1rgPz/63kP6
/WzE2fT49+P25Otj7TwTW0mJp99GzIKr4cdjSCT7JzMLv7P6LV4S7RTifeFSEFBVaBcQS94lWiid
eBsc0srHrxtVEq/cO2J1j2+394ofzuRmGlZQcskicgLrlg4/jsJrpsSxI/pv6hFi9ZUAURdW1lub
GfEdj1lEwmdpmJJkNa8kcG7+b0dpJIE6EuPBKHK2TL1iKHMfdJ/Q3yXW5TFsVfTzJ0ldP76GgYgq
eKwdL7nDSGEEgBE8cd9zKTK6cXEzQGOSanBEZKob+7qCF8HTU96GiKT7h6Ez8IKKWEY7vTOX/t6t
/lvYs8duIP9EqP4rppb8pEd2GQFVQj5YscpjveSsFumABYzQxex4ej1Ka8Ts7cKNfpFkaaLAbTEE
woB4YJef6OfU7+aOLcJ5rbWe1Z2R7g9XpZJntLdRUYY0iskEvqbMY4WsjItSFpvgMi1vegOZbZkG
M2ikPOBCzRbnGut5nR5H4ViRvphEOa+aTmKypTQRlnLzcttJoUV1F3HSGzYih/bQCfsUv+Ob1kG2
SsY7mCWqkN3xagin1MJWq8UG7VRVodUfde5sLFeaX4F3DsxLVEM4zh6UXseCGzB6LCAJ/ppLnJfX
L72g1u4mw61SuZHlIjQfXlNYyxG6gZMnPCfLa0YKY+XR83NbHxvHbUyLS53/ARJ6MAZiQ48/UaGi
GJpS2WF6yDSW/03SgQCZIE1kienYGynEQ7R7csqb0aZPdzT80xJw0r1YFlt5qNW8Tzx+3mwni09a
pd21Xcak9AzmROXzsUPhctFeja+rtFy2tV5iupneToWAegMDBXaXjGDpq3yKi4ydZ6mAigNgprYH
8X4MTdDuNszQgfrKRyQL3ySB3wO5DVQlf3bvbeBWgU5SGtHPHi2Vw09f80QAnLnuhDjkFnFKZqKD
BJhU/uhTwAW8TiNPXTXprpqQ1odUYjFW76NjmO1v3KRPhR2fyjyxV/4BogahiY+gFIG2h0gEOlVb
498IKiVCGlYk5bAiumdujG23OXbK/t2RRmo7KN/bLNGQH+Q/vV5cKqH8DWrS69LuoyyXRd7G4M9+
Sh2n8wC14C2PtXgpBJDxd7fbB7lYNIfJCPJ23pwAybIy5GdzmNkZzW5qg9IRWhCNM2T652A66uLs
b0vB67u3g6pDjjk2CqGU3P/rQSeMMdn2fJQLzte7zLPyOltSOay7s+rYz4Nc5ds6W7aE+m1Zwk5k
YCb87wRHHXRQyNeBj+s96ya9LGoBArhcrkv9Wk9uQMTds3BmJpjmduDdc6ZS4lGtvmymFBEqiJBS
qDoyOcxFVLPxj2V6Vd1v9uU1/pYsewgwKKnBRju7Y0/Re07eyXMk/3LIeKIFVP6VnKd/wDNeAPZt
+rWzUFbWtgQ2BcX/alXpEpbIIpn9Q/SQbLsvZ9qqtRlOFoSJvWd6wpDhv5rMfGU4K1f3jLdA5kjQ
ZvKnVkJjHWt8WZ4CGQV3wqPuM0QeoP4xQsPWrCFAyPGDKVxIdyX5hpCevzy+xHRX+fSVvPHCoUkp
ozgKB/t5ufe8uSUrhJAV1qbebEQ0wjcx2bzmEmUlZyKobm5jqYUlOp7BNRgpW8eEl1JouVJ5MS38
jEbpXuZhSEBYLeHsnskSySwwiALD0ZVLUYSJsx3NJtLabLHuq/sYAhKPfkgycgPKXrdj94AVh4hK
nnPtfja0wUOW3evRcjv9puyAKS9UmTBrN0SXNKE8wf5ZPaVb3SudHBLAKKneRbLj41uzqcbfHqJB
8WjFe4+RiX6vQzrjbg4/JGPSm2FGffQ9vCvYR1wcQy1jpnjdbQo+m2UOKmCH66LRwhsd1pE4DN54
z327YjsQUK76vVYIGVcKLe2mJlfGUppOhc5t69wB0vPCVWUOG23EkdK9FzInY4fM0PxhGzdOTVk7
F1ggil8E2nZXqkni0/0U8+a0Rqt7J9f3bI/W28Gc1OKYEndFz+wa6bTR3JgbG28i5rzcAn2awBBq
uWO7L7Z+bvpd36ZgRYz8xnYX9k6q+CUrVtyY+1TSzFcj2bOtvZVXEKQIJau9fGB4RCnU/6K+L4GQ
O4dJlVLNHlcj4GI/vhJtjmdNHjnekL0zKidgzZ5lAWh8hQ4/t2Aocb3n5Eft200bmaEvgpiRywOS
oFFDSt5dZoMWIB1hzcEL/5a6yGgaUKizERYmhj8FutRzPeqAjxnqgABC2eZeunyRL7afxyt4jVj6
iG7JJEaNfmysYa3jYqDXM18g43vQCxZYpvyYpnVihpYOmlADmk8lCfscZUJo7li6fmN4IUWkKm45
rgrqxiOpMtv/kLe3aRkkd1HLW/eO7kDg6XgEXSxRJYg+vDOYWfJXtbo35ye2tZOcJtdeYsUrtGTz
h0J4H8y/DHkduAal8P534+gTPcgY6RUZkgsL10EdMghe2JjF5kw5okiq9goQuWgmxCzUQ9Pw3ApQ
cP15sjQxo4hFF3MtgfzNaWPyuH/u6mPHOafMQiYLKrti8kK7SFdFDmKEEyZLjpVACzJYK+Fn1PgG
dOomHVDk3np02JlmblFC7b5IuXR/rSM1Z+ZSu9ZSXHCs8rGuKH5xGOf2hwX1HbitMSujDui8t1o2
9dNNrndBzflrYrlWpKuUYpFmbGlwbOTLe88HQ9gfYXWrhcAUJMp3U8JX9BwA5YoKjEudoN7fIqWF
y7kcgEWHhzVIeqegCRCc5zHzd9F3ZaKsGCPB8U41xpEu1D4WNolaF3bhFxD15jU5Lw7dU9lM6Fmi
I2fg6nS+bVt7FFTUY4R2L38ZcBNuMwPHujM69SC/eb3FVk1nPOAAd/1Pl0ULHLrSi4u3WB36Dghe
NSHuAz87R8343n/ezp1tTF+wCkanfBaEZVRGOGBGcRO8G3RtohUOUmIVrtoNlLDCTATT/w/osTjS
19Wxa/a+R0dC3qdacTGPwyeg9cusT1Al1rfOchg8jEUmfG7g4tw4idNK2F0emXs2LqgcMUN7k0Up
5fq34v+M2qRCnEUCdzvQv4FILJpzSozOd6HzDYk3hsaC+j6F/N3uAscSwi24gfYV8igt1ZOtn17F
r1QmH50CPo2l6oipsqbd27JVw4wcu1WroNugVyw/rfO4y8Gl1dSRctAJb/ybP60hUXTvc5EBe99j
GY3zsgjmh59Q4mDEnD/qnVI2n+DhPVXQrFKvr+EvizNvztFOFpXtfXQtQHljjiN7TTGltiuez9yx
8trAcdGsSoEpV+08kVDpUHEn4Ol+aeVYxxu4pYSUSMfGiNoFQytNhCDjEHd7ieicCDZjH8xf0K25
RdNaNnCbABxBzOPhO8BF31W6UtR+d0zbFedsO6EMhCvqpdKEm21x3Izdpfg83eukOL6r8ffuUVlh
ta4F1EwL9VWg4Mcif9IbVXZgfqP02kPhRrT81NnDH6txTdpiI9PPRHW6EH+jfNhVXc4WIkLeArn7
6FtcRrM9xRue+YxUmfgyTYRcvmHt9Dz9RXSMnBTx5V+3FKrlLNgrFoTUiqHur+wgvglXUpJZm9sm
qngq27e2v+4FU67BlNjKGbwQiHUufZhmaB2nCR8p6eCalUxlrGs6/Y/sdYACTmVZpumrcpbRgXsd
sTXecj/LqoUy6Y+PhAIWlW0qWLk85vIpLwiZcHTHzpY3xSXaybqpTxb+IDm4JIyfNucwY94lYblN
OqYjt8xoatIO/JMu3KlI8TxmAZWZjCM1YEUvB/HDwf5giVwULgH2bOslLDo5m/LkHdzRMYY9VnTq
QBOYmMIZZGMqsWIvCIKdtAh23zBhiNWL9l2tk7gSmSH9JKgHYoMX2JECAHFjiK/tWzsVHbD2Bpjt
JggYWaevGpthurMXQFh9VxT4hhtVBtagK/jALwwGvP1t/MJ4VwRlHu8sMJc1XGLznDiw7S89xYzC
8j7EdDOH31Fkpxh5GyKaePiVRJ6NWYacj+e3kmHlweM60O9Zu5D5zY9HvkDJ8J8Lm3coapmnMD3F
dNfM1zkhcnZuxAfNzibOuvoHAy4RouY4LIaCWufjJQGyIQ7HujZNj5Y+pUAsVPT3oNMpz3vfo7Fo
vQhVQyojcHz+RbnQlgfGVwNFiquxzYZx8einj/mOjTXAZ4mZaIYWdGEtsgnz+mLRebkgtdhi+9az
6wyUbEakDolh9FUfRThL+k2fFLXF/tRem/L5t/h6pnbSy7jiLLZI3qIa4dR1RYhcsasZ2WDIAuBU
0kC36BdqUAqcTjbJSOfoka5z9fxMz1FZv0tCsaDEOpAU56mBQ5Qg7UaGiOQJB0WJP3f+DrXfNHYO
Q0OV9v+wGCNqlu6SDqwXFDtECvjSmlUJwyS5JVj3UOTpyOwLTFUxP+wTDYMwgMb8yMTWagxcW46C
XHu/hsp0wCHSMQ7DNeR8ewon5FtNYNknUROGjDG5abSGlchyb5KaEYT8yFB4irCLdSBCFtPa/T8A
OmWvjYWSWhfR3NxMPb/Thxx+Dl3eBLkgWD6vR6cfFC6EP/QtVe/Wlhrpaa4h95lWXI5zRgszaIar
MYUldddZWRU44MJCfqJX1vRZ5dV+aSqvmVThbynQfmqZV/WkG4FdSKZizSt5sGsKk0fc+o+FD7I5
6XoHDlKCC34jvM5eaoHbbGUEiYliA9q2m8nrVESt5XdUpkNWi8V/RovQA9ENXgnWdQAUI5nOQ2+9
SHeBCR8BzawbUYPkazbYlRsWBPXblOG5qylaUhSycLlTeYV2fqRronMxm5KMh/MqITKi+VN8sKLY
OPsCUceee55IaOSLDUOYTNZbKDdURyKPsABqlWPvBCVpOPE3UvZgcL4YCjVtjCFtQvaUyhLy+VF+
Ab3KNsMrIDzFSNJm3EvxOY0PuO3oXsM8ZCkH3frqrnaaksz7NMbcube3vJDl4qjhaxAat/xgAbL6
vj46E6C/ekGD0FC3eRYDlQt1A8tMFxt2PAk7S1Ef+VtYnPPfI9g0dvD3xmbx2NPVdf1fGGPZYoWs
WAkhayp/jfJwE9Z5xswL7BY4AcRDcj38bd4T1OKkbgsbDg7H2vGwL2+duV1boYqreKyN73DK/pd/
iS4pqIBByOcvn1EPrg8ns5LL9MnL4sUxkHW/G6plblOVBqd+FzMDNs6non9QBHVa/shmsVMoJvz2
++ofqhCuR8WLmgNg4WQwh88e7+k/muZsXZChKo9OVKm0dJpVe8sYbe1xCOihWy+pP3OFIwa/grbk
a62xDAOtuk6h9DARbQ4xixWXe5TvndWrso4aYljhixhZuM8fD95uE8HUONOZknDaPYXjLxijg+dh
JhB5fCIXRUz4MDvbFXjJgvKvU+VOa/3Vv3B/xJGcW9WfQ1CqDoKQw4hKqPOMr9hNGn6/FDj/CAK5
nnmECdUNgZ5rZej/UCb2aMze4sxc/OB2M8lePJ2wa5aztYANrd0Xt14+vpMnewl+XrffHYjafZG+
JMV0N/Y7BSPecMnpbUd5P62b4Ut+V4ryaF51lMfBxpWWb5Ubcm2qimwux192DZsfTM1cAN39Efyk
wNbCKcZTvia/i/jL6+K7ig2SFJldSaq6NamK7GzhIbiWDJoThSNbz1RfYfdmLiBcJzK/QJy+UGSi
cvyrkMGhEveZ4vaKnZeaEFp2pDOPRubfEP/6WSqHYV8BsJ10EF1pbxyf4yuzNKxGWHwis1MObb+4
aM6rkY1zBG2z9AOQBjPdHSBXHobPUWVLPBmzeDseBIO1zcgtOXSlB0bYZplHSb7Vi/jJ+MBJA+ga
cVk6AIILapYPQ/7u6T6ULkVXBo3W4Kgj9E+GbtFDEM7fczmDvUxGzUkg57Vs8NvOPzVRj3NQezfC
Lkpuo61qACY8UrPEswBu2CJNbH3jN4DgU6VfIaBlWVNqLC9JVeN/ybZJoCTvMiTnvmH6ZOpuwkhN
GHhoQcKErjHVJNcSEH+l7oRgWCXgpSS2xD7ROnR1wb42t+CFEkuHd4uXgG1/qTtCEava211lfNkt
9VG6ho8LSDga3kbmOuHuIJ7bawCCBof+Km1pkNwgEtzxZUJtHg10Ks0r/SqOSqOr0rD4x9EcpZG0
VysnW+867h8jyzLxNu6s+6CrBuB6zDAhGCeXVAIghM6wVsPtShJ1gxptZ2wHnLmSDckUchHk7PKp
6JwWvSrhA8y0nuezGVgHA1x4OLCF/IL6ksYTiiqjFUs0li+VCJRTRqhFzV75pubVcDrc6I6gIRCc
zd5VqtCZSk/cG9Lc3SU3ZewhneIS7GqJxuJgrvO9EmqILtNKBVkh4bDe2jVRvfcJnoU0oiwOk4O4
mb4X8EqZTfyVVnNWTsrwS8A/BonKPnc0t7idgj+HqnPniIvNcvnfhICdLpPXaKuVBzkPzmQhwooj
oA2CSQlFm6FJYEfZY+GA4s9+QLcyoegWhyImtosWA4AB/YFawOlvKsRwl6GHFGLrV3q9N4MjKTCd
XExWtByJLu0E5p3JOG0/680/uXADYr6iaHZC7ja4wbi6OVzVJDgVNPGp90u6USIRy27/kADwNPWU
sPT2fC8XFR+FII7xjFmY88LlVQ9fqAmQd7jYnIhBnShAVP2alLz8zVEDzjCIkvqoVk7/gdv4Qf7D
d1LGkniExcGYbxt1erCzuD78Y7i5HPH6vW1p3kChg/NLb0RDdc207kpadQy/DM8hJLGf2xUni/wZ
7N654gmOgao6p59FOGWH3EBlRTr1cpjU5DdTiz2YcNpD9LcLtRw0h+tdfknHg9PgmNgsaV3KYvPa
l+gmlMVZSt+GHuOCwsREt6TsrFGM0LKjWbUgeu8EU5HiYY6ug11c0QIsou7EEaoQE8NN7GIeqCVG
VGgxooxJaeTvzblZRIYPa2qNWvZ+8DtQRGi4XcokW01CeQY0gnAUrPpT12WY5pUe6pt6RC8qqd57
J4q90HAlJC/uYGAheNVs1O68XOZE3fiHbykjW7QSHvBQE3+6DKFPdi9L+BmfssfOwJnMhrtff4Yy
p5yv1GdMeaE5MzUQ4JhLjIxsnropNqvzkOESV7jW59CQmkSonzQ4JXc5Zd2uw4dQSwUmn7wJA+E/
JRI3g+STZN+ZCK68vjjoSP90eptS+5Y7XOvPRoN25StVQWom2BGDtk7SctUk8qoAQEzFx3lV4F+o
ocZ6lEnxtixqYYBfOvmUcjPOap+4vQsjx6G3uv6hHPA94ijbxvixk0/8xbNQrHptH0vEfZtlkoqe
Rrq6lRK3mVzjN+PpLyng4j4hP12tE+tKCGqTOIXRK62U+IGXMlKpYq4aQFSb8dkWHcApXH50upWv
ySGMc775kp0iQxMDZ9ook2PsUGz6CJlAYb4hEMNW6Bwm592lGmj2BpdA5eoqMJkzSA2mp4ryp5Px
txFtVye98PU42Q9rD85yyJdJswHUmFRPnK8nxTDqO2nto1n/qgJJvr4IcPCLhlDHga54RF+LhiRp
aU68k2lecColiRalKO2Un9m+x+dc/BUu5JL1AbbjbGW05r72IMODq9UFgXTEUZwQC4eiADdhxvQE
jO3LbuAYkdlivKs6dbu/8GFyFTnYEpcH7cFnaBM3UPMrtQL091EbtiIVLfwLLKHbIfVXtn95mawC
9VPGthKiGGMlIu+6Wt4PqIee5YnraV6Jmh9jBlC6HguSxlmQXZwI0g/nLjGcRbxh4ukj/28vgH4j
6kmNY4XUZT8o/vCKkGScLq26aIEn3nLkdIVwzX4qyBnye8v26RzuHwSHod4kIT6myw+WfE6LjAgU
0oN7kBI/YRbj1cy5JVKYQNSCNycYAzWyAvXCZnrEVT3+4KHCI2DswGonmo/j6vfNEwIdHhUn9x4a
P0RI9E/Us555Y8TZtqmKDQvOQptngwDRbo0r1CejJuVgOFqqBXtOLfOaGA/k2kjzXPRi5HmWyF5H
BD6xD9BxiGbuTUHak1p/w/bbRuBaIFcd8xC2cWVpD8kDjLa9tGxWO2t/MsOg5HbT9QovG2b1qlkV
kpE9AfjmB5tjIbtMRctxxXtHwkH0L3Rtg5Inl4MJDjWagdE5n+yp/eqQgwKkOWi3cLQi2pABdusf
gjryx7i50e5T1e3WACK0L68G+KEpkJfWZWrPmGFBdjOMM7t0KEcITXuPEl/JealpiN0KgMxtuRvB
CuUp6NRJERDifFKnILS4UBopcAQgzU5gYEYVLNkXPWs7tmIBRtWG5btyuQfoR8+t0mHvBIvAS70F
Kyfg8ABwkCwPNsc6sCH6XcUbaR5r53pLjfPgU1JJ9dLYOGewmFlN3QTHOjNSv1u53xFbw0uZnjpI
d20NgVuPdT0T1qcSbeUd3PrDePFMINnbw8KKpy4fJhSsDnsAIiJth9hlzBSLNJTs0Bkoi7Fn86RG
906CWWD1WCxgBgnbjNKAJizYvyLGOB8GYRXA6gxvguJa2hM2g+TKqW+hOohKYJbktGI5WU83XmBo
b+vbMd2aOP34BbfQe9hGFwELbhjYh/J1KR2cdi4g7aIaMV1BTRdcybe3gr4qBl6Zv9+Exv1SMYyP
gPEBbE9F2lq9WEwl8mifQ3mDKK+q/wIgPJIVOvVTj31ko1c5y6XTkBA7IeOCAk9AyuFlFVajth1h
vQNMgvvmpgR189w90ySU7CNWwdaak3IT1454xdhJt5X/7KrlrKWXgljjX6oC8bGaysUtny1jlqJE
wQ2oNnzKLFl5HkCE/Z8XLtGpvfIlWMLyvG2GkkRsMcBGzcTG30X8l6C5WdYwdazd0j33BgIfYp+Q
OWt91fG9OUSjHXIYYhIUPSwLOtnv3mpl3OdJG3Ln4hIzTlVfVvy7vO8p1NSF2otH+nl4Svps/j2b
+Cz41PZVKasYBFUUwtgwUmAHuNafu4JlevLJbiQsDW3/scywa32zWdacGBKb4fR4hqJTaWV7umVa
VWZkya2kDN3BeZbbatVNz8lWdiSckN3D2PzqNdzrKT2x/+4d8ezXm6jgm0DPCh43bVvukUCK30Zp
Cou80m3CeJ5Vonmnbvh8OarNfF56joHx6Hv2hCInRxd9Vy5QhyCVJ9AtSDKEEAvXyGvvGnxneZF0
lHRv1PVPFMSmkINe3ng04gmQT8WCXGYqUSxfiVXDlRilj0hcK9rvLFyim9bJXcV1s7nNsJRvNp68
eDzwmfcPpXVWmTXcgfQgrtLu8Sp12RxWdd5xKttRHAoQNi80f8J7OalQHF8oRvhnCIUEBgv1ErnW
EUWac6SjjS356FTS9scRup47SRrwadU3/EM4bpdxYbNB0eRbnGye9nAxzaynlAGeUsY/rZpV4GiB
1kMzS5eHA6jgMJ8c+k4iT2H3eSQCdWOsvMEnnj2tOiOBmc8/HxcJ736N0dejeyCxymeQ2OL9waIM
0vxdSxtfuBmLQROK+LtCSsAyw0U9aOwltpBzIfQvayO3zTT8MBEIcnjrJucR8HjgZfvNdveDM8lf
zuDD608jePNSkYNQlqk7HYwGaBl8I/IAgw1DQeAHlb4VRQRR0xaIUUTW72+NnF6bcJzobWnA9oE4
FA8C/rXDFyvOK8TYkp1+fxtVRpFG9jYQAOZATltlZnKkPyotok7ww2/LJxe6LPEn+2DytnG2pg9S
t173uvwI6ZumM0s0aJFpvxXAF3MsmBLvrkO5H4zLatRgAwMfr1qQTeuWRWNOYZpXdCx5a+O120/0
2iH9JlPbSauVsupJZ8G8KWPUaCZyqXw0RWJDkidV9iU8or+Y7t3lcAYPN6xlG3BrOQ0sbVgLtszZ
ANIPZ6DRABz31TSc9/as3MZ67SIUL+SwjcAuYExWs4hXWBeextiyWEdbAiaJ97QMzFdacZJC7MIy
BSYVWZFCzsri9FCcc+3cu6+XnkahzYMJ+AdKV16WfppxTzQ5f/G6+sR132cnDVMQaSuCbgNQw25G
y8fwyuMoEEziAqI2BNsaWMAZjJg4sDlyvhFSFps23QjsWVBOP2pXAEi8qHh1XXEIqnO3Hz3ZlL0f
ur8W4H5/e8XKMwGG4+W+FxuKNROkvvNm6iqnsjOKbrqeMkNHwiOPH5aru5lXAL36sI39v/vsRaq5
RjBg21iNc9CEc66dAlFGYyDdPC2pL8LVbY6zct9j93ywgZ9BLhgriOs4d8jfzNFeeNcGFmsAolm7
L2JnJaR7nxtuSE/OGaxCR8k876GPXettlxhywyaALx1IQoZMYKQkODHdgq/dmV2h+JauU4RUCn+W
DXKi/OOMlGP/ThHnP2Vz6A8Wo7ZM6W0XEszI6orQu+LU99j3a3DINVXDe3GsMfYGfTUSsXDAgB9r
uf/ixytM2uma3crftMZl4xz7ii35lwId+9DqO14wNyXxzY4G/hAPCAPnFs2d5AQjXkROeMh4f22K
cKJg0ORq4oXmQlUg9Bk6kdQpDjHMicHDxSVb+C4crjdCAKFeRZZ4Q79M9D9UgORoDzQXbdUx956b
MLvSPeTSdklkmG2TEAnXRfv3BFgXL2kq5v/uDZ8tU88v6yryVlyXcBplAM3dFDi9JqtZWlF3Bu+h
N4YR1RMimnZR1+APUE6zRCzALLOI5iLt4rX6Y4YG8owiJmNKoT8z1bzq09aGpH8c4+ASzGeieY2/
GyLWgujYGQcJN8irnV1LA7uigG0pFkYcFxy+3v0txyujyTdJ563bkGtecKSpTBO6o8LRGDukJ0nT
bI6QHkfHOp1L0OQ49XFa4Xky4IdM1uB/BbJPfbjabeXlQolMAXj97m8arzqu4QeW3DHVcmrkFgIQ
ZD70H1zmvCww6LxPAuumxgSjGNu3FvLaKNTjO0dbUJe4T4OlDdy4fVyHx+dhNpQAux8L4qo7zbGR
o5NUEEXYHUnYXz8c1Dj19gxYguAVmHi37n1mWzQtWEaF2Sb4owrVaLLPnlP5BkPstj9cdiTcnFJZ
RhECUrxe0GUhRPjWYtSIddk5i344QA/2VRAAwpU2sVUFvpkoH4W7KHpK8OqOWsBuRxr826d5ybd0
0bDDtuVeTdJKH6o29FtBT41z40FwwkW7sH1s+oxMvUTEDxkiOrTWhk7Fpn0K9caksSJ2p/gyLs77
PDuPNGLN6Sv3WKP7rWbx0d9GnN6B8XFlKTUV5jZjY2PHfyKiwJDxsXrAZ2WJu4eMlWrIcZLbfpVU
mF+a6AESNr+aPkgwUSo3IOZWlyfePf44yl5x69OIE4ycLjfC6Y/syT1u4y+829eAv6MFzMzkRCoz
jyrdv0k9IuBhmUddcD9Imo0p6kAVCfL2T79D4B9Kk3b/O0o2Q83eYdEqkuGVuQ5uf9UCPBbq7qRs
B2HvHvoR4qAlmLBITGg0+ORVhmuHIdU6HvN2eXVMDp/u89DKN6AanSJlzNMXCztoK3bMKcBvRghr
WJutse+RQ/SawHfrhe33dB1Pfg5jL4YW1ScCkQh1tJXB6dsyJ/WfLKezniBYEVHlPm0GYf4IFfzJ
lTHtEjmGH0H4Puq3/EPvqNipGTmyc74xn2qMEnurIJuaA6aqTPpFzW57S+FYOwXenPQ0XQD/bREn
TysDhxvdMS6RvOCaCbuAl80LmZRy4x4nimja0l9gQcWd5DqmWa1r63wd1ZWQDmTTeE4uyas1vY5y
yliOMlJQhiiJbkyGS7lMltvcuUjWiQYsyvD/FUdpjt9x2qv2hbbwmZNkp6rXWmdpNZWZblUB+zrv
Rqoll9gSkh9GD3i/hcx4/PCRFjDmAqb6+5N30NWmol7ywc+LfTooMtYdeXuZB2fn/RCKz+70xCDh
8UGwBtq5hYpgIgK/ByNAJwiElvHfoTqi8ymRxVk41Nx9NmzUYNJoIvyc1w7Li5fUKPLbtw02e1Sa
MdxuZtc9IN3xQWaqaSwJ2y7c7v9sDdn5ZXKTkzNT154AfWXr4EywsHALxrwtOJjLDUx3YSCzwTeW
rvU35jNhcJzICe3tHMgjHY0aVqeiTot/LjEMjTwduXvkAUUUqqQT8ZZygmNRPmVRz0mHmK7Mh8p0
TdDt+ysLrx3yp6b9IO5MG4OuWjNemYYlUTuhAjzsp7UvhuzgxXpy/noXjzS3SAVDUjdoN1FSYZQy
BDiQHFKGqx4lsq7e+pRwBzEN87q9ddJHydHepsqV6oOiAgZh2Bwva5XnPDbzcy9W/ShVenPiBNL9
2RqepjiPDelH3B7+vhry/R6g3Sk4QvO6/XXekFbpl54zuXdROXgvbdyj4gxgOdC+NkuwamoYUZDR
AjUlVbaIhoUPgWS4guAwoREn5+S8rJe0Bq7kBCcyA9Z7JmqVt4gC/NYdFq7J9k5jrHPaILwN2YVo
OCYuJwNTt8vjRr1iiSErW393No0WyqDS7b1cjd4DtgjVaw3QIwh4O6QcA3vRS60GPPI95Z4K+i2T
Uf6nGNcd1L3nVPLXAEE+vd0UcMYkPuX8PAqklUA0y77Q89/y59HSeIchlDAcfB4iX4nea/F9kaVY
aPJJ2xplsfBnI87eTRhCswrVifsNUDqzCLTm4WjFuZGOTA17pPzQoEUx0mg6VVEO+EihKKMiZL8r
+VBL36kRk1HQfMTGFM7blviyJlQ82ebXRq88yVaGgVnfzruFBSPWdgF7hFm8UjaLizvdHUKtUXev
quGeeh4yS7tUyZbAOAYCaeBduaHH+emqsv0Hz8K50l0OPVKV5xU83FBL6kPr8pcNYrhFtCGbm3tL
JztOWB2MYWjQYxB7QhiHZjQw/e+l4tuOB16e+44t8OAnkghVPJAIedPMTHfUSHCO6vVRak9pY+uu
WOmz7FnpTnTVehmDNKJQrfRbdTB0crForu8gRGj1pq8AAQO83F+WsdaMdmpXhVU7lJuD+qwXAVcp
8XEMZIjj6j5Q7qnGJdJPjBY6TdDoMubudd4BNVEcY/+jIQGACbnmZMunHzXKJMmdq7hGoa3HsI1G
et3k70JLuMKEYIboM3sDy/lT8xC8xiz7XOuVQlWrpHbynCvUoQYLXWFSTz8iClxxauQ7ihDPa1Os
fvrXiw7hAG0ouERTTK6zb8n6V1rMzCpOQcUgK9nz7e5PVJ8sAqY9IHQboHSgl95pVNNiaJ7z4t0H
wVFwyiLNS+wJSk6jmvQtZLA3aEP4AoTtTfLnSkgfaU8qdgHEtJcGeaJ+aIQGkKQ5nZjI496mUDQC
mHymYmPllXGbMApEKJudNusQl6d+QXbrHWmLj2g8Fz3I+TFPBHvVtlEa5atixy/T3itE5MZavmC7
F5jq9KW0vUk0p4xPSBx0QQZrwNcNi9FkIaUOKdifvABqBOUTcHk0pdBLwPdrZyhPY7l2cV/rCo4R
ZSMdYdyyoaScLDtE9x9KTNAnG5RmV+DfmhaOHyYumIRWoKjUmacUKPDHqP0bvt+6aBWqtdFicgy9
w30IN1tSVc23a47gIDoqsD+jW6zussQ52cKs29ASh1+G4LKyFqcfy15UImxOiz0BmI6ZQ2hkpHEZ
gQOSZW9xGDoFvcWWQD+ggLSP+ba1ryAsWuyCVMduhHsvPBZy310bfp3sg5BE2TxIWfxRZugv52Rb
5o8pGyuDOOM8+CYbR0UvHj31mfwE+XTgkHjUuLmuuWfoepN8BO3pzs7ENHCLuPUWSkVbpRauKe23
5tzzrbfMNbw15IWFOJuPYJ0Ujz++jdXVxqxnHGuaScovJk1JXqE0Dqg5t3349xRS3yyJUQazSgZQ
g6C/jtrEF3uiFvoPOhbELvUty6PHzoOok+2wo226nJWfZ12WnlLalZJq5bnJULneJWrGcCcCuWFo
um+BREniw2Sj63yrqhJYVQ+JTqNtcWH8ePKReRUfbFFtwYvoaNaC7V/SESQ5uSpkbwA6DbnF768V
pJIsWIHxc28xU59sKcKaXu26UV/Lz1tb2P2nDP3oBRoR009Q8sWm+Iv4e6Fx/pGT24D7AhedUQ8o
WjQvGH88P1mn5BqQIljx33picEzy97MxbauON/J2JHivd6Mi9Ga15bOIQmkzk+eOpzqyuGfZStO/
sdkJHsBxu5MFPvnrxETvh/Ns4kkoarGwvT0hNCOY99+LukEJ6IvUQN8mTrnEofUZyyX/9fDnmCBD
lzyBa9jfpIkepaBj9Zl74Cn0SR6Yda+WU/STwEMze9Df5X7QTTdKNjBjB5EkqEV8jay/85SMJ40s
ipL+jCMWNXNbp/AB/oP9DT9sJMWPc0g1hpCGiwfDh1GfBRaTWMESLXlqXSVzMhXu7B4KXjUQQa8u
TYpFrfWeRnl73WEki2XDDq7RA9RbRgE2QLJWLb+zFoxej4wScWlZ0vQ7/XxKMseFycoxgwEQg4+E
v8J1UZK30PeZNExWByCHTXppafr/17wyO0L3v5Yvv/jc5V5JOAqHpRHY2Nqq+xd5cdQsbGVm9atS
r7ctw8xFq/dEVl5lAcjudJ3F7ejgIi2NAznyELEExfF8Vxm77duNQvimy7iQlw09JMIBZgFM0oL5
sEM3XmD0Urv/R3wOfRN/I/B0k7hkQzLosJ8aD+G/9L99tXej9jVaRJDg6keJi8EAE5vq3oLlc8eQ
FLwBj3wG7gj9iihUO04rV6faOsyxROcwS6pIFXcYRdH7i1pp7YOLQrN0xr/PJY1ZMKKl34b9yqRk
f9lm1m1B6E8uOlNhmoBmJqtOoIAW8JjLOg5uHhFEmUE2xrvfYescLNfUVkjecrpl1TkJx9EDa2ZV
Am4WnusSIGvj8l4RT7qt1z/6xdb4WauH1Z4BIYdknqJjqXOzl2rzQP2xiFtpTrtfYzRjV5iKgcfp
EXNIgTlIF9Qp9VatLzR+LC+DwiKu4MmVE0xSLgHOxJnmgTc5MlcmnnpInj/h6KbRw90/uuy+Cwbv
JRZFg+rcmGsyP/Urp6C3Za1Onqza27QNGysf/mxodEyTQ4WMFaLMaHj8+WLjyfXxY9wyUAbtWbMx
C386j3zQd6emTR35ZMxG2FCfYXc6rydkyhQxQLMTjeeE6zWkO8cdjk6K9K9UtlomBgKSXiQuDK3Q
uOyhkj6pAmtzdHhnrDmGJRO6XvRoyanJGhYE9ZW1pJa6hjWrQ/Nt7iEwewcuFSOFhUHAP4BJ7OhA
p7wWhlb2Pk43ux7MGlZcZ1FJfi1h8qwAYG+HhysfLDkQfEFhC1J/TbFKxq/QMrsC1XjmkAHr8XH8
X6ms0MCArCfxXujEl10GRKS98Ii73Xsi6ox5JY3wqukh968lGe1II0W+TkaSaOJz++8iKF0JBBUd
YLswiC3r58rp1SVmcf52XHVqVCCZ7aF2TKPnLtop4nzsz6CxlVqEm0iDNHFHkXFhJJ2Ij8uqcRJC
rd2xQv7uDafwpS32J3SCCWMB9DeV4v6xduJ3P9EfT2Up1FdYObGHnqf4fWWx0rcb8JWElVvneq+A
PCCFsHaSXGmQUTNTFUnNvy+ygPX6eKuleDaV9INT21B/v6z1T1Gg1J08ZoyGs4LstctEdigVLw3M
Nxs+RzikoPPKOX7kg0/Eoj2LOJ4hHW6SD5OTvF68nYDiz/sOREsLm2sKzvY+dtLx0bsOM+Ek+NRS
HNR3wd2EQMXDVTuuYJTbJ9lgODkYmA8BqAbyGk0P+7iEUgdI2beORyZTLjQBIa7c8LdNop9iUvtN
3m3buRXC+R6/2rU6K+dG+aFctdS4LQSjFlLUFysDfjDnU3mZ2Zi0htYsyQepj1wecPlsWwZCTTOS
8bJlRtQ8M+HkWvc9iZDRmgWy/K/bFyXLvskfWNFP7t451DiJrAb9GPztrKaJnY0Sf5dT4aEyFFOo
LjtDh6HJeVvp3s4OdAczjZ7VDzHMQo9bBLU5JxsSqdVOtYslBaxvVIF6IojKei+utW7PXZdJgS0i
PSG88TNJlxvNd4CqyOCZek2+SfD2mAAbXfiRkw9alaeQOhWyt/qUQtpb2g2vFbnIrbuBL2ubLZaf
azapEZqTFr4nSTCitzLdLd3HCe5hSCuVEwCL1qAuiEbhXBnF/z3XFat0o1LJdmNIYiY2A7OeJsQJ
dkR6i3jq934DFMWCJWNbEVH41peCtk3LQ+FpUcwQfhb7mX+pKynidklB6ntv4pT76b8fAS3Cf4Y9
U5yaXcLEFi2lfGy0SGXCSKM1W1eS/FyBuoP/EV729aikSRAkZ8rrvcVe0B22+BHy8Wq7j1sLGsMr
r2hTJQZ+kruenRGNIfmOMxX2PdMmg5kkMuZh1VziTNDRgKgTl3h2QJXzYv/Nlf0xoVA4ARDvTFB8
DSK1yDMhXvanw8JnLHaHFuAbTGs5x19Y+iROJ3YbM6euRviJ74lx5vIvFKSCG3a+bSEMirC1TnwK
L5i4W2nPcTtSnxk/xK8uBY1CMCDmWp6suLwKkT/bvvB/ghlfYSMTPYwRfxTtsycmUlNq9kTrRRVd
9GrtqX7TCPtSqk4QwcxV2U3IHYMBzyuA5lm25EO2PqmQjpezoQtUUzoXsBO1EP5qBOQ6z89jMZ3H
JfJ3oTqUXJuPIN7xhG3L7XyGhuhKGYZ6jrbSJ/DAPpgSbz2igZrtGQWOi4kYh9TUa/wak1vyHQ6y
HB+Me6oWbNkx6Dy2sGh8jMDnK18w3hFQ/LEDmtBVKW7XrwgsgNzDkVVkQEjOgJrL7A7ueBi4dU6U
rPNvVudRJon7ZOR29A3wbIW4ncKOxqGG0ScrFreZns/oja1cw/BJqhs6tBOfZxzJPntQv7om5fu2
AaPQndaEPtUdscaXwIWuVTpqRLwTynnfcQhw0+1D3KNnuWnVaxam12fNSaThYjkaMx/jHcHyDCTv
48aOQZiYFuhpg23clLc3eW43jdipiASDbjyTRTWjGSTjmoC5dCW/3BaUL0stkXk7pLNNbHp/RmFW
9ZkjBXPemQHBSxT/m5+MECPrWs8l7Yg9EO2VZ27Tv4xOQsAS3AJR27U3JCFB6iZ9BX+9A6YU+8oD
LXMfF3OJSsE1URXnEtLrkJex8UeqeyXAf1Bfy9nu06F+Bn7oaIk2F2tOmXzG2wLNSfN5egLrEOk7
i6UjzG41t7PV23YSBrBnA0WidoH/eSfx2fXLD2DVGWhhdvHVx/nQnEnRuQZK9y71jE9fSLKX6UUH
me3FYSfnNEigD4XjlbuDXEIWwvR+AJEPf7mHqO6DmvfKL34aCyzlS2KvnwRI5Uy0/kPhePP7GbGf
AXp3KmIbqcmCZAIyPWpfTjMwwRzjRYsIT1wRkrYWAKeHRbMJGp6yYAqsZ9ybkD8VRsSfJuG+Zvt4
uY0NURs/EYzWNTy7pkNUsD6mIp8kALn1biOOns509cTgtJlb3YOKUV6dBAMuIOsgfZBNMPO1ZbT3
OPwCY4agZwXY7Awy/15TXfCIXnjiXjCHMNke41R8muGZLob5qVFZU0B7I4yuNn57nR5bebvxvEph
4F7n8nIQTZBnP6vKYw0OxUbzcV8JJuwvq+QCvFBO+T/3j5zU4A7J3kaGsUEA+TY1tmD9zXeAqzxg
9+5R+m5UFjMqX+bSTwWpPy9IbKXlWiRqqjEwVUmoTKAtyRcuN7wOOACJiZipMnWWG8uG7BAh5UyD
Jj+CqLMXyE4vtbta0ALEyw8jlSaEiq6JGVN67hOZRMXnlDZdicNsQSeYxD9u7nzEkcNFrqt9X4za
NWQdUjIzPgKB5+Q6yYFsFLp6GpaSLhVScqJ/mCWod6BNgIOifzKZjjzokR3mvFKDZaWPxdqq5VBK
J9cYtvv9uf9j+U1xUYUWW95NJiJjhbEfD5kFqiy56X3En+gxAdZ8goUYMwaodpUXWOz18uzYfj61
0v+ADfsBhJb+k8QCrnPe/oZpaj34PGYCMGIdb+CCHtSKFgHKiozAZoMy0pBb+Dabojr3DfBHT1jj
pKqA9WGOUKL/pRlfHccEgkzBz+DAQTAiRKwnYrl4y2mHytLq72q3l/I19pPXT6Rz3Cjz5O0cM6Ne
MTFLOD+bKLo7BIw+yqWGnyYj/zZrtsrObCxeNuaaSBLyz8tiW9M9ANS+EdZ4qezgbU2zhCh3yENP
evPEqQAqNWMRP4t5WS32o1uE3uy7q4YHttzbBnWsX1Bd6oLHr5NqYEKVCvuDc80aCn9ddLHDD8ld
iCNB4NVd/1Z6YY9bBg6o1WLQoNfGs/7yJQbUcAQWhatXIegpSPBc7sdfhaXkhG3yf9oNBl4O/ily
DTKcBTrTmkecdxuP1PXYw9p1PJGltT/NhAGKIpbYPlXquOlquQy6phl8S2fkt8CorMJRAR03dNMF
L474wnG9i5XfaK03AdnJKNgxC4IZyE/LxcqupstXODE3H1+BUwO7Rf+3tk1Fex5jISSWzQMDONGF
9MvKYAibhN52bgbZsquSbVt51y8PwtsKSCKcHfoBRx06RgVy/RSqdhMbJ2Oc8UGRnlFB9vdTMyKH
MlJ0Vlj1g1mIVnjwF7fcWXxAcoG3l4BWVW8VDlhnDrODhJ9nV5bY4sOm0aE9cr5vjhIILw9/D+fM
j9xSLa/Yd86At0OmWUsLYMddKmkRYYLuVrAy0FhQuwivvkTjYagmYKGWtFX1Vh9NPrEtTMKGMvOm
Zq+mNEs/+ShoRsKjZ90ynEuKBQTtEZXf2xXVioIdhwCd20FAGDh/6197FJ7Fg7lgWGbM0XY9IPJj
M/jQIzWbaxi6O93AqohTdWpHybtzYrck7eCPmpN6dQXIvCn1WJkL66uMU1zIUNuFqVTJG7/3yv+V
E1AGECy3CXV9JpWe0i/3z1WiH7CUpv4F/Mq//UZTCajjY74YbDYWkxFHM26I1OClQNudIlH9gIIJ
eSWG+rIV1D4cxs4MiuUyBTmb23SR0kTDvcvVyA903jwEHrwA7eBYrLvVDcWSYz0A8k82Q00GXcQN
bQAi0cS4dR4vPfhQVMr0XL8l8/pxlwYEWL1QgPA6UDG9e+xCEaxq8puKcPattg2VpxUK3F0lQHng
Y9eCKHkIhRhvMCk7cILzAZQIftLoeG9oaCNNCpKfNXGbPQ5QWwqJQP6rXqiSZzpS2HdCGK9ob2Ts
hp5UiNprk5JMKrlUR8lzjmjybcsPtUvylhXEFhfWC0e4SnlLXvs+eElS8BU7XvDuF9KQPJbeA9K0
MjXUKsTZrASnENjOuv5xka0Ju7aru5LFYy28GRm4cZ6/k+G8cLyvJZLE/I8As76xBVtyN18JMw2Y
8vWy7BW5LJ2FEcuGUNFxKpD57xbxrtKE3fu+sQoLR6a3wPw+i4c6bS85QJhe+weOIoGau2CoMKPW
XDk6CQswA/MsOwAuKhJQwCP4+jlr7J/5uuKZppcYScklASWppCCUNg8X2KfmRwJkICH9Dr/Wfdx3
9oiH//VZFPi1wxM3kvI+dJ/H7RIbha5slMrRggec0vhoxT/xHw8yWxVvLh3m7oQkuLUGo5DIlgGA
rumX92Rwy90k8QR1ya9leRsK1Im8pVDu2eRItLku/ZZsOThVPhaWOiBzVJZ5inTQMWpAs2Cx91va
h1xnv4OPqi0ah+rKkUQT7VbYjUknfPxWxg5fOx78LmqUnHBNUGwOPLtQa1L7XMkmLnFgxlVUVm4k
Vyv+vjqZqczGpPEzf7M0YIrIR2c005bQAxSgE16as8X2wFizSZ9u1rIv7XHE76AvWKaGASAfUqWM
xoZ512CH0TimuVrRg2r9m61BOmeIkx+hyV91ouJO8Hr9HrSzSeVoZpe/UvAszfHvOfoTPJkwJEwt
6A3Nje2EP8Jd+vi3CIXOBjZdq6Zx/kqk9yV12pa2SFMVMtQpnecXhDqcz6lqRQd3wzapZZRuSdnH
RxjCkRsVbvnkackiY3pvrXzm3WwjiNNLU9wyAXi46GmKW7PUmHZpcCCYsCHIUK/1mAG1GRND+0MF
Rn1fRTdkGbpA8BtQiVGFy5AgHzkZDTUY2ivbj7sWC+Dp/eC6t3LaaUl10t9+2SWjCCZ9lXUCgIo8
KZKf/T7DmrTyrQr02TZOwhk/KBHIFhXu0NDonjpofLgCwGZbtJaXJLgJKafCjhDFjdZLTka5DNC7
ObVm06emwp3E2ySTYzdg4hUbLN18bIn2nxQwHOaw0bhlVDvGibBfk3HN+5bRJXFI6vptwj3zgV53
fNDACZAE3OL7Nc1ifsE7lQSsQrOuD5X67uNAfZzvModL8DMBKveFo0AVVL/4kWSpQ1s/hFlxhOk2
iYZ3nrearw4jlrSpQLxo79hk/MOqoMn2db25HqKZdAD3NTwkrtjUKP2bfV4TaSXHyOjv8FkZ5FvY
AI9KQmzeTwBEVzcsp6zY/BLp3OVmo2lzC+0J9T3RNFBqojTz1+FT93hFlLu9PSqRFVa8jAM74xCZ
veE3eG9AlqCYwX0mpDlTyXeVZ6LvyguZnPDKfGHHV0kC17aIkJppHvHEePlw4/CvuVAIdQJ3CWCX
jZnrNcm5w9ioVKqP0iMP8jpCwFfoArTRRhwsmiZHUJDKPYkm6lnJUAbMHdhAcnWmsoE7E8gCIbtF
kPNiZlSiRFlz36OEJSNVuHEnFsS+xO31e+hapx0ZfbgG0rMZr9ttZ8/HaLaApfJGxGWxJDpr4ZOD
82YARMhS4dxbamtZZkwpU2zz2g++mtaNmSNuInAE/cA1Wxshjlpb8mUU2i5zdPEyGISW9avS5lxl
YtnItmTQWerBEeoNT76YtWc35B4HBT9+ngkovmgwRdt9hg1qA+/P3QBmGuM0lPH1vD2yXenrnWeS
jskfBgLXmqZW0Xlx+msAhATv/1r1UlNJVGCkZ2ApSIiyJGE0BI+R7HL37zhKpNIXSS6JzwO+q7/h
tzEgXaJvUuwMk8Ts5dsnCPpqCELMHfHiSJ80UDDiGzXhv/c3l4tvHIlU2yKhYgwDBVGRTmiQ0ZbR
/Ng5YJwkLj1IIVgsuotFJTpaOvkFQzxua3qup0WoaCWiHtlWoOvaqoXNEPJ7J2OD3DkS+sRdfSYF
wkvRZIw1HVZztJELE0AyqtzRuaWWx3iPbp28SgVURghxLZloiZxMtxhC8HQbLoblcDXsCH93zB5A
P+QlRVRKk1BYku3TR6KKxcJBlt3noSfTfimW2N+MQdgw7T9p/P/uUSrrJm/6R7FToahC8S9X6ogV
7DOt6nugVyKq81ijDSQx3/KZNJjLdNhISYGEk5XSeWB584HcfwuMH5q3TqriPHxcDzmqR9hOgY73
CjWkS+0f81t3RDcD9wNRQx18gaxGrhTijgmIiB0irIs52ySrwOYVMhawWIeFqQjxb4vlOabzhDvn
e+nT7yr64dV6KmYayWC+FtpNOy2/BoJPP0f9eRxKh9eCN7r+1CFX5MSTKvw4b5qTsepeijzwWfna
Yy1y8d9DprYWwEeQnokUL7Z7nhTz8CgGHfU9intczBRfbYlKofiebnlLtsEJU4HGLY12O20/HSZk
MsaMHA4OX18iuqD7GU8Ohk1mehf7i7lrpipLIg0iEdzOGgryXqaxT7li2VJ9zAp6X38EE3NKpsZU
AqHNKbAOhkf2LLmzwItPEfQb4Zxyb6t1PUjXXmL9O9i5aGj1Tm8BuYlT6IGf+ePPylv1P8hwA0AW
aCv6DLLoDUBO5VYlRhShbHWedYeIstIyh1DAP76NPnDlTsY1env/bEF0oqOTLvFcljh3h+wyLCka
K39MwNec3gkUsbuze50vqnjrZ5RbTkE4ujjNWGItThcaq7oNDjzcVquGg6WQ+C1buNircrch4CAO
ct4dJ7E14ojGIpqcgIhcwEqzuaZel+CWtchw/aBaK9ETlMTGeLsB7XKA6qyO25IIk7B5eRYsWVnQ
zp62yYlqUWTidyJn5LYKRb0EhoJnllWExRQTHMU3IGPADaOFjB3fOOVAPKk7WCjtBT070nfAJQzh
O5EDUMUvsV7NgWSwlnlk3fq4EnNXJzVir2HD0rv9Gkppc9WzhHOWixKwCUuk1PRzmXoJw4D3EMQ7
Y8n2lBEJOgcHW55MTid5EW3Epkv2iL30FvD/e7cYi45GyQhfLHoAFQu717T/OozE720VL76/zCi8
dxXZdU+n2khusT3MA78P1DKOh5bUuB2tnJJ2obkvBmSbty4aw97jG5+hRZXzDW9yL0uLENnwMOoP
8JDxjKOfFQ3Seo2ObWcNDn4yibNIERUu1eg6MY49vok3vzrfSb7+e7uC/9oOmVHj/xuIxQBLaDzM
OYl6r+rjsHmtKPf+psJkFMD8kG6jRCXQn6cyGsuR0rqhZ01NY0xkrFGs3FOTitMtnQdpV80TTiT4
KnUQQl4VEskEPL92YowZJ+F0WGGyg9+vl4epF/DQtOJRhsIzKaYfciAjzIUBYeV2q+NL4UzPBqPh
tvmQGZVNzgfYAlVE0EOlN52fEtWv+9Rwk8lGCKxIlqKECBOovxZcCw6y8QGiguzUmz4fFnRbGhK9
Hp21IfAUBRo4oaqAbK3XTVG+WZDxOPFhcYnznD5q3O0qVOwrMa2gvjDP9sNT5ttoyBlHeFk2FDzm
3qz2vCPdu5JkQ7cGuLi+Hc2O1sf69LnIk7aMiXVa6HzpbPu6Bel9+17fuc8I7rYI4H+rH+yERxLr
IFWwDaEuCeSeIba+WX7JdubpMF1k60Ix7WA84pOMCUlssQk+/QtN7nU7OZgkqwVa+WRfr5Sx5Dpn
VZPkhn7bn8sduFpPLNCVu+Ut/t7WyqXZ/HupAOTpl4PO8XmodneBFGjKqX+lKH/aqgNVyUeo0Voe
Diho//g7knK4pby1eIyo8iwp4V+2QWJxXWvruH/pC9w2NT3rL6N96BUDKYUE6hDESUZ7mOswsX49
CzeE1ysIe1AvmbIO7HrajZ+c3Ow2H1kxqdOMcxuvNQKBf5OKMwsAbiJpQVdM+RnrWqYhsXr7B8QA
EvJeXMTwZsB8tlH1xehm3V2G6BF8dD/IayRGQQqgkUpEIrQcxdqVBgnjihWBR1gzp4d/Fbe3mNTg
Bq5yrRGXVvDY+buMh6WWYZnsmtrb243EeSsSf0mcF5Kad7A/sguFppyr9XbKZ/GKNwHczX70z+nY
Ma0o+43cQSlTUUI55jVAET1A+QlvI+xYHgRWwhOvGOsHxHeN7prBkkhsDP0TiuY8BY6iztqSUsFO
20L0kTFued0776CjeOX6qwYUj1yy2nwCZtBSHxdxlEAg7WacvuJ8K9yp3NgkpNqBpZkM6AyUVpXS
bQK7joAA1AnDQF16Mnz0T9GO6oQvCSLXcHUb8u+QL0Rqmc5PPpPKVNAA1ZWjnWmj2xyc87KBjS9A
XhkA+Ok89d7hVMp88xfVMw8CmbOqULMDKPejjSNiHM+s4PjOQsQoHcfHuLx0Hfc84Dhz3g2Dq4fj
A7Nvey/7f5VfhVJyXM9YKa3af1PFvFTOzjIL9tkJkTXUgYckcyyoTG6HsAzjhNjcCk6zRza6/gKJ
DlPyvQi+oI5W2+tC133pYNsIhRvZVyf5b+OUPKzxP+M/142oIk/Z12pBXmIkN1IgnOhZGeKlrDOy
7BSPXr7lWIMaAPuskRoftxZ3Pv51vqdt+qgi9ifaH9kXtektU5j3BuxzaeK8YB0dpqf0eAc0oxA0
PzhddjiHJmoLuC9S7NXhTHsniqg6mXvzhkxPh8MmvMeAMUx/t5wQcOn/UwSyGF4guaJcW19SmLsp
Nk3UIsxRLydaEiz9ym3EAepGE056ZgPv8JYCQePCGEkonOatuADt9C/MWHUYh40v5K96ARNmb2du
cGFYU7H/v+eWLIEulqY9fMjbpUJVfkKtPfUl8QyJY6LGJMw65nZiMy8EwfMw7bbUUEXIlyfaWQLR
di94NU4dV67wdGS+ZJDDkSYQEChi+Fjn/P5pZUXq2Mudre+ut8YjYxolKfQOVw7I5Z7thGudjimI
WBfSfRcx9INnGz3H9sJsOaTW2vMlbHXm6uM0V49/N03hgwe8n0iuVnD6mJX45gvKZdlrsboAZh/J
CgAVIuJeS7Z2RgsXEqiKYTCBv2d2f1ZE3uFmmINmELYq8L7IDV7BS3E9pfKIOTVijPVYAwhsePcK
LlWOJW6q3XSkZkgy4LCjfPF9ATsWCo+Wm5DSsDb0Y55h4Ot2AM/CpFY2B4ieknssQA8Aw+RtruTc
DviU5flqM8Kivd3KdkG81aTZldfCMnomOX4aRHPNs/ftAT4jcYeoRgUgnp6xgVjWakyKQQmE0T2b
UbqeTNnuRsbNRIgakZdHBAgrAF85XwHwvlMwXcMRPpOxXFMBTqzcUiWaURm39QDbmYJOlnGIhE2x
xo34VbJv70Z2AMg06+wFGylMzuZoRmxXjTY20vDVfx/ED5HdOnWIjr1qSwSdb5FX93EoqtiCiPvJ
okj/rJIwuzAXP206Lbq+X6U7QTn1gQ1lVA8qfzl9MgQRkPfj/4swqy7FZ8ol7v7iR4GFBYoF3z4C
taOwbAGW5eIdwqy9nwuAhD/f+/bQSa4q2ZQ/hIU7ROzVHdu4sR9Yj5W6MrYtJgAqEjazT7eIp6BV
M1FdY7ujbTbXNIZHjjjMrTeGQIBIFETOzAgNcnbDeoSscyawb0jYYp07pFKz/yWc2A+an0HzEc3I
JC5OwfbW3TIoLg+QOXsEQDgj7bBqN3oBwvfZTQI8XTQtXFBEz9Nmu8Bthoha7NECTAAAplJOndvU
fFTIysntcvdqH1mc2KTwjmyLVpEQbfQeXyyVyn55neYhF5RamWwn6FHDA/R4lpj5gAdwAvOkI/Zv
jqj1uxJwV8A1t9/RmcmqCHsJZf4Mdyj6sA9UhKWzEGMpERr+fOleEUUCmeac77IxrBwhCciwBsUs
Xb/s7QSyDZbjWI8B6ojS8Zo86TMv9ZxIBgKYQ+AZO71sO488zZwFF2kI9za6pU/vwkhp6BKM/Lkj
lkCvrKC+MztJJ6iuMNXY/Bo1vB5jwnOyIyRD+vIHYUQIe3yIfj7lnzSEkKFN/GWZi6R1qAx9+xA+
qqBcUYS3pGcvq3DdYvnr5GAEhc+m5vXG+IjixOXHjarOV7Kqwf5CY94wzJw2sejj4EQ78r0e0Hio
As9yBtTBuxFXqcxecdrRRaxt9Sj520G0IIenf/7CV7cD99tDY37n7m3yxSJbkiZuhp0oi280PNbE
XtSSyHf7JnHUaVCyxyngRV0BRyiIhNdTxAm/+Yd3LlWTwy4HFPOdM0C4x3mW9RfK6GjWtxobtEYp
kN2dUZJrupo8gwTE8snvS1SyX+V9/VTQObNQa0VccHdc4uJNo9e8RiFA+QC2J9cKCsCXs1QXIaLs
wcx/58b0LZpZpPHKCeCZ3brW7rx0WlRAIj0Wv+Nwy8YfuUsws79ClexHZjGf7rGP5ZIt/ZQ0x49p
92kRst4Z6UJP6Ea63ZqUG1wKwn5CvXgvmSMaHbg94i8rNIQ+lLBWIWJ/RpQCLTsk2L1Xua4SuAsB
skmqANbvU7RV2m1gJ7qFiufJ2PkLO2srG+sNvPOpZKhbQr+td0OrKzw87+I5lXSbyZG+PBjrsIsl
q17R281awTJheZXoTo6VMEFPIJ46ZZYRN3tWlS75MTWn+15MSlwjCnxBEYKtuunRXuxVGPz+kXtT
MjEIZz3uBlECeZn2mL3NUdMtd1sLKVxhY/X/GGmOCT33MhcVxcMvXoIP8WaAjrdZn9gD5V90topR
wS/uYDEcb8AT7Mr+FJlvHRVvSpRWfQu5SJgOCCCcOth1aF/cM8NeYukfdizeuhyr83P80Gk6jcaA
eU0mlFQtfg4NBP5KlD1aXSkHyy2YX6oIngsPomtZdpZJqwMfv+Jp1y+tq5iOZfzm87BFTAhxT1Xb
v32TGw8HHuc2+wq4sGmx/5RbQwEWxGnPsucUAckcZJ87Rq76oUS2nxm7I8i7MrvKUXf85eVcfhmC
oVyIu8wY7l28kz7Xgvr3R7Pl97h2VKqTIgbVzdWVTdU17AdM0oijTTd1RvjePjP/RaM5TstBA9aq
KE7Dj3s0dIbyrYN9JF0E5/Yyy9OZyC3acDRUZnPDjXVVBJWLYA7ZmYR2/pk3YfBmrpZn+PD/b3/W
hKofnuk+EXrskcFFzTcQldY1pZbIidEjvSadWSaN2KCSEg1Bp9ECNB9lFQ/Gm1JdXUuW08hf0KRO
xEvrGrdf9/frLkrw05yVw/bLXFK7j+WNSgtZPsHSzCsoK2p5MOPGanAkj3fJ9OaAoi5rLOZqcYDR
MabzWLTqohXbx9QO5GUxkRu/rxyVvGUDWkzWndqWcN3UY+FQh4a/Bi4RygM0R2rIEF1ikTd0Twmg
g1Jb5ppVTOyLGbnZSodX9Mw1owMcUMFvDi905PVuvI+WlUJzICMXlxKVkNNV4pSidZGvV+VHx+9n
oqogV7dlYJ54JeBt3sSBDY4d5Pyb0pq9u+mO4D/een46+xinRReFnCL9bQjXHhqnm5FUBvC0fA4t
nXwbG4xf69zZPUbBmw/oO5MasD9KtHHYThUxx7fmoDe/7CAgRuf3i4oYVIU0tAU4szQpnWbcbbat
xRXLyAgFbjMwVgWHRt60se4WyX2gEwD+Pu6jK4lLKUMKQk5o8AxLzAPR7YAQ1yl6k9kIetQYm+F0
NAMhJLZ4oA1nyXPxl3yt1j1VlTq60mpB80ZaJPZUWJ0Huwt2rOrfvPZm2L6pBSC/WE2D1EySMJ83
/+CdL3IudT2/ZCLS4pCESz6Wz/jr2AmW3Tt3jqNH0cGiBbrQNyNJTaUQjjkyb95TWj8KUqrTHG65
iQGees/mRbiEKXWex5QWyls8VmjKRc0bj6JZDcWwGy+MtTRhGcCHk//1esipBz+sTt5X3DUqw3GL
pxHFLFcPHes3Hib0bMgdZKsSLRPu2XyLsxeZi0MlDpGBHHbwOGoI8jmdrLVkOPt6o4kNOCmUeUww
7tq4ZSn1AHvFEY2nSEmvNvjUtez/tMY9TbKSltXsD+zN5uXtNnQFUIf1bvD9QVPhN1KQRoBF86u0
i/NGlxkCYQzlbwCxEXlM8VBnUNCjVGFH4ADRnEFbz66RZBv2aFBpA9t4HMrynk4reNRL7Hxtp7pp
k2TMlilB0D/k/eUMz88DRZkPcANp5O1c9UwBhc0+DjhL8BMbLOUZllrtkmY0jR5U8xTzuu9A8pya
FbTCxdSDmLafXIdkM4/W32Tip/LIi8rYbQCEcjfufpHPhvhm+CtaKHW3GHCZKDN1kQA0OuHu9vZg
Jhb3dT57fQDx87+DIv+k08TKoYkjQPVloeso/c9sp+QTMJj+dtrBr4Q3385LkcaNoNJPnrjHDjCi
3hNqb+FqxpiFbHAHogPwYYWdaw+D8mXJ7p7ls9Hdhe/8nh04QtObEQTeEAQPbKaq1mo7b0XYdRCb
ekn8ucyPR0zJSOZ0W8ogugH5rCouWc2YixRsSATc5Jjgv5VkCmJ/eiSVOEws2iJG+cE/p4J43hOV
F6XyHD6JKl/BmCS6qHtyDq9vnDensb/ykKgIbDeAHQys0bYpEkK1mrPC3pVFpKzDnYEV15noyqsW
TWNcId3Sj3mb5bfLv2p/BZw+eyi7mun2Ll/wHmomB9tqAkaV5jzMnCQcAhLw6QQpJJ9HAloFfnUt
TNvEkKw2e6CJE8yS/NYE0/pVAeNrZNQIy4WeZ2umYXr8Jlu4L1CNkVRNeMS90btfnebtubK1NPiS
FR3PTlRctw6K01h4YQb1+hXGAZn/7s6yskw44fhdPWE5aDIKAex5fuwhimpnNiQGUNmojG9QUJXR
vCC/hEx/8E1spnNUPGhMQJRc3nfinjzSVQm/QvjAYwW0nsRTtr3VpvAmy54IROv/Y/qspMTI1HM5
TVD/eTfPzLTaXdRMjFKu35eg7+3fHgKzO+8nCmxjVG+BXF3hDlWHAmS24duwN2zigyT0s3RxJBBM
CjUdC5iTY95ae56x/vencYcf5mRuPPn9woIydrKKxF9GojSUwC71xW0M2Q13O41Ib1xhtOF58hMZ
uqj37JsJ7eM3aA63hm5zjSiiLVh/9UfdBxo6fP9JctMkc9YeolCggp+ds9fxMNwfN4+1Zh6ACE8C
RsE0QUQiiRF5+tMy/9tF4kLPh3r65LHUZG3JBr2lNRAwAqPNRAGqFoUiXauP4Xg7+Aa7iCnyEjm3
k2OyDZ2Uk8wEBg/6tjTrMKmPhohe5Kza0TFzH1EGHKkXa8H4EO1Z9s8rllqPWw6m/KlILI4Ti6oB
ILD5t78KEmIYInYqHgB1L/qvi6bjdAXCLEOy6t1ZbdZ0oXiYO+N56Zyj5TRTLlR0nvs9QPBsGUYJ
vzRBDnVUF2FgZ6UiEEOHOMqyxDrWmBg8B9ckK11dx84IN+xdkVw1QVIJMQckMS5A9KMvZ3f4Y2Dd
kRWpzINAutL/HolXsNlfcI6K+XjK5VfYAXrrRTjrPqDXcXK3c5lFPqOMMfqjveEIhee0KSbzUAi+
q4BPk5FQJfIBqEv6+G9JMTXRaliZPN3qN78KyHbUYZ6Mhr6tgw6MzPCwNvv/Z10gdwrLx91QnD8w
R6aSfVPwy52QU7GF8oyoKq432YVQlzgjHK3SgwiH7CR/oEqg6jfzT5KfBetFhjeWEq8WT/QzXUs7
KQaYCGra1kITzjrTmCBE+t/pfmJejee5Bbcqg680qJ195+1aUWrplsFpDN6P85GHstnOwyVEH3hK
ljGIc6RRPN4M3WiUI36a7KUD98PpO9qsKQc/9vQ1e0DLhgrHz0CZ9z/pw9uv2J4NCVaXrRxo26Fb
m1EZEj42GMZf1jQuUuhiBkp8oCBpV8mWMPEzegvV7TOI1PU2faFbSXPgHyyNJSIXC4ODx2JAB4dy
AhnO7FQZjQJCusmUIjYD63k47/rt79AcXyXmDNAi/HpxWcbHHhoC/rjF+JVSXB0sipS6MO8CV3OU
37OCLI9/aAaURghJtU5UqcgUxbJavIe5xo0rVETf3wOI94h5eHoDUh/Zticmls1+b4aXIR8vlSgM
Pnj0rvNorPDPCZ0kP2f/dmwhNN4vLG98RwXoeVgZl5BhbJi7b2h4PLyf5kk9IjaOAEemQfFpn1Rp
4Bo/3CD6YW8irzwDbPSiOf5RXjY9sno/OzXGYryh1VQKHlcTmxcR6bhaTDwwizE3SpypkSaV6J6p
B72bdK5fPO+w+jTsszqPWl1pNp+0NJc0NwXVr9bwln41RXv7QO7LHhcK/BV0iJUFJRh8d3DFxjwT
fnG8CHvKuCxFJ7HseewIHpqJLg9Oe/SDRZ0aGzYV97lywr/LZ0u0XLewoH8hsI8a0hPc9avq0+mC
1Z1UMwStOPxlH0SRU/YGEFoy5hDwXjUM9P4RIoCgcSLM2gnvdnOqKnOxanvziOonEZfJK2dPvcZq
eUQV1ERbVO6OzStPjMAG8/H/ttZ9C5sOLEyZf6PsEemgkQaUoKW9/V59W0nIGpoeEs/GEYuExEyI
43xDbrKnORaZBidHXMgXbIdkIEf1nogIya1hoJLH3ib8joiEkphNZkgZrjTBRTFf5nSGxGvr9cys
bL43tDNg0KrYJUdtQ09qv+19pUr8X9zEfPeTbSwJwPlBPm1vcCXg2B18Z6n6mmIVo0pNHhonon++
ekCy1yPE5cUVVqhcSCPYDAELZfFN/aJz92HgyhGQEFBznSg1VgGtgnJFvJP8nTZePrTF7Y77bjmd
b9hV1S3/RK0YsB5tTZV11W5jphA1mGDDwZBPqRufxN8mTxyltBbfYqwakwj5o32iP0+jGCEOkAAk
Mehgc0HltTZs9OzS6I9lmAipWYQ8LFq/cKmm5k7ddM/WEnHNLy0UmSnm/ZK3D/rb7G2NJfYIYNFY
Hwa9NANjjjT/cnn5MhbWUFfIursG+Uw+QV6aAhS3PycVMem2vGNbCtTPSOyJ1996JdFNvdm0rDaX
d9qe591IfRoNDYogj+Ct/KJldPJ6v5+3Wv7pX19kKi1yeLf2uKbIqPPlDuIQsK5GuX+lIfZXBbDb
FbjwUa/ovOSuzsLrPqgQWHOMuOfXLID1SEpG4FzJMFochcWUwNZ2nCWucxRapGCGb5HsvwEcITL2
3OLeSP3tV9Hgxkvj3k4OrBHI0sMmSlzK+euhv/8cVZrDRJ2xG8vhCX8WlxsU9cRdCYzT0kVBxtBA
VqgTJNeipPrxtakn+Z35Jmpl44t4cgjWLZ6L5q1V5SitNvSaFrYHhaXD0q8swhvR+S9FVUl6HMVv
7+JH8OEStdpMuN66i6bThVpRDQG3Rcvo9bseW7nYQTArVvTGcjzU2RKEYtaT9cUks1e6U3SVToac
k65hgyX3NSoZkGkN7Xmf3/kApTbnXglTl2Wl5WnkcvmSRjr0QS3p3TgyxE+Ag0qD+6EmHVHgBL4I
B9rlC6sQB2PCW6D9sKH/rhWX+bjaODKdSzW0jDtatDOEstBPBAORABowjBqGGLVwOydX/Eme83dY
PDmtWitwNtGMxaNW3zZ/ka6w3vUPAMeC6/p+KyOyt9i4XezRdt4TWXyLuzGqumeVgla0UCTjqJZt
dqOw32mavDRSAuQl4wQiUW8JZMrp16kAFrD7QgShrmuXLljOZbPczz1aKZAfNzNqcL8jwAmQ4UuG
2hjH0a14RQ9E3jXrZ+fA3hkQfll+ikjd01M3db7I7nCtL5xBsJmKH5NJjytyI1ufk+GhIi20g3EW
zsC0o11m1v/xGs4pSCL96pQaVHPBOL2/qdu6qMnxsKWvFPlOdlTJBFk1g/9xUs7iSHEP5WmqDGKO
veuPy/tDnBDwOffhLKvvB1Vs/yb3VQZYB6pH0ekdFV/Kd+idTh7LLiieuzDRUnouS1CbBG7mWkzt
taFjGzCRft/7/d7LmCTjKKeQKvgKp2ii6YByVkgTIkaJvQC6dnJXJTSV4K3MXIEhMWM/ga5aSAA6
2uVlhoQzcIbuX7EWkFSPmGY2vLp5GdE+UYVI7l2cSPIg14fl4L9HKJEwA2qBsgvwqCZsFSzWeJ44
qkDhRbRjB+RHExvnYZmMz2Z+fzkX3Zmg+QbV/juFSI5ltzdd8V+62/iwk8erBIkFRzFVPLSVphpO
vdT2FGmlmDzyeqW0zHdCmaOnWMiLJ589Ic+ULab57Zh4Q1agYQQJfEpuztDbCJtslt5tANk0Ora9
HyDPjIF68zvshioE53WSuvftMLVzps4yIm9YKG+ubzl/u8nD2bSLH3lTXjtwDr+VrbT5YOuqVa3Q
TkYtlVt5a0ZrMV7LYxZMuPxG9mc4CikyYJbo3j33y3NV+bZbmNOs2eEACYooRHYWgmFFMmG3Earx
6u5BWFdXw+xU4d5hNO9ySrPCHt4t/sq8vSuwRCpw8MLwXlUk05bFGJ2KmZukoChpKi+tUKVD2BtR
DKOif2MWfHqQV4y8bZJEF5oSBiWDAVI9yLP8gQN3HtHYf/Bf0bpjCYnOB17mxUVd07iwX5bgy2Kh
s6mXNI8D+hKF0TAYsUxFBFAgSa9j94vgjKSTYYrm1G9efjMt+fY+vHwJh6jO1hfe5J2UtCoKrLpf
DJvzUhZ2+82HXgYLz0Z30Gd28d/tLri30wo/gNplF1VVLGFXDCTykqV9mJFwdStJo5SdefZ0Vq3d
MgmJHfvppEzEbBjMIkh+LqIVNDe+s9reQ4OhpDcgJga8fw7/9a0RbH703YfA0Vy4z9GRkx3Vu0+u
9Mky0CwuI8HPYuy+S2xS3EmrufLHxE2eAqXeosxLcgwJz3QyUE+RMWoXQ1v/3ZxwrU7ypqQQcr+3
HsxZS3axzWJs1ufKwNkWPphJ0Di1LnZ+jnChx/FEZ6inO2cHA8E7OHMl3cDAbKglM/5pAsg3tN7H
apuO9ZG+pkPBnpiCvM8rezCuXb2hz9c1dUgF7QzVZptGRl9ECjl/hJlB+sejoqhOfdmb93HybB5U
Vjje3ZdldVebqYapzq5iRAdkCpWQelEJWGzB7ie5exaSr/XjXUXAJ9Bd0/3oBV1Gehr2jAIpDDfZ
GmUKW7C4+yme7vedJqwMx6o4fgBjRz5qLvUDhNHhPyRMRyj7syuwJa7MwIjCiq/Hb4BgKYJMS2s0
3unQXq0bgFcwOM6nWrbgj7N23Vh28b3lzGUGchh1dQhfe8RDBwyTcBlxKcmaFwY251KHGWlpeYi0
yFl7Jw72A2RcvePqyaj1EjTKCmdmkgvaxoaxDMmYEz7AAvtS4Ycj7Vm1htl1BPvgA8//Qo1CCKRj
Fe5U6iJzB8bk/jIJuvuuUwanhzDVPXcw795C91BVadiupRAhITZt7UFB5gR5qxOnI6H7oZUdUgZ6
ZrYdyjRrEyKM+gkSBZWbbbQ+r5pNXQa1ct2PWfihMZ1SbDOzUSo+IVDJZclm556fKl7aqHjsYHzf
f8ecfUUChaZxlbRwYqJqPBO3qi5Okudlsf5eNK8ZVcsRQmWITeCirLZP5G2r3LmCAbKg1QMdRPEX
4/BGuJ82nfOLFmsEsZyMwxRyHEFjRsNKNhBAdw6brLe1WS7AbVIK6zF9FVXNZJViSsy8xzYQFXvH
DFEddDgwd7hzCl6HyXOtUwdzSDdHDyf80Olja8oILxWgCc3P/fKmD6B3KXD8ReccwnGn2mOvbtdi
Fuo8LJakpn+dWkdt/wXCSSO97xlZV5atJgu0t90r9jCLUNnN1Ko6OpDHZWHUIgxZNIYx2Zzx+IzK
s30EN7I/GO7TYba0bd6CYJBssuDHo64VqBUEQhOhvwgZrjAntrwEDIhkdvBoUMFbUrIE+sHBMBuo
WwTPXucQdkaXAZh5PYoAvVwH7MLn9FpyWlQBGscuLliwxi+rfYew/X3h/rzwUW/uxhbaaGF4m0KZ
owpUQxYRM6gisOUtB8uWd52Ipls9LK4zwpYLAMFmgwZX8ai0oOKiNjSdBb2rYASZuWG3ugqsCiYh
fCM20G8lenGGfm7Ym+lp6JJOYPVS/exCVE60yAxbwb8MQsNTuwpZ/sCO4UVtrCbQ+Eo8zKxsW7hH
wXpAPDSN1zYfc24CxOD1VNYbuF93W+Lmk/P4/ujqrejkwmomGZdUh0wIZb2mjCct7QsYuPKwY+BN
hvhxta4ya6l/2tepshnXu/SL91FGIbPef7m1vQUSn3KSRAmeuhu6inwgd2DTnE/PUBVBdIJkKD5a
Ta8ocsPCUP6iP41D0NltkzKIQXSG9zXde0/4vwyy68kNKyLGNZm/bwIFdQNTdOrRJ1ZZJ5F+K2oZ
ea+WaBcVleFNiQIdmrWVrI7VvPmT7FUwHp33B4cNigSGw63Q2mIQ1RtuNI37PInBCwcJkxt1TFlh
RwpPRXio1an7F0EXXDHlFPPxci+L8UnYx8DDA0j5sOWF0CSx6osXlvkAty+/GS3W+NOrkPb48jOb
oPx8dQGCSETHxDSMymfDYygzC3EGHnJDaD+UclGYd17N4vaagaghoptbBmyYvQ3DwAQYQ06Myx+4
ubqASMlR7ysrmpJhHUXBqSaxuLnbXDVl6tU5a/McMtTKnAv6m+EbGtrT+XC51g2ix6tpXI5pt4/O
LknfheP3o21vz6IFVGbyxmaBejcACN9YkEGqvus0XIDnCXIwjHs2FvpmYR95SxbV8GqdYYYdmuxi
ACCzcUeRtjUcs4NBFvFmAJqqIGhrNreae4lCvNMI8Yp8AzbYWsCOwGWLQPHf+dvNsGVkpPBbWV6l
fRVBJSXNtmS/TLETv6PT2WMaeCSxUjytDAIA+HLjbme4sLqFFGxlukrZz9Engq4hsOHp+x7W+x+4
kRiWPmm2dAlp2/7wvvo93GRUxb9erT01ZvFs950q2mmMPJQU+GZNm+ekOhXkGuEX7A4rvIkv/OJr
QzUK+X4zi0LH+G6C+D5ANHsFj/ibaavcy8ti6Z4ZiZSGBKOthYi/yZzvaHd6SJ3izgTnC1N+8TN7
iOqUSPpX4ApOtAq/KXF6WudIchI8LUM/RbR5KFhSNzs8BDZVpMR3N1+yXsjsHk6WXGsD43wO0Z60
2q2aU41tM9jmNZyCb1XVbfWu3CJgn8uSKhSuIhd+l11dxZ2ZG5JYMmYuEaThjNbtP/t6mM2nI93f
JNorf6j1umlXq3n2DevYFBZcxf+nWpJG3T7GfLBwM0FBZ0+TabgueaKT56rOGqQ0Vs3SAFRYIu4X
caEgy2oopt9cM3A5ckvxnKiscjYuJuC0ERxCODVmBOuXKZMI9SVV5zgcKK1C+8I7P1xQGbkKwH8v
it/u+7xSRMjsIdY/hS61dtKmHG7HAN3vzwA4/bpc/ZNoSimSk4j1Ul3rpM2gEfUGmPojis0eo/7X
2F0+asKqUdq29tHYWbYJmVY7Z0mxg0WtArzyj5jaKwqMAuMsQ1FE1RM/Bb3BwsvYGvzQXtnNJ1VB
Puy6XhHzwxuaRRWKY2UnoZ8FohhtP1P2/9KEFf221tdVEjkRIlgLr4zKBeOCx/ezHwco/P/BXytV
QPUnRSKFxeJZmmHJB1tJBrF1xStSfEfcYMfuKMIBr7DNPlo3xCl+ot833DJEqDGpKV5vDizCOUhC
a9Cvs+HfnGNA1Rg2XvXVj88EUjoXCpL0cNjWJmqadI2e5Kj4Ak38n1px+f5f5nSIgRReK3G26exL
eQrU6NzdiI1lFkvSOgVq/TztxBZsosLHwziRXkeBnRH9x6Oq/EJDlHPjBM94MnbihR651JHeT9Fn
k6xxiXad62J1qU7eO/dQ7X2+VO2K+o+kUzi0edtuOrI6bg+2A7bLVlpFWZbYph/RHe1btS6QfdGS
Il4avKpFQfD4xTaM4E3qoOruwkh6gjFkyS/OqW9DU+wjC94hoX3NGDPE/e5SQx8O1iSi7bWxBbDJ
01s1prcitIoaEl99zLwQDVvC2tAbRcWQagCkNCkLoJAZ633QCxdH4MuvHYTh1Jz66/byCFKLW+bx
h7efAtrwSdglIGAjH1UjM6u5BzlqTqFIMgAt0poaBE1fjlU3j8VqboADgiYvEUZhBadNgR7bcVpW
vS5LooW+zrtOKzkIVDd1oY3in3po/8Xpkdx9jG4OBSoPtMg6MaOzabMR8wpfTAxszOgVn7izDFch
tQLr1Uyv1zor24DzrOwc9lwjwOKb5juMYQmxKrtxzPLRv5T0N/THhNcABfIB88ZmSmKeaL2tgrO2
KE7LMCfU9esQ8jzIN+WgEb0EaRJDkv/EMqz1/qINMNYOqXDQmsE/AhQ7FMDnFypkhnbAY2eXEVNJ
smW3zxnvMK6tr2eIKBa6vQepilPmMj5BT1mds57B3SwaUPtgB6UL0MqTYrkuNn1NiGKaQPUQvVbV
BUH16ZVznmEAotZ9ArzSVKVn0yhby67nLRdjPbqdIUDMhVbA3fNq7AjFxxmp9JRE8MFC5eGSyFW/
Ye5CxZsY8huqLR51MFF4zjffspiX10b0ihguyv5NU5H2qAoYGBusiVXtRhcItF+Hpzn9F6sJJ5fV
g/5oDTnLVthY9s8hGaDsVBvqSpnfwF8XuSD5HfeelX0KyOr+/jbFnM6FTvrH5OZrkAoL5gS4zdeq
jdreXfdm4mRCCyQlKKe0rc1PKYktXHcksj8sgfYveKjbEL2ktEmk06I1ubNVV612j9gRnYGFjWNG
rLQNoezO3291KR1FzojqO62TpsTLogAHdvSUsnJ+6C+SNskEbOQvqg3DuHJ7ZCEumJHFWN6U0t5L
+0Xkq39A5v8bY9mdlS/gZoRpOh6CDzqoKKE3dT5y2uyzkeQHcgoWvm/7q9Pav6DKnBT7qd0h+WJd
VIB+mt/Ty9Y6Y4wEdHUW26t9GCAzmwGP6rpDZeXAufBcodTPowyAeOtsrAIKooGBoaW/EOe5d6cb
JnCrw1cLtLWKRf/aWTa8G/FiLURcSXOKZAVH1h6ca/o7PZ7asojTveo6KA8nsLwMc6ufkaG83pd8
t8EcGND6dUiDiCGZAtBSzonw5qJoPg1tqAUN3XnClIhQu7fVxW/JkVEIuiyiSOIjY1tMfZue5NXT
3jOJT10uopzqPNoUCm+LWc6YNVlsU9YvNZhla12DurjGP/u4Oj54AWKojdI1M59LLN7C3Nqu6IqB
tVrYgN6/sVzo3ZXtI9F8wTm1mBxJE+40vew/NyC/AH5SbyBpT7cqyV+FZG0vm8twVL43HbQsf31n
cexjDoZB3MSHdMgx6W9hNEEDQnHwZfEKKuD0Aj4VFFAYEiySCBqkEV9w+/btpZCVldPr3PFamVU8
Mcwb+eYJaam6h/lrtRWvrOmOxjfhXhaSxmzAKrdwx0bGo9/E9z/gtyThXHlSvcaKJcsH4aRXfAXv
ldXrTCDLxckNFaLrdy1CHyFcfSYHw0+871DG02vdmBX53Nn5eAelghCaHZ4LdLqpRnOCX/UEliZi
WHBH+bPpCa4MRqI8xi3R7St3p/IikksnhQhSO3EvYacahMnTkP9dFsb4FwbDMuj7nm1tRqVRr0vq
aJAglshXmCcpmzTWMWDs/JgnDY7+EyJyT7Sz/cEVddbRO0v5jIW4sNzTeNg/6fTq3569azdkuFXv
hbtGcDc8F6lssWaoGCVsPHptEEBEbDJu2ChbBd43GBfUbiLhJBqcwPEGEGDVlJ/RNg9m4Ijv26+2
RoTi2WRJXJafl+ffAD2bU+vJkpLR35zgSibC3F1XKlLEZIFzbpKIfkq5DHj1iH8dH4TkfYW1WIrM
xEkQRaQ7gHqH5FeKogDgH9ujM1A/mk8aAYZhXLCEtj+8RdOn00ThtRCACziEF1R6VRBiM2jB91Ew
XrMqLKJcQL171x+R397ZMyYvsa3l9eXOfwTMTnPGa256rKgA3OgZVngeWR/k7oikiniarA33isXG
APRZwa7+YkCSVNhKrw79e0SklOwGhUv1O5ardOllSk8hKBFaUR5NcIZDPB6kXFyEqQWY5M+DFO3z
V3SybXoD2CIXak0tjdvKXtCHB9WvgohBZ2fcmGDINIYHMpABkdCz3+iK/j+OSvsz3GYEoG92EQDO
PKfkus/RIPcmb9nj3DyYWxNcFUbgGjqeFgomJ5twbPBIFniH4LlpAVVGUUx9lht4A6sqNhfSm2r8
P9lvjVrU+zd2OqlApfTVvM/QHLbDmlk1jpCDhqBFutuZ83b97EzYW/tFSoPl/FS/7g0lWWV9YBxC
zBf06vZtcKdTHHdOzpA/UVcHD3Wa4PLzKTP+/Kby+0s6qAc8gKQxOIRsP1zJrjQh1Tw3aF/QLxYF
mEvXfyVWmIm+l9yNrBEsJhb2v+/XiwHCaSWmkslqXgnChx5iFDIX3KuskWqAN1kk8zmQH2eArGRH
3mWJX3mYtReUlWvcxRfhdJq9NnJQkYyEIH8TGAF63MH0jE/YXt68nE69kMX6sNKKGqM6qio+y3CS
Xl7dbhahr+KBu/m5X5/yNP1mjP8IWSemB5RQBQDcrUHtcga25d1u2eH+THuroNFD4LCsskaBjLv4
ANRm1yzwg6cOdUyFCO9EaHl6jbqk01THzi2FWai3V37nACw91Rktnt5JXgWjQdUv9jnIDsS2f6xy
ZSXceEmfOg1mKBTxAryI4UeA0qQEB3kTpcTZbImNQ1UaNzQDbQfQJaD3SEtENXhOA5tJN+LqwYYq
s0ZdxGvpflJEGtdq5afUyP/KhohAGpjVhafhWpI7AvcqEaTxHzgdVRas3oMkF5GXWolTZ2n49oQF
OJSH0OJafIQWiYrtrYjfxbz4AGJJNtPQL0vyOj+ooW8sR25DkrD7HShzozLN5UFHCbzHrciPW1tS
mRT33f/W+1jsqK6VHZftgi41a1TPbH8lC6XZtDXd4Urzz0xtUN0tUiHGsjuqADn3Qx5Ci6x7CWJG
ch1TKsvcksJTWAYTGCjirTG+/QhKNfef84pgN4xqxGXBC/+16sntIiWgM/sVd4evpwpmpWKlQVKt
UYUmfJ7yGmWqLyX8iM7jsmQmcFp+N8fjAImJOsZMLfwV8ufVkhkuj1fni9L75mURCvqrFYjQuhtp
1p2AM4dOwpRSHMlnVcNtsKTgSyR3OcyMswJjV487tjG5lERuHkLv1DtL/h3Tuo6nrLvbbjjhedDz
n/nLR8akhn29/Qip9bda5kAH10rk0pKkRfsft+FJhVZLk37w1+f52WnPC+Klg+T5RDnD+eQWPCgH
k5RmXoysYEaQF702rgXv58E3O58jCegah6kuS/kBIF4ddwVbKU7lLEgrk2yiTe5jsfUk4qXot4hB
bDBFErnVttw85xNmBkYnQbo3eS9cd2R8BxYHr9LRR5y6hUadHKOIhdfG9PXcNS/XlFuqsve+awtf
msBTamGj+QPV3FIUYtoLSTXSHRF6nILCfPWGOP29cT/C+Os6m9+RFQA0oVAnZUuQIN6wvWohVdCr
Wtuq4z3uKmzIflrodK6ytXsck/Z69yA16+2hIkEm11uVRZVYz9WbnWIQBZaRfx73FJYLzwjK8w8t
TUgm9QJqxRvCEpsq+zmw0vn4G53itO2xcda9SuslLRPd4MjMgZyIzsPL0rSbdhR2V3Tl16TZOlkZ
KzSl1DO8KEJRM94AjIg8AyOd2vCg76PWMHPsBgo7OfvCIUJGNHAN0WZXo4x5x0eBWsHaQHdQtamN
TWblbQ14Ci1WcT6lg1wLq+B343K2KT8yjI1ydRaOjGOFg48k13tOssrNHwKzc5QpVFL64dL8ZnnR
xyn0WG0K5CYFkCaH4NNsHxcJT3D7SU9BkY7rg9lJ8nhWAmywqfnl3Wdy0Ynk0zsoBiES3aRPg/CI
YMRrZ02Qtedo34MjBrFzUFVYjBURlpVsDJ/GWi1XEWOjN1teUtvl4fXrDhljxjVrXmjeibVmHXV3
QUUDLf7oNVnfdDbsaCK9tqszRCRfgmgtFTYmxHejjkua4UpKX+qiToNoxg5HlFuHOeJ12aTPcoEB
5OooM1fmoTFbIEz6Gv6YMpDhEclZHUVAKBHEx5kF4SLdK4weO730SyMru5mW9K/VFNOMtLjp04VH
MK5nkDlv/gvKMSoyDRiAi82WwN1nAVJvNxE1TsI5fCjIKCTynGfAl35YlmgzrrvPCLqZbAOVDm/U
HjqNaIG7CFi01jamkkZDGHbv4hmAzkf2Y7uVYqfksc9sb1E4LtiH9xpDFopmDs0PIzPjAn7ATPET
R8mywGFDkxV+yuxOZNpRh0ES51SiAmRxWWGaWG0oJ/YJ+Z3lcuFkrzBs2J+vzBdoqukKC6jVYKX5
jF2EZKiu7LdvKuApV8AcNgjKig+DxafFHX09C5ejh6/aU7bB6v3m5Gm924ayYOzWkxyHiTQfbN6/
/j0sC9efY4+bamW5iE6++BgvYjWikNp106P8gkSLlkEJ6yxiVATP/miv7UbvUshk3WhbeWUzclc8
5K71NnFokOK7/yS5I4CxtwXf4jXFCYA3TheOGgObPyHwDuJauCpQfb1yyhiOt05ozJlp47cPOBE+
ZrBp/7i3zjHkeASJiKfi0XXqDbLSZnT2a9cHHweQA0B+YiwUOjMlTjuoOMjJ5TwTDB7cw11kWBZl
8z349HKqFTPOLiiISlo9BbHa+IFyfGAbJSAdxoPGSayKYpSENwYhrnUfRonJfoFX0uwm1StrwaTx
reACajegQzBGNlPxjA9oA1ztJtS4eTee/LPfIu7Xx6Kxs+iJt4QY68mRzKVyYZTlml63OTeDF+wE
cuATeAx2b7/8XqoMCxsBIMgK1Pl/Dw61kRVk/LWHC60JFApvgcxsby4prgsZFe0aoMc4v3WWX4Cy
4KSdvDX81xeyuLGEPSzM8FvQViDKbc3vvTImIubwHI4wwjZS/KjtBjE0iHI1c4IozgEZTkL6bDn2
WfRlp+lXZxAjgS8j6RuRr4af0tCzkptcnBUsueaokqQm1VKWxxlEPNTtiYMkz7JluJV3S0eEZ/DQ
cHMZ/M6h+FstJLf2dsGr68V8XBJ0R3dNFaqnXpRVQbrBJc/5uO90iXKXb4Vym+xYieaQBYk46fzO
6TIGknmtrrgg8ksmrjOfQoezUPgP+ok4BaVon8zFE22KfiAtpv/w+qjNZI4cSH4SW2DK35DIekWV
6iUgkdYriPkfrvMQAUBoR5w0E3Crd5Re46ZLYbjxuzoBxdbd7WrZp1oTFFZuDngS7lUL6k+LOdeH
wq2aovl50DdrSKAZmLdrQ5VLNEevHhvUWgsk8j85Z6StizP4PUUNKrElYF2+2VBzj6qROiPYSiID
RkoR+zls5EYKiquOVoP07d9z1eHEyUYQaClMhFhSzYMmRQWLJPq/9UhHIrlPHIdlkcBXCGwi26/y
RZu0+m/cy4k44DnqoGCoCsiWs+rXWJIdVDfG+G3aEblalbMqaqT5tuVl+U99U6gEbpcZ8OG/m3eu
1CJxUV23NA/WBWfYlfEKUn83oJrLbcXBnF4BC5pc4VKk5BVIY4mtgBT7b1M3ZK9L8EF6bmu0e6Jh
KCheL6O48xvShU+ppt5Src+DHcrx0rkY6iHunrZUWss37Vh8Co8GxaXxEfJaRlqSKl+KXViDoyut
iUmdvVudkq0ZW4urnCfwDD0mysRFoQmkaO1aayAww5DzOWo0GH0V4Zo3E8sUXqMNWJttsmN7etDe
K0w4+JwZuYJ/W5/btD/cidQP7Hfk5zpvotEJOCWk4m83pWIt25KlBhiwF2LAhlgMT7HbvDEYkrgn
p+yma3tpfwaAJae6o0IKM6VZHbaLlvX9wtxEOHMhiSoHcDrfPp04b5Cor7zALDFkDJklfbKVcmNW
hAXnyR2CSZBF1Bq39e8NjYk0/CiRC4k1jPqruO6ColXnBsEWOiA6+a6RAD35WXFJN0hUZYruNq/I
+OwZGZKalolFUaY+dTzo48+y6dSVz0rxPifJIGK2XJgMaxffrz6Vq2XQ4CWU5Gce+czdhWswC6ah
pMJDoPnyQAYswaF9+WOtayxwcIX4bp1afZb2qlIo+9A+LkZ+FJ8BaiW+7ZhruJNlNu7Ha2d8Zmha
EGM1zNC1TvLbhFCjrLGY8uIhgP8BVKxhhibaJ+RIpCn8wNAL0ctyMGwlvrQI9biFbPl/SJ4T9bi7
8P8A8RidYfsaN6Q4yA2lBwzeXG42TxugzIvy/GRe1cP6qV7JJCCZ9mXFZLEMxnAPUh8D+85taxrY
zWMF0s6VirCxeg1wA7UWroiE4PZeIzMLyKVUkfXx4EtHCgoQcJesqD5Ec4vsxKV/AEYj9lE8qUlP
GQI7dT71UvaZh4b2ddmbjRCoiKbw/VYMLSE5u421SDaiVDacwm1z/ryMCMkcDWfs5FjocPYuyVh3
dRS3DwOFgc7TCWVBDPbR4D+4PvXOfvdV+KQSBZNCOGtQMYpYcZaBEMBfp7js2aJpVmtpKtlu7m7d
K6dHUY4nOgHyaKwhq+TsgxFRoETMZOHKuwd++SWVpDySYaIEeUkgGH0fnL98ggKsHcUb1145nR0N
ftf/W5ul7y9q5mvyLOwfwnvZn+JjO1cNt57AGNjd785SAaT6D7PVNYM20j4xExg5QOeAS0fMx9fD
7AA07mV+RjUNNTj2uQvDQ6VvFsHgI6wNtCd/RrPIsGPlLANS9q6EldnoJHzQBtHDMJLWRoKUNZIt
D6Ym3A7HNR3n4SFNFOrLxT7niaADSqvWkjmvqd1GLb7zB3iZ3fxPIojFkp2zma3LSZHnpUefBiRx
sasR6gazc+qfRGK2FjgibYt/icKAtVfuT8e/PKKYsnkpan7ykfrG8/OCo0VSxProYT4ppK4n2lZQ
dUsG22dIXrPxdWMmAtkPQPYqwdVfuj2sLqIMbFBgGnvIbeb6aV3R0OeY6XhjQ/wJfQh6innRIXjn
ayUMW3555APNAst+zOvgQz6XJ5u9STa5d4p21yCAuzyAQKQ/3L0exrc7io00ACNj3tyvDiyYJvMU
lR2y+cyh71FejHgZ4Rn176uc4Mqr9Xi82X4/4GiQuRVOXwzlIdeG40iA0qv/GT/HIt9Iyelyyhmh
E3tNZeP2VS3oLXgVcB322N1Jx2SY2d3+DasoE3Ljjuy9ROxjx11EbMfDdJIky2wBDBVvcFFpaqvZ
iGf3e+YXKA33TpT7suUEDAc076CP6vuBXzd5+Pg8+DXQ71ALMltr9exlclX1C75kcYchBJOyLOMl
Ns3+qFdTZdmyiI5Dp1ZHt0W8hjISoWC2KldcvfAkGOr7BCLplVEVx588MPYw6jgxMtM33JVwuE3I
HD2aimFBq3uSNEwGIiQZI7q9X0kxcsfnGJJHZMOYO4t6Aw9BXTIWc9bGEB2vAMG02LCWGs0qdzC3
eBmAd7hZlaMkYSHzqqKCb4HoQRTwVFTFahBpN4KwJ1vHG9q48hpg0Ko5PQi3hvyztE7K2RB3GM3Z
/dAh13673PtOmNqkqDovKXiR4BAo3H+6nCBRYxhAkeaIBBYzti3mGaXTg4vpBGUhV03cYKI2uh5n
vgVAWjQMzd+HeyCChmT6+rRoGzsGSJeMK1P0Jzh/ii7uF3U/7xdHr9omy32JYVRplx4O9Ktluhyu
JpnyurfFKr4Ie6x+LUCI5e03VvPFThFy6eW35uKq529z7U0AYctUzq3i9cCsk9tCPjsY1NCt84AV
2d6Ntc3h0H8IdyRDfHavQ4tXyAzOKwA9KCYm6HMB0D6Q66kLsx3TvkfpqtplOftuEbtHiTJLAYp9
xUYYjCAh4e8RswTi0P+xw4XK0PUIk8CLSFqkd5ANpKoXrmbkHosTInnNhYyoRjG4rM0oEQxfC1tx
LOlnD+aoyoOzt/+NgSW07AjGIG3MfXtAkzLO5pjCXM9K6DQ1RAJvuxBSZEPpuBr3BlLl0urzOOYT
U5+WN0tQmRH5Kr1b31VAR0xoMH13NrsFc0kueEjMhCJFLrVaOTldfUt+HhbYf5R3eyxebGkiKTwU
JIuNIn/ftIsuPTTex2mWWqnejz9uqxY5IFcIFzr6KJm2v5ENxFls6ftNSea4UpHZ4m3wOGZDmmOY
b0Y1ZQ5B/dWKBFJD3WQdtnxwzoGuMySQeCXgiDJOtsrkRxA1KEGkbKwH6Mm4qig5WulprS/tLSs7
TDujbzKlz503Tz5OsX98nif2KNF+M3jEKV8lsBxHcHyW4+PAGjhYGOnBn5T8gbp2Z4VhMqxkUpyj
PDWgQc6eNGoBCYGLshkeqCJArU9HVnylsQ3o4/liX6tM/jAyzRwzE6/xoCM6EeGNmuhrSZb9G6hl
7dLJDNwQrBua7hGAZdnRnRGK50kUpGJ6cPVWrJJJ1wA+mlcjQCi5orBkEjbQZR1On4v62k8Wjx54
nx30P3iM2N/5vVvCOnfRCKwB7/dM9ZpTndD2kxgI4YEqvhOToAsg8cdpraACwt01PGIo5hh9KoeH
RQb1Iq2/eYXncVe0vQPqxQVsH+AzQq8+lVxjghI5evd7GARVPgiT2y7z7DrTgws7LksP8Bv4FKin
zeFHznhvx7g0uirJ8nOyK9lm8veM7d7a1+ip7el1GKTzpQ+PQbsJbsK+v/I8qidCxlrepKLh1myJ
/5fnj2PPtCW3gNdqfX1JTHVkbMJlQPM/jbfWymv/rP4Be8b8fF3Og9KLLnj2cqfK5c61CGNX9KM3
PVYsOsxI9Ly/hU3I0fI9g3iVBHZmnaNXrfRHJgihr/WJhUxe29ZCTLJlfIwAACZ/56/r2ZtC+iFh
KnD+SCwxsZcrOU6PNWOliBZtArQ49aIK8J+Vg4qO1F3gSlRHsomM0Y6ulgpBPKyLZBLkFuW1k8l+
EH89qMSM5uD5UR1yfn9aZLPteco7FCrtP747pZFGg35ROFeLoGAKmflp83/pzvRVc2cg8JpiJcuU
FoC1OiZOn25auW1UKtAaoum54/jjEghRIREXWW80AMmBAdGwE5KopwH2kFScr1g7+KLUZBZ0yP1f
Plac06NrySu7XRhZ2+udzr2F6iHv8t8U6cDGx+V92mG1w3XBL0NSPHDH88/BbPu8kWEi2VOmT1U0
P/pHH6IndcSHcSDL47mwM2CY/1zDp8FX03cTBJRDbnpc+uS3AqHRha0ZHze2riVN48VBSXdayyTX
k5UhAf00S3RnibA1qPO+0rDca1ttmyr0khSWitNZjeBrimLQiPdElPPdQuh7yicFU4ImolOaAgGA
7X9IxITuCI4Cvhx6kThZs7zHE/ujoGbjV2B1R/fegDNdnrU8s/rObuyEe98+btjgfqwp3iS7XnZu
QYvtGz1blAi6Aqikw8cLXuG4qyJZmfa8Y5ZHWKNAZXBIIx2GA0AVG5VaZnYFbNZYipG3JjgH8G5b
rcaQ3FWRkDnAH49ihSl1ZJOsjEcBGJ0YO5YO5G+jYjv9LG4XIFHr7ZtAPBOSfFE1wUb1XzUNSYqQ
3MFQDwnV/5RvA+wx6laBpmQkc/RMfhLKSpohmCP9/za5vKzDzz/h7PxUeJYQM/D0GDqP7xCmHX7n
Rgo9N7BRLoasjFh/LyQONUFplirt76QCrGmhdI9Es7ZjGSdDColspRwjwnAWtIuycmAaFhzA1yXl
SA24QERt7W4b+5UTvjb4q4gDh0F2H3gEmv0856DYKHGIt1oYG4IqzeDMSYUr6eNvTgSkYGXm1vrj
uzu9Se/2W7pc9v1BbKGALyyEKfwQayUZCMhzUzeKu38GL5E4SlX6xezllsBwDIBosGtR098VEr6a
ofpylyy6qMmujjkGMkloV3TD2gbkyNAPqWViQHcNWz3knCYdsLfMmtGJwtLUOaAARrzwDUREFjVm
LTgmOkE/72p5EtY1mwZw3u0AhSaXdz2DxoCo9T/sNOC4s6StEGNoHUc+j9JPpvCs6BmqC5QyAB6m
zrFh772xu6N6r4SGqE+DuNhYpzWLv8wojP9QZ3R6mldyrWaPpNeh0rmTC89e31Aw6wnqosbyDQBv
dmedvkwasZzLqEVCLw7oz8169m8tNzHZwcCDzy605Qc1XcljX18J6zET3zrdyFAmX/G+IfbjDo/6
i1VL6qs7xgsczXrrDqLEgmkLNJ0tFjXX5xHAezMjHPRnyRxPjYvQAFWEb5AC62EWq2GwwZ0DHr0y
7bAUEe7ppg6z996Kd9AgUcBZdAo8Is9LH39kCHDBKmROPJZbTyDtC573Uom1NSJZIhh6dUazEJ5A
itTwJsp3q41yNkEnCz2eB6z2Hw8W5I1ddAcnjbT0eZKUzmdxrMnYjdZmLg5tJGTtjqZcN2T8E4k2
B4uhTbH5ouVcj/I8JXaT4I2S4qpQgylSdpc/3W88Rxadi9f9+u8kIrcN1vEu1EQVtw3wnmv/MNe7
RcEOQp1Ig8jYwAGxchtePN23E2pzIBltkwm/6SFhWlHyjM/vey4y1G3qvOG1uCGpC/wso9kEH3h4
KCjQ9Au/RDzkdsSC4Wd8ghfz1qp8Dy/4Fz7aKBVwR5bOXTkjWRh0zc3qIwfILahORP1cQxUlrMG6
nHKJbJe+7nf1b0OPL7HLOvANC3FeH4BaL82s2kgFAuybqy+4QZynRCcjuQWAejfqtW+UBmhF/vol
fB2V/I3+RTTZ+rIDHvbi6/pyi7rOQZ2D7IVN93VdDED/7r5BP2Py06xw3zFkCcJWcen9xg6IkrQo
AvcEVy7PUfhsCmpZ/V7AMIR0ubAZ+sAHLuSOdcvpMF5yV846oHEHdyxim5oUwqI4+UkqbZzuhGTy
kkxPLLj5VqaypREX1uHqXa6K75TIYeeAUuvAGlXDQsMt0jO0Tn/h3v9zFMamdGqldfzspYvDTRvV
OmAsUEmlzWag4dHnEgZnl+EyETYF8IvjrtumBD1gVpHDly5aOQZVaQ62OYyMFjoZY/ic1r+a9RAK
g0zNnZEthJaMPJRKGPIBG7kbqblxvl+0Uq/Trhm7BWSrcS3QgG4ZxyBDkDPS0PoGrdlDvjwcmsdk
9kiLxgLOjnNuCopGTbemcaD18m6FZLZZHP0J59STuTxhX7FOxH9W+Uv0s59SbvQnyVp2Xif3elz7
LWvCAMUaUBBoCEDhLcDVvizQAtX7guPtoYkZIShFn7I7k9LK5sRood3f20N+taHONOx5wnpk7YZF
l1QNxXv4ZxinEWOxgLJdgL0FUGWDdzmWKZUpdy6de7ZNJxK0dXc5mwqsUyBtiKf8QciBoWfTZ0KF
kvR47j6sBItjdm8lCgwvDQDJRI7cpNQIO14tP6FXRLT7Ip6m499371mOOCI8G+GYhzYy76rdT4e4
maWAZ0/bIj/ftp9Oq70qNKCvLKCriMb9GhSHscfFb9BHY6xJqlDq1N+gnSBPuqNrrKRLpV4qzk3m
FM3H1tP1qunodDKGcIjMbOJztP8+pbypR0qbI1YueUpQ5EBhywzWyGuuPoNmRARXxcyynKIg244F
lZ0ATPmKWftV5nslPCfhCZ8nApZs8z7daD7L4cslrPxfO4ECPcSHz+ad8UZFlYNUO7iXIX6QxN50
7mTw/ruww+IOfy/0KzWjVs9BCnEiZVgCqbOAsHGf1/DZpGlrbr+/Y9IDyAQIpwvhO25bAtWdGS9u
gTcMHykVfMv0aOx1UY24aoG7wGUh2OBnQA3aExItGc0RZxU7CWfXxIiCLrZj4uDE3FWE8lTw0MCA
lBLGMe4B23CNBa3okhkJoqaHkmFziet3qORpBwNx3PaToB2nIjtsxP6hSlKXt/+bjRt6TipiNScW
SJ1T4xsc1TvXgrMyvju4iiS01F0vWBFSWoSv7g4T1qtD1QLE2J+lT7zKstfqueynLN6stHGDWTMZ
c1RbbLPOKEAG+9O2g3cyMntOKGn9QQgdI5kBeFQzPJBW662D55Nuh7o1Uz/8K1jbN+tNOb+h6CWS
XFPMAdZY2l/8J+gNXdwNiKi7z432t5cBovoIEsXUZWuPmNHJ7n2USdUZtANmKICpcDsiiTKG1Cnm
38TQfijYBO+cgflDkxoLTDpwB8b4YOHz4h+voKYCcvbxmJYqm1W6B4kwVPngXGtqd/Y3ltm91Nm1
rShqWkP0ozoGgK2Kjy/IMxNieULYqt5wrNGdfQSlB+5+SDSL/rhbWXD3xQPauVhkOsc967fhrbdI
gM06T+xZ0Nn05e645NXZnWjt1seWZ5hGfQzA9RdDfQRlsGXJlEMHb54qQWl8cJLRU/wS1MtklVfO
WV67GjicjBc4CxME0FSEUWaA8fMCdQLrS4FzdF9Hjj37EKY2Qhy0mM+nmK+RElxASG3pXcFtxbD4
a/vIoIWAouxAMGd0kZkP/tK0b5LWLXdgjWf/uPhxYvmcuhNkHuOCPboXEIcAY+SAZLJqYkdkqYiY
pG0uclr3lKAzGlsjPoor+TJSv/BqMBETtcLf5EeWCfD6dgAC+pUdT8dPcyjvU/3G7EASSE8McGFU
kjplNQOQ2Lw9jATdfJ/KNU7qP46Kk1DCBhXoUMucI126ufBA2lCpK2+V3JfXLweyquDJ52YnArEn
vs8SLF+iqMdenaRegJ+IIsaZuJR1kcBNKcpXvMGwZ/hXfkzC0x9+9z0IaiXkwsqv1KrGQEwn3Wyb
drswFgh9WJ96UY+dKRH+1611K858vtRQr+SjJrh4sFIbMDQEkY2cfoPTk78ie4NIFOcpzWlq60Ao
vWZblyIrm6Raas9K2uCNyZlCx/W4kFyfzAQAYvnDWymD1lsh1XUpdI64XFTA++9qP+EqLEhPGhhu
icOqvoYxwz0LBdL1AvQMFW/5Ub0jzxIDs6iNflQ8d4nTaDLFZhfmvCIMKaYNLmv2uZimGeLZYiz5
OD8fc/AiPwd/U+OZFE9CqIOJlgNMa7Fq79YMyTR+p4zgqU3IlWjh7pYefNTzeunJRkf9dLUBTonL
XkmCp1nn3Sm7mz7H8liyg2r7Etv4qu0S29K39CFwrTPNX+keNzef+IyG4c8svxFe7UtSlDCEig4g
ooFwDTMKdUeXVVySbcRHkjxzfGZ3tHAv9rbvzM4QwBIyU0Wd7tUxEgMIqBxBuhCVeTDhegYFXRcw
dET7DsXqJ9zysot1JKphyCeeNsuHyN9W6YBZN+PHlbueFy8dRhQUZowKGRVwWJoZ9pE9aKBmiuEr
kcNVhe27yrZIlZzpfRtLsO2l3s+thQpTbYbPz6uXmfSPa+iPTcB22RS1pLFmERzrbikm7bKu3z00
Q36Mt+R9BKIUOefe88vmEsIyzymX5OJUUNjV7MGSIlcTft5/i/R6TuENsNVz3pKaCQHZkcSvuhj2
2eOr5rY28gHtn3CSU7/kVfPPX8AuKjMEPNn7GkMd+/RL1DlXSnpd6up0QdS9Hn9hQRV8rMr/w5ov
4nksyYd4ARpM+6qEb1A4REA6blwMgAVhlbH2dURqXZ43pchAQpr37hKeP/BijLZDTUcHCMVRJy4C
phl7UKoNUKI5R2Whb1hTKo7GMeB/GR2bHf8i6h+aCitsGo2bgHMhtUwgLCiomIvMBjkFcIgkfID+
8wBQQ0KbPF5dfzky1o7Lc04z9agUi/Cf8+xPb7EEX/RvJlZcIoSF84G88OUa6SiZN84U73XfXg5k
m0Q3jOKkRovb65prcbKkWlvnzUXIdgWB4fqbPHQj2LBN3XmZzokwi7cD3qjK6OFue03v+rVvZF/a
ObQ8RwzHBLrIvvw+F/YXu9c3YVBTYy37PLqza5Ho+S7t/XYkCPmmjajwjw00SOx8rYt0AE3lelk+
b+XtsWeVEJ/8Igt1tdlKJCI7iVRQ1GAMQ0wnOIU6uLvHI6znYYBptqBRarqMh/Bgn3W34Dy/Ph3A
IjMO5LnRw2cJCaALG/PV8/xFbRPqRJvWqQFqzD53+AAOf8EpXkjN3SakHNl7xnMk/uZaYPHO8p1A
5LNb/wnIiCGZLsFDDMVfv/b0EQ8HmcKD4oE2dLfJOVfEE/8z7ffKJF8ftdIVQTK5Lw6Fq3iw4jKp
3w0h0dsRHERBG51fz0Nv3LrpnvrAiiOVGY/+SVfzPz4QckKraPnT8NWDTMgpydrmfFVkh1t+Bboo
VrGz/a8P4RBt1YIEP1XhLxiwUemxoUszfiYOO1ZGS25PciRm4fPsB4g8k0vicH234nWmY8ACwV5K
+uD30B9IVMrpw+Kw0XjwFaXCM8BuCdCO3Xps8s++dlGnihAzWicEX90RtTO7UERxSvEpO6lX84wh
Xzfur7S/7K3x+R3TFJLd+/4DTGN1T2Kwb+Lt6CasORFa4YprO5vkae++1enZODpFEyrxZ7dUvtRy
chemCtSipBqf4M/hDDeWFqOKFNadvMmXQ+lUb/mtrKNgAXgK4kZZMT9mALnRPyzysv29ZhXDPZVl
6XOHa0Ji8LiTv3OrGKQI15VlhYNFvrGyUqEXA1dbdGMtiSFD9vfWyx21uKySOR9dPziHtxOQM5um
2bsRs9ZNv5vqkwHh1XNB+nd1e0gb6o4caPoj8on8hWOu4YhQkAmEcwcIW3vOkAq7VBF2feOyb2Hl
ESbeIvoxmTHoKpZJ6e85LYZK3Ey3dUu4XbTkDRA+snb6HvgaBMywi2eglYC23U2cJ16aBotfsPCH
I1x/l1vb4z0BcCZms3vqQlZyjD7J89MGOaf1ax9giKnvVuDfl3ePeD00s5/T39KGisKHaRd1Ddos
g3QdVH4S1uW1HjQ1PG+4Wb4FXgvCfKJhVjg/HlLe9Kx3rlwZhqyw+DrVed3fhrGOfLJ7Ub73ZeoW
y1c3c17GknW8y+UCg9Zdg27qNdS1943FfoBQlr90jFsIOV9kN5DNtWhP8gEjAeEkNJy+7TNdAsvj
toWiTbMBpS6Mbezal55OD5NF+crZujcsualDq68tsXDx3P/XmrD2n4TV1U33IRLNZsArKZu4Iy3M
KXcdVGv2upcDVITdtNiTSdqH+cDEXyrZhUAaE4j1JeIx0LFjmMtOmuuXLWTZgSK0TNPtxeEDSJgs
y7zPp8aiAMzzMgXfZ9VCmyJnMnNA4MFO2ALB1XsBmskikcXdMyZDvRMOo9PuyI+IQBWPumIH9Ovf
1E1G+54Ll3MMF1xzHMB9uS8nW1VZt4KNRRQokK2S9+dW6XRHEdfSsTE5VPSEsvbHvp1TWWWeOCho
4VxY/ZVyC1gPBVSjddLF/bbivecSrSb1YH1ttWeF8kosyQPuIf2une4qUxTcFk46choetFbzGReg
Gs0ReWq+G9TsQM5rsRP2Os8n3hHKH+XZJvQi23s+s85jtWeBqNkpa2gkEwH4i5vF4LhsZ3J2inyy
R4esjd2mEHB8ARH5Ol+nPh3yv2wvaa1PKuIX0PWnsCJDTl3tYJriZRR4kWt7WmJQzW3xKJGuJRSQ
lHk+Ki4wt3Z4DrCCI/TBT4ac+9fuhKXC6Vd9XjyJBz+Ykw7/dtlPrj2WgU8LiaNo3IpUq7ga0Oel
3DOoNCPCc3ka6n+eoAYfXGNPkzNzFpYzuZ4PVb3ZF1sSzQIQoS/DebHMhpt1IDyIvng3kyE2xoJ3
pa5qLB7CsQrq1mEhWPaX+7YZlaiN9hme4CzJOG3WPgZdxXzjViavPWLQtWQ+QF3GjG5j2TYPkZ37
H1EPy9klAwsVA3/+eDvaGKa51hF3I900ww6tx/fN+km7Gut5JAULwk6zj7GtnNNH3RxJe0R7QISw
p/LenfAke60oqut0DMvkCAAtTwvl1isKQeQHjbRHdaFWKoNGTE0GDgphIuNfm0LgOIMhaWDmrOwe
hZkIXDdaj1fYlw5/xCJ+0WcL80p51VOFyT61QChDvzFbdbtbmz8OnVKKUv9weYoNVzOY52mWbYd2
UbcxwSXakcuyL3ApFtALOaOsvtOGSASFwQM/jWwCiW7rbxSRSJKfCNE8/mx8iaU6bYib9AMKxSXV
O2DiAAes7yLCLWbj2mIC4jZLOSlUytWynUm+2/GTAxFo1UPNtt7hCLZTwEyxC6IxhcizozVrQC3m
uzggsL1ZJJYxfiZsCbymk/NBUix+u2w3ZUl9uI1RWdStxGqs83BoSkoT8xWODx5oM+yMQGdHpPQg
697WRDfcCBvMnnpuA9k520H0SSdULyNLO+EZROxWwzzStzUTIxtnVJ92ICDgI0e57k7unJ6auX7r
r+1EV36f8S4283SashfP51uWITr6igMC3WxwNIFQARY7HF03xM73gwon5sszCp6GF/f7BSz2KXt+
3zJFkukTSWqpouTRPVBOXJziMKD0a9OqrRMyKYEQy0malICv/DbJZ1Z2chhfhkjqnDGRN6qLjS4s
2ogU1aoYuFmw8V2LKLiB1yTtLlISXIHO0rsv2zSkUHveq5uf+Jo1aQTQaHdePTNchRIc+Gz2fe/d
PWIMtsB31HccT6/7E8WU6/LLQqY5S9ZRNjFSXNy7B0+rmc3ifSSg2Zn3SbrsfSMPZg3kjfm7Ouet
bSguYtT3BbUxl5JpUu86/tOp/G7q0AblTUHGH/ZohOuqxFowuwWxu8oBMx382D+GRUbI/qUIfY7R
YY7WSMytarpBb4I+Dt/qziff+44eTQzKEJMYm2qFOa3MNwtovqxbrRWN1qVtmao3OXKLNIQOMrUK
GsAiEPZznNLuoTv4UYzwcLXl1RY6PL7BfTsmxuCvYZdoq2jmANO+p2LQn2b9FCX4ekne7noZ07Js
1/41jAeIV6DY0s2V9XWQvchOl+iCvRm+24z3Y03mHnzpmcKxkS4mQLLaUossquk5+E7UQZVzJpmb
iH0Hnfu1hhFpYCI74bpqg49HT175l0xk9EFWKr3cTvnFGRMzywtS/DszzgD9IEKfZhVVzJZcmLPl
xUXHvimJT/+FrG05hf1/mBDXQbHKR+3aPuc75sdfe4OhWzymaAV01fIRBV590g0MA1CBEJeoadF+
u6/eBmaw8P4/nQJCp0+6Tp1ER8rzF9YzL60vYWZrEz7wr1jitUzVrsfbEXMu4BGopjLBq0nLvQCM
Au925jn3OAlCp433ORcpqJRvp7/CgesRvog75hmxlAppZKgKEzExV9YigEJ0b6IbuGUsi3SF6BkF
QoygNGeF+n364vYbhzoVf5hNo7arJv36P02DGxLrBWkdMSiWhUFB+wQId2l+W5tKxAfmHQtD2qwi
yNPxSOG5FebYZYdWt2eT6eJVa15ASCyMx6buYBmPZvTFfa8E90SwHO7VdrguagK+kS4TI3gPAyJX
7szU4tj1NjtCBXMxgekyhutdk5ClWh4KpZpf0mJamRg0gMpvXvx+SIaidxf7GRKQiZ3jIBDF5S6Z
dIpxl4FSfNFBB7uwIaj0Fg5mt3P1MHFVxBJXMiLubJ2tjegiRreXfZuDxUx3hTwgBdnDpwlV5pvp
7sejv3PxuX22hKixkMNFpCsZYG3E8udY9+PYyX2+a+DEPsoFqGXHPvuIU6IwUZ7YeC7Re35d1vKj
Zh09rhIy/g12pv09CJfb9+Vn7PP6AbItWMB/u+RONDV+901Q6EtAg1+qFZkREx43CQkH1rffajLV
KQdbXfqYM4FATSFseC01GuzIwMq+CBH8P/P4ypLyv7Cn7wjai+/YlSraa+4tuy4Fmrpi/f5/bJdo
y5/ja9WHpc2V3037yys8/fRNL6glkeZVoF/WOvBQCpJLKf+PYCodd6ZIFg/oJSDsQzBGs/LMg8UR
RsEhLj1JVIMa/oGf8iL4+zSXZ9AqPv6UXL1SjJVbcLLilDqTsnwiEuppAjVzJ1ak1CBa6Nh4OqSq
phF9bG/ZXUBXmKFT1QVwYW4MNx+gMZn+YeqFxQR3XpiAOkNZRM2cfybYnSQUMBWI7nODQRhbp0cH
rzkVcobwuqxGwAU4a4nS8cqk16NZT/wWJvYlG4ZhCEA22zVvhczajpiwKhLrxeFqwnY0CH+fb/LP
hyppZbfNTd6H7czqQ1Rsb4R3kT2sbOt1UYxEqljykSbOwtM/FmL6PevzotvtQsA5HcVQmRz3kypL
pZUhN3oecllhCtmEGyHAIPTNvuHHY0kgx2T6/X0JjpHAVYXVi3MkBEA2MtyQauSJ4AtKqAfeOp4P
JZinDLiS/k3MIGFkm9A+lQKwxTfQxVPVQE679eSEa6rsQeLGmrUPJ5uWg1XIZUJ7CFWnd6+VmE2Z
tNqdHGgpBYkc2alwzL+Gf1dkbUUUNleidrKXvmImQypbkj+zbtr2DW9ciWlK8qUAxRn9yj0J1cGq
oGxPAut3HPQcqCdWBTgM7g3O7jcMmTqth4TBrgNpX/r45zcu/ju3G6aVA/UFU4xmkhr/gHSNxGK7
uJFPcCH/LAqHVI3Bdsq1q3SW+db/jDwDXzM6yEhRSNOhhPRnJqE47djBtL8W9rcet12OxbCL2YXM
LKqkDMu28WHFMFNmVCr4K9T+jMQMrhtlRkpejUbew1cv9Dv64ckBNFun6pOLs7vgPOY9Nz+7dolC
nhiPiboB8XKUDGIdlHiNF+IIjfM8a/rR/65etjjgQRCbPvqVxNsOCctuBUV4SiSvMvzppSn2Em2r
hXA0fjsxPwXR6o3Hryc5oLn1CvqkwxutPTOMNxB9+u6PLqaI4A5TUgcLxYMbfpnvbqJ+6JkxH0lB
XdfG3Ij1iJF5Cz7GwLJisQVdHJVK+3T9vmohXOK86xqMQdX3Ziju1pIoEBp5EPJXVw3RgOx4qILR
Ebo+c6kAS3msX18akrqgtRjUqkhngY9Wv6c6OFsX6Jzj5//zW4uFUQ33dOCObv48R9g1dPZQIBAH
7yc7/YlrLrVl3kpl5R0vafH/GLO7ps+3g4Yeb5amlOcU6O/9BD06tyqJGvYkLFzqek61T6aC8JEG
KtfuPNbrXZXeeJVSHdr47cZZZNxaEeN+3urPnhQdDpiguXXujEuP377ghHHkTKMibfvTJ/sf3rav
lr0qL4NCZ5vrBzDwsO+G+bBMmmVESf08x0MKlNE+PoyKTN67R7kWAG4ZDQXKYGCgVfWKzfwDGdqK
v3qhBw3ja5Pk3Gc8hdW/8vL5UhXjVapaU4HPhondJy1uTao4jxUT9aSgQ5VcUjKuXZC3fcV6GPWr
CPEJvi5oEEQATquu3yxiivGNhkMY17IK21EqF+o7/S4iubrNq1287ELqHL5gNhc/CXnNNXqY6oqx
HCHB/QG5oETHqsKPeRTdDHX3yg1zqoekBdPrcNas1FTPdZV70asE6nNz/8+ZWvRURBLk+DUBlIey
c/4ES8r1Ya9BZolQyxQf5HAOBIbThJzKhx7Hfb+BHs0xy/2Zn85MqUWZYDFS46MPic2VSiYUzqBj
vHspnjsN2HfRS4M7+8bpGNb7QfGwYgswOXgGhGvaJ/CAxch6cQxunXcN4dNOVLDNrAl+Ut9UQrW3
DrV5nqIKOQEzSuHKfO9ie6BqPO7HXEanf4iXgPaPtI4e2q/a88xm8P2A2B0kS+qiJtoFhK9YxTi0
ypkYf2bZQa9NmoS1YmnlsjEI4SD7OKMHf96dRR1mwv6Q+h6gHG3cjOTnPVFizGopPXujTqcCzuzx
LZb3J5rSv7iUaBhjum9uT18pkPRTnMGcLPRx6nr1/wyHX/umaow2At0SWHvaKVtqZlNSbqwBhccs
5pZDwFHTKpnpI+PrSdLgexX6wJxe6zp4B0+thJnqqBP8/I9FGev0+z+TXDm70tipMZYq5XYxLY8Q
mgRf001bCFdWFzYxjyCe/toJR8aWA6Gfnpf5rw3wHtNCcFx+RqCt5DPQ6CGItKHfxgl5YJ6d0tHm
i35KM9Ge1HmHyeU25471gVvUw5AZy3RxtbE186NmkRk79lt1P+Rp8YQo5g//wCK8sv7tCcKfV/jA
TVdQSr7lXb/bElm8/wh90mrdWMtP2BBM1GiVtTbFH5+frJg5uqbofqbs+jLIgmy3NalCjYd11Fnp
tFs9ck0XyYtMnx4bVK0UnNgQhMXtrvDw9O64yBljr2kaDjmn4KoaodZQhmU9FXMXaZczyPEWesF6
FTQJ+PykViYMrgO5WhQk4ZLghEqaQ3PXDNs7cG2648HKAvdlPGWHiSTVx8+1fLURRqVfeMRpbxWz
JBNVLsXhyYg3SesKEw6r80Y0Md/In2CSJWrAOfBXsJ02u8Q5m26N/w+X1H/V8VG9UZgQ+wAMthcM
flY0CdnE1cPn9SqHwdYIwy9P5bl++3wsmoMiFYuhVVP6i0GLQZ8WEuuuwIg8M6Zf1mD5pCrL9IvA
PJ6bTZlQruz4OehbEh5eGP/EK1C2vfO3TvAKo4gpLAw+awh5ok5tBbw9fIms+aNqeJd/GjbMSyeS
s9KYgWbzMgFHb1Kh7NqeKJAbnaiqkadIFxGNsXOTEMG472nMNmICYwfKNlUtG0SJTX6+QyHTKCh+
y5J13r4iznfKJKNOvAKcdcrW025prpLqdnXOWknzGxX7jWh089lxoNdMoqvyP/OoXE3CcoOojCqy
0h+quikoltwrgQXYi0bedQiUnSXemOxAsEjqSJsU+HcA2yu4ioqgNlm5fnWdZIz2M2hw+qgwdU6d
ripkZ0sZaOXRr40DYYjblkkropNGCiUs2zjFf7f+wLpvUZKTjZcsUisiybfbSJCpEnnoU142xGEi
9ytMgXaq2GlY1xnspRqmoNSwefBQNwMBj2xoRQPPD6HcSHwEo8Czmszvv2QpyhjZ2DhnBbjepYLt
9/SFaK6w+yibCcJfaIUF0rFTIuKo0aMmI9UR2v3ZjFhqxmi5PkmFz+8scHNNG8s6tY8tE7TL5IP3
kGSCbvODREnuhRpDp0o5/8SluAES8Pxp3Dhzm0n/3QiR96x0rJDnKeHUoDUG7EadVPVTIMCF6VI5
svRhROtroZo5FYCjmKdIcD6BpTqdu6Df0NnufA7hNlSBiYww1vhUXecUGX/5IvWjvEWrD+d6Dy/t
4ZjJULBDcIoVQZuJY9w+XlXzKZ0WcCv1N6jot+eigG0UK85a6axY+DjzTusNG/A6M2yHMrhHFQ5b
XuE6KGtYicJrkkKOJXELRZAls6kApPrTwrPrTjMHCGptHJhUu5gsVu4be3S0C23SaPuLUX2TTSGt
GrBA5r+TjAuXWpnX8/byAWrlI+TeDrfzJIB596mzyiDRFhJNpHw7yd5mA/2T0x5kzH2hvM/BeAFf
h1o5Jwhi4GVTqViUdnio0VUl1FWOWCkY5GWqPKwr8qmnorBjJYQZQxyc4ywDzlJA9k9K249dldH4
zORIGzagsfvGQNkS6bGMMvz1va5P67772vIqL7UYxHWP/A3tQTzbjceIHWIFvJevPjpG4qQa+BOO
Y4vcZJQN4b+xXlRE+7QDIblPPti328TeFYpyZEI21WIpMAgXe0Ie5PzOpEWYEyAmuBT1EdMRHL2u
BG8Q123QepLow+zY/hhMHmb7OZDV9ufxgkwpzNfXazbbDMF/TSpVtcIo3P5c4joo2cSvCwoGXgs6
emALXARffl0WK2lIrsaYLNFHFNQhIiRdmr8R7RdcjIpIRY9DB6vQtiR+dYqXtx++AdLxsf2tOJcM
MX6LXC1tum/Tk1y6WZ5VNJYg55HNMOp+SxNMF8lFimOmGcpFZ/rMZApfvAXtuh+kT+I7nWeXsGq0
gJV/rut4d8uz9hSYCoUzJFn3Sn2uyYUTtvsSIhxGbwozwRyZZ0o6/Lnc5tpOZA8uKmDzg0sxcEyy
xPrEZCBW79Gz+PiZglAYkmroaoWC4JOqTZqV3vl5aS5u1ikjjoRD30069iAt6syzNxZes34kCVJn
kFZth7TQxERLseDh/efFVPjxBzA1s1thBN3pezrQ8lnapMQ/uWJZK0zP6r57NuKu9xn2sKghgNAo
oGvHV0QFKS7CmBOGjRJo6A70G3zYfxoCc4crwzf9YW5v/AmEEBBYjvFuBMOzXVzKL9+Vj4/4ptZS
30/8BwBuwmsS4W3tfXLgbLKYbqvKSiF45seLWSX4HZEER8qJQwrVV2nlTfhXknfhJVU5xCWB9ZFV
NBy2RxL5vomH0H+AAuroRyGdtypvquIBfRKfSKScmd9iUbj3YzKAkXs34xuT6Po7NqNvD7KoouzH
ty4m8Ce9DNxPiobi0sN/f45tmglv75tkT0zxp62xPLqpZfxOzWthdiI3NmL1FjeJoNeVcdy8jYn1
kC1xoODWmaqCFhRsY1iK6vfaMmf4XyFkw/Zirib72DNSm0VDQJUDHPIVLrB0c8pwSAppQQGEtLLH
MjPsnuOrod6r2U14HEuoHOnCCEoITA7DbIoeMfXjuI93c4cn79VEM9NjYyLZ6T7ugAJA9jcvainO
m0Z0BnY7xA/2V5vGS9e449O3u66InM+VLYHj9jzdudcC7dRX6/jvrm57LR3OYDbtWQq3esX4/5yR
rSA/7fjOg4Ndyha59cIeMVo6mOWDyZu3f3R5c5sP+7FcbXArdYa19yvzHMBPwHzFMIggK1I8htnk
V84rkitPokYuQs6DLRFBcPYnqL4exfqm30Jt8xa1WRmou0PMgHaPzvkkHhnqgKO+54ZBCFKjZi07
A/vUmkHrEEaswoe8V9s+CzWYyLjIZH+0JInH7CQefAdjvhl6CBBBFtlMLaqXFfasA8n4G8zqYv/3
kO7LN7bAvFgqybPGoSvBGfMG8ozEqHwI7DqXg7jyAOtfYhPdcfb9ylKb0X0oWlZ2zRORxHbofOvv
oEjvU5LWDcPQ3gwxE+a1WbjsiMIqkA1YAganO1v1y9SDq/IxkQrf8P13Zsq5KrEQxAIN7MDUggVF
VZuUrTe067+2wpBAHStFeiUZYKGWdoa5K2Xd8AoME+2Q/KslSNfHTdCuwN8I/UL0X0JIVJpGI0Cg
PeqTeCoitj9yraZFhAx+KgWZJSCJ8DAXJZtwhoyszDdlWEnbsRXyJN3gjlgOV0sZaN6ix5Wb0T16
15T/9k7CmvVwXlDTIxfsmQkwOcY6cE00b8gPC4q6K+dgKVPHOb9BpiPdmrmUAW2FUBSzzwIBzfEV
dsxJRGS6ukcNdFAE9YHT9LRAlUqIIFzaFVN6fzjfQ4NDst0LH6lh8cKcEUkaDTCheP1vyamNzgjH
kUyv+QIoDsWw4XKhcX7ZJYwWr4jYY483F6tTrFMv35EmPkT+dzCvjr1x6DlFaXIcT3v8frwpFc5Z
Eksi4mh1hiBOxDaS3xbL51PZaJB5aGaktsJutIMXV2xFsJ8VNlhnytxJccrB72Ji3PrFciZUD3sn
4S2ZkTGdqFjV31vLmCOuZO3uNAP/Putn34JqlERA6aERq7k2jrlibzEfiCBPmnYtLFOYL0ojfle2
kZPoL3t6At29X+QSBqcwwHoNJGTqw3EhYwpKkeUlkkjnxbbHgnH/3RgPOLya05SfMt66b9N1wlah
GgZY10pmSDCZwFe0sUr+OZZ24KeVyeRNacg9MvGYSkdPqJ7I5myepc9snzZGIpN7GIbkGmE+U4TJ
KP0qMA01zHUUqrRnb5umflT5Qb7jS5qAaIWokosM16sdS3/VCtwV11sjV8JBhZbyfEMb8qKY4rA1
hnz4DwR11KbvJbbW4AB8ur7DOfTrs8Fyo+v8+QSZf+M7oRuaILaYWiiYHIHAkFFEENvT5dDbSDr7
PRHZLB7J6zptpU624LKzQ8H76PKAo45Nspl5F+YBm6Hjb2QJuwTcFfEe8rXhpW9o0bvd7Qy2DGml
ExqX4tFZxbZjTU4OTP/CMjre3R8btQax6CC9p3hL3JaAut/ZAlzJ8mj8JHhJt8Uao5kQu91DBSs3
GzlNrBToA6dHqp+TBtWN3m3wbRYv4M/5R38/o07jN3M2e+QsYaFLltvZnBaoeU0LKeG0UMLyY5GI
IMcC5eTei0cORZXq4XHcw2n/ijmeo6HQzPo7oz2WO8kc5c1Rvg7QBKJKpRXlgZjwr2950Wjbz+TB
gMJUOqjYVP+Sz1S7Z62elCmPsd6hjrY5tVsbpV5kr6T7SiH2ZWoc9WoIMMqpztGKYEi0u96pDXB/
4KoCmSzcE15RKLgrBY7OQxp8aoqzSQm49HxHq+cRziElq3M5W657m5rzvfcaxa5X1PrwpDFUijSU
TQm3TXUk1lL07nBUX4LSIIhwHGXXpTVzpg2oC0wcbdAnQTGx/yOmZxeAr7HDB6Q5qUb/dU+nmKRg
dUCt4hhz1ITPUiWTYdjzokmnah7NzW8rHHA+sPkY45F0VkZs0YmMLBrAfHlG1WRTMwRZV0vxdE90
i/fWdgWK112UoyR8+WKoSp2dPe14E5iXcqnqLQHKAyVpGy0XReyq14cc1YXHVDPeuESFFkZPm/Kw
SgZxoKoFaM/NWlYvQsp8lHXue1Ppt9k7G7gMN5sxX5mxBxasHTDAgYlwAwJTIcMiloPYyWzJVqfR
rNkilh30OspJYZHMPAxO3zsghI7IRRa0HKSZMXCIdWbQ0PauYBi+f/VPXvRVPwT+ZahF+EuOq2A8
/GsQ4oUwLzfHra+wYGN2r6Dw4KHVyTOT7O5JFKvB8HTWrt2L8EFfIGBrA54UwZ3v+aa99s07UrdL
p5M0+i7khHJeVFSTrJ2+QR8Y70TULSc0AaOJvB4yxtPRHmofErikeWuXIc9UTjelfkk2Y2zd/dhw
sCClLLDUO1dlVsdEUoH74XAtdguSCm2hYIr8bFMc/1sNQwaMDDNA9dUXmiqKRGKqx5VIi9BgNS5p
Igq1h89+Kq9s6wTUnsQ26idXmAncoPZunnCoHgggnyIgFCULxHTBvhSJPt7PFRfsDD/QhBNGlDcy
aTw2VqtOl40TtmtHACpwib7A964WXu/EZD6HVQu3JDY4UG3GamcOH044zBEoyoBa0RzXvPP0mp7H
/jSFMdZF2zPNxMWdO8A5e2gwrOfNmX5A6b05RmjIBsMg/jsMIeToZ9cm6XmMj6rkPJ6uYyHKE2Kz
B00JOl1I/6O/GssGOtedIxFTcwpu8jAwfPQ2T41nPwWo47B8pmYcOh6yc53GcWC4YP9s7t5yca++
w9Q99scMZ0N9BUA8WfPve5yPAMQ53P5GHDg49FhciHZ6b5BQgsqPp6Vh8w/SCsjcq7rUh4g/2e2I
o5dVLILTg5qFwjUODeLBwg87ElZtJVITBhOkKzl4YRg7ydqBpc5Kyql3pFPv/bE+wj8BJm1fOXPR
+F8uFj9NmBPOkoFf8Nm6VEg+SwwFEkFp/98kQiQIgOnbyMR2+/OqiEDOZaDTAHu+RpClfZY31k1I
RChRNO9zd0eBH+sBG6o9Qne1ZQm9QR8tJXMu+gWH3M1riU3l67tdD29TPxW+qFBqQsVEInu8oNHK
MgsSKXL+WLSoXg3g/5lFam7Me5z8fQHUdZrvW7vBU51dfdPbTvztOsaXPpsDpfOtWUYHfDaiwnMP
VKRfxAfrP2EsavJfO+yZoPOLv7cVJ3kjKp2afVORT+f8lxWLaVkSMpg85ca9D+qfi0FgaEknbEYW
d1h+znNZkbHPr3pTYRjQkQo8YBC5OW99PBCIDLhgZPCVhFw20cdSFkuu39S4yghhrmvu7nyPaqIT
Eo8U4qySbXRCeW8/EfrVPyXCZj2WcHExnK1Ahcf3RZdRjTpxJpvRPebHnWkJ+Xeh4S2l5hVnTwLF
RsLXg/YhbXo9ivBEDiTrh2PARPzj//Waa0cOAtvvLvcSe24lbT0ei/IWp7y2U2017gtjg8TYFt/0
5bVDPCULBoaQmq8q7Q4gcsU8vYPz8rqJ2Z2A/RZWHhqnfkDsqMc2yt2G0GgOS7oXc9tEvJoGaSxk
RcdIZ1qxe1z+4dm0U12lIyIubwEu7gUJUuXF5+Xt+KzeMY6HR4MWeAns4sxcq4LiwpPCnjcoZERg
ODl14Ynow4PZ9pViOQ9l7gdsxODpl61/xRfVFlFcaYt2TfIL1tI6DGsHIIhs6IOCHWUPnyvCCrEF
u67HMR+6QvJCboSsuc2EA+IfeiYOTm1PmrKbJP0qLMpmLFk7SbUb01PWwuYPmeYiiRmOUkL6lVQc
/6z5wtKn65r61TT8v958PF8OcnCIu3VLEbgdJ02jOpfkMZASSIE1sK5WJAtBwwvaD3k0FjTLQsFu
ty9Ws2aFYlmEacz0ezMe3gqWvCZTTToDfJJeANSNLM6DYVggK5OqNPfTgxFICmz16eia2NnlbK5F
uv5FJw/4TYAoRaYvfg7aDBA0AwvNi1Vt+9Qh82hgbNAgbapxZ2kR2EFP8CB176vkbUVZlNCCh3bh
1bUrrMxVoqo2QeokkcEsIkVgn90smsUYjRIKUlY8LhaP+6yAtkh4aexRyo7vN12PB/bfBklcE6xv
LKxBuKbkI1zDlELuB6xoBx1twf5K0JFSRgUwJsHnAJDO1Fy2nV3MTopTdCDd2ykiIsFW2HJ+VAIV
5PT7v9uvGHKQPftzoQurP5fSK3OWgt49x4gt6Mcu6Ihfb+2LZbvsR11eMyxMfYfqAwZ+B6IlEdGd
4BZKPcXY5rBXv7lzg8NsiLkKjYVdazpbtClof3gMp5ATbjycS45dDkpTW2RimUSVcZTsyJJPrNdp
wUt+L43tZW6WpIYL4IoMmDyJhOjr5wFN5Fp0mtOW9Smt+1SffNdEtGhVt7sKHW7xDmqU+K2aEJuX
9zSOylmmEJdQDMJCAWGc41Yli8jtZMHkbPcpXPwF0FVfg0Zxvb8ws9/z5fc+fEBn5ppSxZt0Ez19
ByYndrs70zFUIT5KTV4GWEuSyvR7Rv+9q/XocCas92F2kSGsQAQ2dksS3H/4vNmjHaaKSTj+vsjx
p6wv9Zp3EikSmBflnomiDXr79Ju79H8XxLzvgENCHTlnYLI6VeDQ4dtucX1D5uF5H0rtMDjC1ny+
m9mReTiaZe8PP95QkxH1S0bwyKPz90eoBDOaMMjEB5v2+Q3gkVvlTFQont3nWY+W5WrOXD/s5Hfo
wkKquJqoC/6xoFx6yuo3tLAhl6DBU+IkLtA7hc2mBrbeLcVz+3xgDgUZ5swaWCReKYxVAUs2N6n8
uwIRvKKXgeF0EgE6i+FMG7cbONKJgqrI30EBALgACKxv4Hlp8jSlH1jWGzuwIdoOl9CvJeoXQ8za
qTwqbpUmq89LkfjCp8Zwff7QkYSRW3EjJtSHoMKZl3S6O/+FUfZApkM5a4bDYu0MREeywmD+vzhL
DQ/irTm0uQeBG4qk+U+gusm4QULjRgPzqWzhhUU1iyMFPBeF2+OlfLVMkHHVy6eOhtECiFvCBLGT
hHpCU7qnT/AtPL1UBid6nGNvXnvR4Ref/S/AoeAOPBvlB+UKsiLLLxxxM+AHsBV274yf7wqN1sSX
ZZAEDZGXBYhL9xMiz0dmPwzOhpqYk6orHA7MITGWes9dEQrxhmro8UaEnCxewbVyAbNHKCF57wyB
i0O7ogLaLM8HvZmjUJ+gpH20yEswugXSF0b0xpcKs+InlovjLj5EPvd8GA79Cu4MO/WU1I+7Er2/
gov8VvC2LhB3lE9Mx1T8TAVfdAva/DT9K8rhm31UnMaAPEjcIlSu+aUxyuK0sWC2L+FN9R4zVQIi
eKa4K192ef3h+knLxcppkcOsiyNEP6CSusXiWZbnW6u9YT1oDK1P/VRJkVEQ7N5wMGaGJOzfP4Pq
hS6ZeVuvuHq1kQZAzD3Qodxnt4yb7hLx5O50E38sFS0xTlQLId7upbLO+Dt7qNNM3rJMsrOGU9wc
yaVm9vePdVQ3aflfnlSmQ6JtzcEzx+dKkTgkQpZn963Zfatdpt2ImkJAFRHbD613RKcjSXeMrNoB
V1kuZJh27jirOmZuMDQi+9rjAk/L6EBJHiI18iWAdTBXc0zOeHvE2fX36Pr2nF3mSIHE9bHvacvh
E4RmjEFnGkJtVpqJdaZk18JeXMfCT9/okIDSRAkG020Bv96V+EmJZoB6x8aQzwhQTspwbynH1zED
gHFXscbUldj2S5zSMJC0b0OTJsHER30B7qII2cL8Z9Y7FEKVJ7gGlAFdi7wisuqhVe2xplDSSBIZ
hlUVFKWcgSNr6tGrh4GkyDfJb0VDzmPrQr76/SVl/5BXJDOxf/uVH/y+5Wqv1LgnsL+t0Scy7Zli
TPNWOwP5/XYIl0ZY7FVz+qdg6HaYG2u0jJVNnuYoucwuVSHvaguRsyG3Ic/tj5tvY7e5mjkNr1m8
xlyFvI8nDvlP17pYGGOskEYf/KhqFPSwIvwLOSxAms5X3W4ItzbTujXqrKkz9YkeCZnoUYZB6N7k
jkZFK5t6nyCTFSfqYa7Ak9rCo5APyKy/MwMfhYz8WCr7As1z214uBMGCwaVKH5fpCckRboKHffPU
TpgPZaql4XvbC6bsH3bcqSoQCUtepPsLlKTH1uod6Rb0as/kMeBkoCIzCNjBIGL1IAxsQbb1nPyX
CQVLm2FQY3eHbGwsnCXJwIakvK3KPNI2wYS5D093pBKgs9gj0X1wRHsqZwqrp+rMU1oBse1X6oH3
3g6MiHyxhxKdhHnXMkjmI2cdQze0gYb13RGtqm+M/sgAkId+8OjXxstMSUpZL1A0/d1+mJ3p+nuO
6LNmQ3gZArFqBAzje87/ucpZUJCMU0F4WZRRFuGK82RFHc4ZLF4DzxxPMPcMjeOgu6jdJVwA2ppY
y6LZ3/fMpxFUxLsm1J4I8knyglvjlVnRQ0RRZVhi4AjtxpOBw4MMslA/ycHsLEpqgdybgQI/hilt
puUeZddFn65XDqEkPQV7b4BUYrVWcCHKkXVw9Ahf+wxanfjmEKjGK+MzjzyROKw3dTh9R92cj1T0
+ayku7uo7GgXARNfqBykpSG3kT+VofETXQqIZOe+kpoYb2Am5xpmprxrlAHr9RJKKsnksH7Jqr0W
Tj3T3SDXiNJV0aAFMMA+rypEkmiGJSYFF2Fp70pdY+S8NiQkGgZ7JtipPXhZWjanbfqSF1nm2iuj
NWVLGzP0FkezQUbUs1bwfu71L2/W3ier1+dF9+HZXd/mFOXBeGfVmiViGtszMyFXtQ87kVJhYiOo
T0719bhInpVJ3x9kOQsYzhCK4mFuDl65Y7NXhhepZbpz+pAc3m//qyrBpXSiXN85xk1EyeNH8v90
GR/cOHcR4aONOjRPeJVcL1Cn7NFAEVhdlPsqNgZHz+TVz2YXZekRoJUEb+qBonyu2MPoZqHHiE3I
jUxA/SMTwi7HBB/Us7AjVzLh3CEpy1FPklrk5CLCE7+gaqElRkH0Y3aphQjac+WEuN04O1KDDUHH
MGPWJeqvnH+/oZGyZU4JIQGCe70FSlQfI1wDtfoKiaSXXMl7EBhfUnOwDnfHS0AgqfwJrf6JdKhc
LXSKMh6g+EWoWeCKrj9wcpuCF2uRcKyAN2GtFvxvBqNlV1qK0JE4BJ/CipKsYeNYCPaT9+MM1rGD
fUMtac3qHjag6Ny6NJefi1Zuepzsr5XnMJrvsQfq0cWVUjMnmtHnzQDBF//88IxLMVR4ebGiqaGy
QMPdB1YlHYtlmAitjLeC4PrHQHdd35vy3HmJW7m7HcVrMoXxrDZYeBWNnK5y1AMAHSJxnmfkVya6
7/3ST+WdTcohQG95K0MhZ5OKAUHom8g9fdLw4qTVZ0q4tdaWk22XKxXiNnRI6/uuIQH/pscS194Y
Z+OM7YUUDq1jkSAZwJdXNvyqqgs+5zYyPsdCR9JrMWMv/M96TOTU43iKlmcq0dY3MhgU1h9iUcIA
cN9JH6po10W3fhcpXTWMWLiUgg0i/8zsH7v9OcFUjjL7FaIlls7umQcTv+DsZGLE2ylLHTZUEYML
cjV5SR+u3zeWadxj7HgXUSM4Io6/wj4CgQ4Vj77+FIY0ivrh93Ro7P+rkn5uvhpWcEIrQt70Ft6Y
A7qX2oG6/SPPTnwFLxf3AusXdgLUjoDn8jdkLRqiRnAeTHxYkMoOjYCl73V6y9z3GD7VRprG9/l9
arSc1Ah1sFZRH+DyCHabiHghZeqb7pqtmlo9ZmHJ4A4b+5yXR+Yk6WbNDK6KJp/jm8phqz6aTGPp
+WlsXXaj5FPlpxXR4zuXJjVoZV/yIt6R3tYZrAicnhSuncMUFBhobh6NMgjX4jl6NzyqdSsgmKES
YhiW3KqKe1cFbcVjvv011deURPc/pk5S4XfLgRTPZC4pdsOHWYsTwJr5zaZ8z+/7sGx2DGtoEfP1
WIGG2k9hodFI65ctAkIB/Qque6qFi9AFvZFJamD5PEWE1ELdaUg1lHibF5hnvr2sA7k5loxMtEYg
ja3lw5ABgF4C3ZspA1fKjtjD5p3e8DY1pB0MhR9sHcr1MKFFElSdHA2LYat+BEseRuq3qmet3Vg6
HGFdaPlEslXCGoO88QZ1Tu3DbPz5wUUj/iK1wypq7tfaY3M7YCCZOmU+3RUHJ0/A83fUxhNj3DOG
Tt8cUnaClJcdGa7ZtqxU53y6lHBx+q8J7HCUYnQyFDviCj9xoDvBG81KUakLmTx5NirizxW3pigb
gy/zorple0sttRP6XRlWYK6jzZvA/ufDezv8q7u3wXcHospeDQuD3N9nwJ4RLvaW7Lx/WJHXSySH
bMxNsUstpK3Xwl9G7zsNLVVqFXf97a3yN+6oApBddPEG5StOhjmakaue+nxqcaFNXhcgLpMTBzus
b1E2K+zeys0cEQY9J7bOKzV2K3amcApxdzrNXghKRB+ro46sitPWRhObotp1Cn+fY8fvFr/63ssh
6d5Zhzvm+Ipu/HRqwohORsrFHOV3nEC7Xn2xZ3fSLKg3XnTi3VVYOxCL7Rv6/BFQly97OCFfOkvZ
OPMErMLcr502BjF2i1t7Dy5CSJI52JlK+rW9Qws0zFYiSOsUvhbGx2L/z4IDDdcvxPe1VAi9pNeI
Plj7xx5vpNc8kqjONu47AKIaEsBHX4BHOf7yVOBa+jlb5qnze8hhvWCESroLANQ2GZlL/60L3q6K
XPrHF9kB4WeUkdvdLocmlKtRKb5gcsQbwLBeRbZw2kC7l1wbN5NYUkduc/x1UIxLOhg5pWEr7X0m
GdLoS1Ivq4/nxM44VU5eadjDkT257PU+N8uZgEbTZrHjGbvp2a4oUj4xCXRDc4fbCayd7zN20Dro
p2QWRbwmd0DoKeDV+T43hUf/nFKmzw/cgwEJ/TEwT1O2bvD3P6BVBB9CJKZ5WeT1NHczNluQRlFf
BObr6S+1FYDT48WKNpF4Q1NfFp9fLnS8pu4HrcsjrFFlStuEgtxmJiovV1Z8Pq5W9uwSC7dXSCTn
X72pHWTfqMIymV9pYeTCI/40qL3b/tK1ixuLbBToRBTu12ilVSsNRxHY2qqZDolnRK8y/llMYGKH
0N+e8fPYtHuGF1XDLte+jnukMYvebTZG8WRWhvc6FN8+CASR93x8CRmrmULc16CSC3am70i6nboG
YyYAL2hmP5kz72fW8Eq0OehzV363W0A+pKv4qG4VOUIbDBk2AhXhmJVtTlTLt9r1TVSCnB9fG8uN
rtaFvVd6fZdH1a6CsxI1uWCFvfAaMMaeb7R1AINuuZ0zDC5tD+nl84hz+IgQqSxLJ5xXpGwFi1t8
EAgLYClQcHRgA7T/cY5emm0gXiTMFAPWQoScGEzjByQ36uqegxcZAwrZrFDkrfgqvbbtZfvbc8+N
AuY25f/Kf4x/8Ou7W1UeEfMVarwTOxlhA22RM2KCEZfHg+aZzdEoVGa/UVGi7yZG2500dSmVQcPG
HFPI9gXqNpLIK06Zir9cHGJLJoOwFAqQrBshRxD8C5Ua0t/lSqa43HrCw7OU8mnV1feEUbMzqDXN
FExZofkyKZl9c5cW9Qxxsc+eto5EjX0TMbfj6R9zNCprewOCI+eMJ02SDRCa+jxo+AFo2+3/vP/v
KZJS6qr+ImdO2Be3MZArp0kD+kf6hgMb0XEjDVHh9ad3/un7GIaCcEhrI25dY8dm86k+Xfb62LRS
h2GDLMKvsBdQEUYuZ2XhXrAn3NSt9mtkDSU0M+Cmp4T6x6ZOCcg+wKGOZa8m4/01jRJKw7FRFlq/
umN2FISgrVjxTLLoT29oKUi2Glpsk6wYWzB31uIGnkg6+VPjTsT6WYiVqgqy11eGlw0ZJGzkeHzL
8M582FigNX2lpR4K4iO/vuXRySpcOpwUhUd/N2JfkPGSA/dVN9Tb0tx5d+D90ceHAi7HTwSEj/a3
h0e8p2ojZ/Vh8LVRBkDfjFulb8DK44vyAykhyKWjxceoHS0Y1b40sM1Ww6unRBZ5ScYBZnPLuNsP
sNrbqZKaUJJBSuXzw/MzIcvfE5lniWkQC/fHYmbVfdEbY2sehuxkDGF1oVsPZw7NMd9ZvfTDbgEq
fC6v+3lTzool9JB3UtEBMgvqJNeNue5n8qQgVP3pBmxkyrn6ztVbGlYr6qevp0BecGEVUAW6ngZj
DmnlHjTgWRNWIwkc/zp8LsGABwCpl0EGVWnlLFTvmkttefrTs0A6TjlBzTi2IST+xzbOFd8wrhNS
48jN5kSEwzilJ2fdKAQqJc5r1uUe8ROM+Qv4sBGLVCN98mR7BPJMFnm56denfkw7/Zd2fKSgAYs3
ALMWl8+TAhRcuLTvJlz5tBzE/uvXSIMoPIdLs7pSk1ZHwyU6S3pAGcRINefK89Vytvc4ve4UAEc7
HSgsl9k/yZpRWuZRRETJZchq2+0PyCJjEgZZCNFJREq1jzkF6UH1k4LuSyosJ6io6Vqh5H7nGjZl
VCdPGdByWkyvmpEWxB2iH2pw+dFtik2lyP3hZC8B7kzlsFihK0rPakiMoRTrtBlVhd+Np12cwp80
58IQj4xaSZr7Gs5MYVn1vjfDIy8hrY1iWZOoGlaDwfjm5fusOQFakg5q9zxwH8bJjnEy6EpKy5z3
GMYG9ZWm1fiPNxuWWlWbN+Rb1p2HDmJqWJnwKrDuVSfqVvJ206v1ID4g4dD1+6PI+qWH1JtBohzF
h18/TjbS0q7hGmGxpjpTM2R22sF6aPmgB/T9VXmz0Gni/nJBqeK26U5sCIOfxdehwqOgt09+X2lH
eYEzodzKep2WHk1f50OYZVZbEpbRWdcz+cUd2STAUKOWnH+NgcnjbKV2kGBfwRqkcSk9V3wEU6VX
O+TsZid0Mkz2kSw31sAWoRMjLKlmP3xaQl7UiRFJ4hqXN/WdZd/rfMfC8sGbhYOqP5kJTHcx28K6
w7YY1zBK36ZnqaHwddj+1/ZdTMLREHBQocHftrihlbVRBBp1Ex9w5mAmOiIxdBqBmvkjOsRjSyUh
lu109euMcmr6+OnXvxt+AdjX9Z8zEshlZUERYsTrzTWpnX1XSKIh2NkNzMYNgjFM4sK2ZoqViJ26
/XguNNU66tofSKt7c3EgJ/pxcXfE0pDXQ+p5Gu/HAuyWJByGo+shsElpmKyUE2t1T9YQN/RFfSp9
TFtwQsIUiYqrwxrVXgsNL0NW6pUY8K6zhJcprN8+lINiiCOzswzff6ZV/ujVPzf9Cyn1ttlmDpZF
ijkSoE+XIjpXVpBHCXW9JGLeoJjeH6nJpftqwEg4E7nioyJBLDPMoJBcUCQa9XVXp9ienn+elOTY
HGNe2zGWR0lDm6oY89V0M7Y5UW2QvV/ei91VgWRanWGfhcKDfnQ5IKdExw54hx13haH4Ydms0MZG
9YjTy8c59/A+j4RtPpgCd2ExgNmGD5a/IJTVLcqz/3Eje1gOILThk94Ib/pYP8WluNRepn1r0i0y
3cmJcA+lvCf3A5mEltKJKxpKivPhS4U7OiSx59Zs0pc7oQNVedbh62A9XKicjmpeJolOJVvrUa8s
2b8vEtLkieaSkOtsf9Uz3KCln+OhkeJs4mcc9YdnJvgT2Hxs94I3fVb1xmzl1MHiE6w7+UCno3xS
eTvWa/bfi5utkSUjlNJOyDxn+JI2jbbgRLx1aJbnVi1jkiidDo9O/k5mBKTUQXxyjoCD5J5PopyE
FWIvtviFxr2zdSVF2mBEXYZAqRIkAkkn54hAXo0UFtZhP3pWwrqxMjPyXon7ts9ELReccQu5R2XW
5OV4aDUiGJNNgfQPgQsUgQMgOJfbIrhvpT5MQiRmcU6nlCxI9lfOuwdLP9vh4YMaFx60a01BGYlO
lGvxoNz19OV+Ou0ASlpucHGFAnK76CIIC8WU895Nnpvun4FFTdnEpUjotmNMuRzgcnZseGFyCnN6
lI41MpG29WMLSSiJR+nViZJi/vj3W4cGRNgwoO/NkuFGkSIcr7BwExaBPNoCYsbHp3yrH03qozmV
VJb72lhPhCcHdtnZm0dBOC/0w/w4HEYcMh0elEajVyFQRCnT+CflQNWGcFcsHjyHPVGUW21MiHSL
BAnnrbSpnHmK+BKlZ2sh3fi6qctfZfZo4Exc7WwpIpf+xjcC48P5KE8TY1vFmlKcxoyaeYYNtWkB
LIuEsWSJW9RTb+yTnA8A2+Tk9odyvj3odaPO0OoKOi43Mk7zVkDMUakzavbbCKZz+4Twvf2hemog
OUrUoqnQLKIl6VZbRxCRIztVAKZ3/yn+87WV406XLGyac1fSm5AktaxCRemfby5i7GCs9zRbJLa1
0HILj3qqkiFgJ7bMt13RfSGWRAmAoTv+pZrkzx4HoIvfqtMlPnqWIwsBTiE/EniCWQMfJJcHwcos
drpFcU58e/nIdMJ9v1qbqujmAG/6kQOPJgU1JtnnvEj/8dlKNnCnqZrc1hAAqBN5YY8kVnjVFVES
rBOtsnUmSSi9h97diob6WcaxSxs8lIGATFO26uRVi1+3UPm7J0xBOT6FSoYtndQbKPT5p1T3oo8c
y/bIPt5VF46sU+23C7Xa2WV2WHPf+4XzNmfY1hc5KoYROL+UjSHJg/fBUHrGDbByl+RRKGAhIZiC
GnWJ6Bpg0sUhmtdHGHH+BNWansY+i33GkmLu7IT833vMwTui4F7O61ZxqYd8Ej6QQtkA+HNvJ64O
wUvSn7mqL0Xd/sXAWou35dLHSMWLqYn9f+kil1yuCX6Ay992DaJ0wJL2HEyvoPxaxvI+Vpzcbi/N
y1tC0zEA153VJr+Cm0NQKSNH1SKMm/TJnsLgc0tTttI/OndYpPPS66ZnmknUJqeWuX4oAeLt3hHK
weHS0Ifr415Tqd4W5t9yZ4o5VG09nrDDV/EdqdZTX87mgvJW1vgH+zuSKCXlggekVlUmQ2u/Zi2S
WDIpE0cx/DUfsEd2EutGQ5Ica31LQYZhcCdS8JB9fUQZv8+6Rgj4WB1G/Xv34ZQHEBkfRR0qdTyR
vcEROd+3bdCiBxRn/AjV7eBbQuLuxb9RAKbIB+lIEGEWkydf3VleiR1fCWORqXvLYObYyIhXKThJ
kT/r1FrC5ZBvv8x7EN5S73fL2VvNPsuhDVhyyBdxZ+R3Rb+BWIzgnjfIv1wjvyU8zGVMeY//jGxB
cgolk86ATvNMetZOHY7R4ZKxaKjJ9WMfhxOPeoM3TikX0OcPPcU08YURp2/88csAqmFDn+LWXar7
mlVyJ6CgDK0zI1thfFXI/zAZx8x3hcnq5Agy4IN7af8mgwkCVzB9DO0he/tg7z+b1aEl/z4nMVKD
OgO/udET+Wcl2HlRCShKY892xA6iZzCOL2EUpMbS1OMWlV/+2lcn27alxanmYsO3HEMqnrwoIWIR
poM9RQTZkNTkQGHJkWIEDe9wKnOTiIXl4Sp0yBoUdxmt/TejhytW8p2KNbz0fpnXvtRMsOSkehiE
AeygTrxSP5KmeC/GIO4jpRBIFRZ6nDN9jvIDDsWQV8TKFhGh7TXs2eChbpbGdVZezs9HPphfFJ8C
2fbr+1ocGCqJOu/9a/51sJhK4nW89H5L1at7A/JSALHMkk76Hhm7fY0/QCULfR8TTICy+afKuV4M
iwkbHoI1p7p83rWZAUZUq7T/a54HNakc6DgzK7korTzxN0srpqPIdAMHTZ9MOJCN5kumxWNkFnnO
NUNj/mMbEegVpQJC+T9DGVd6i6boZ3D13XdsdYLlcOTYeEUmPAvzSP7cg8O3xh6Fwvsf++1yGKZ3
/XDDJdBuZGQmtVcUW2uMMIJVsAGtIaKxGXNtSLtGAwd0jaPq0hTxqjuH14F8ptqrt9+2NaK+fw0q
/z1oyUFlZ32Pth30GDrerOIF6ekUwSSJXCy2xZtnLcEHIRFFnAhkHmooj9Ko0pvmzzHKFJSRtGJG
q/6ve+At5RDx8jTax+j1kv6eBgr6ioHYtm78esjgqxO/wQy2yTUxaA/qR5KX52Vv2Lthbo2yRNRv
Cuh60H3GpfTxKw974a4CkA6ppOlYQSG0Hoh33mwRpe+9oGyvzJt9cAQxD+WJJXbNWnZNkivod0EX
QB1c60biQeSk6g7pcpnCrGE5X1hveLpiKkf6hlc7f3HzF38AfxpOAcyeP/RZvnsh0i3tnB2RhO/O
HE4Du+QP4UWeK4c/h6yrn3zOsAyjrvW8982pimbe8dh0bwEU8Z8jNp76B7UV3Z0q7sgMC+fFLHUU
JcSUR7MG+5cuHka63SL1v9tpGI4BrPfA7wNnQNsCqACdZniZr91MWtNqnfl6eKyL5HGMb+37Mlow
JJLMrFU1dqo7EyRhHxDPKZrMgnW+peC5H3W49FK46cRxGlHyBa0SlfgSKUODsm+3mEUhCXzgP60n
1CAuouJS0Y/ARPDGFK+dzj7scaZVIB/HLIL619/kCA7HBfDNi3HvwZDUSbM+oxJbBtSSDtXxiWbs
/N7OLtdCk7gJyNUX6c7GHjiBC9rmy7pXHq7DAItyulpgZOpcf58xkgtTsNkW30LtD7FHy1mJYNqJ
G3pCMOd6ToWPyT/pWUiNb+Kfk56UmwuIcbYHvHj9hSQkmPZTbE+FEgDaxnxWvLLmuvqH5HMOQi7x
eRZMf3ZuQ9ISq5v8+k3poLlhvATNTIHTYdnhokhsO0VxIdpGjVLCNkda+wDK7q3H0pxt/JddiQ2Z
nQcnSXuaIgcsQ33ETsDpujkJzVoUE04gk55g7QagAhZQTgKc9fliFO0Bp6CRtDomXdsUmRi6zOF4
2HLZP3IFOtqEVPE7S73fGHQmLmRQ/SF6PhIgYJT9C/cbjsqMuKymRidMwO+euYZQ1nZaGUWouMg4
CbQddcfmtEmCWg14Tp/r1d32NEUNV4cgUr5WFy9DhPVcC5h9cB75tJr9OGPOJBmDlTsr0khAiiN2
jT9FP4LfvjcpVJmO0p4+iximjcovAfhVt54B69oHjXrqydHPYlY+u/kVxLtQ7IlugDSj1eV5dM6t
iVUYrHby79k1/g41jIZUpGH6LoiDZGq499hOHIsShYLGItU/6IGbs67ZNP9aV2uglrZiC/sJSg8v
FSGf4Q43uAyzjN/RsS6jADhwMj1T9B6vpDAzz0FecVnQpTmzrjXRpmZFvVKHxbaEQY89F+bnqIEv
yJMHIHUsUqQ+QjEBZCIOjPeFZS28DzA6qEpS4HCi8HVGId/bZ7iFkAaFsn1l1XMKPf45A1vuHIu3
5luKsr48DiN6KIQvvp94FGb/RYlpArDS5Jv0WZgzcGG0J3V63xLSY/8GMyTefQ73u87nN08DclQm
lhErRS2F6cDni0xaYs51wqoDszsUSpXu/LSTlo9wjfCfhZpr6MKDvzT1CY21rIvsjKJvAQlenaXE
TlkNLRAkMZcYjCn1M4FxCD5gINj9uZWA90Q04QlIU8WAki2HVxYtGdffCwhEK85kkKwpnc4oeEHA
Ddi/AQlUjEG/3cVhcoT3RzMvW47laCREQFYGr+qXs8IsNQ+45NgqcRKXjahSrjTFgZI7Ojjlyei/
b0TKBamzreTPC4FRjdqw3N02Jz77/ArDJIjrOZwlq8Yk4lg0vQzU+wkfc7x2wL9AnPGNngpf33LH
qIBWSb4yo5Y0qRGr3vPwqOaKanhEykTDMaPv37Gmu9ZUohBegfJMUzROMF03nxxVqEHcZPS7FQwv
yWDt7QtLOtMp4OpVrbFkRRZq8wWLkusmLS4gW0VzEBLW+Ku7njxgUqxNJBNZSSYFriOIj44dUOpm
nj0k/D5RIn1raqHVy1yexY8zZj3yU1IN+3/w56V0h2/D1AJAPFtJpLtwWaiJ9zfhkoVlJGPpyvuz
MfqtKee8qkJuU0h/rsYFQNPk6bhZmYwkCRezcGC7hV3g2A0JvTYOGYM2H0lIcfOs6+olZxyyHmSm
LGiClg1isTTW8A1mUQ52WLUd0Q0QRAGCv6TfQP3Vam+to0T1wUGCqfoymP+5IrXCPC4L+Ge4n1Dh
Jhr6Sz0qWixPUnMyhwyQ4Kll2F50jVPOS4V7jzG5UFp9Wd/WlxNAi3hNyEE/0wxavWJA601jmENz
7ptmsEQFkKJ7ks9rLt7sp/AAFOe08On4cCh88O2IbhN57xlLWZFtbaBSk+7h8BO8RHkbWk2e+Y26
52PRXtC+suKbx388loBKFbaRro65XuwXpJS5mr71avmxudgkTYzwoTAP1O4QNFp6zM60YH/cBTNZ
v8c/ti4JRgbo7Z6+7cfGi8BDSGmkPFHeLdxQ7QSAZbrLbRV4KEI1JiladuWe6sJxOebX/vLJzbWC
OtL8IC99OcxP4AxHMdz9IsjmITNgvdUkpHuEMDvPlJJ2mta7zvxzuKfKvZlZdmEPdSsupfgRUlu1
8hBblvhaodBAzUHLG3lKHA+Mgkql1q30zbNW6hBWda9NrF8Jky0QrBHj9b2lW2TMJevzqHHBkr6G
2I1uIY/CrAffI/QBSZRLFS0RdZl+x+hRLO7DavZxvSzI5Ib6kpezMJx6GXnAcSDtMsJWaRS7bNtn
M/akXTtX7mEIY76GqkK9arbBbGg8qV53FIAzCGvv7IXVwBiwJPyA5Xp8ZTW3EipRzNsGJYlyVMT6
ADv3KpdCOqKzujhJnOpW5m4S8RDdI3iVbPrpz+Fkzen2OBf259X0PEjBsaxHNcqiShf5vfpvlb3x
7HSMRWClf2P8GWWVxUOFiN5zJZW2jc+n6RYA5uZSmUnMCh2xEKTACHcCIUgtzBhkG7dHp2hfQWUc
GRUjhzYIMruXhZmVMEGiXTqpOkajkCqhwxMZtjaDyMMmdWGxRKxnwKCJl8a9npZlvD+G2moZA1Od
4d6rpZMkTeTIQX6+gjiXt0/+QwP4b1/kPOhKolAlVY4Xh+WgHblT4q2bq4vBjL675ZidDcKkoH63
xTG8sLafJXJIJFQg+SJzSC5LWvBnqvlR45gEYuSv2FsVD+J5riQ2tBTwjpkpGNDyy9jL3ua+IMHj
bRGONEsm6F1ExlR3vF5H/zkn/zDNm6V6I7cwDvU8emER+K0ssCncT+/9tt6N0liAqo1FugrljQan
5G1ZvhP6O5PVrVfYfaZ44mUwHts/ihJsWtQm/SljBBEgh3ohpJVNpaLl6fEqFHXadXuaG/8gOdYN
8CtT39K7yF6DV6gbZkV8Hp0XQqajbXzrDZyxUyYijaHOtyWtuKZuoAnWn9lqQq1clYSA4RDdozIh
ZLO80wFNDCQ6REc9ymnvLi48KDBC2zjOmDamLOzZ2wROQbM+K+2D0zAz1mCbXM6ffVLaT5ku/pjX
M8nAQr1yg3JTOADBBAFnwpZ6WaNxMJGkWRrS3HgHK4z4/6AOoOlwD4uA19VFymDQrGsDApQUqozm
f2glYjEldOjdCljlb4X/KHrrvFMjNt2vckMgiqAen3rIKgrvSspk4sC/mBaVgSztN8+VdgIUCr1G
syKM7Nn92/Pc+xXYH3vKa+zRitZlCR9ziLvKjhN3sV+NI4fLK+fAy1D91qlrn7W4Mk8TKTsRA9mI
s14HmT1SCpVGOpKpSlv7ysPdaqdR/U+JoOfDsZz0S3HH5Da8cvra4fCP7xA5J5V/bf8I3V2gLTsp
RmIxkfzkNgg+vrUyYRtr9AJ5LggbnfsB6Faj9D8Pn8wQPvdBTGjc0aNZO66VVnrCIgBu15surOyf
p46rhUlibHwVp2sNq8JNXGn48Fvoi2myTXtpGjOBDn1e8Jj2fu10U66pc+suTS+Sb4OTfEvE6F1A
kOsGqkiTq/EHU4VwgFGXnCa2yIRclQY0bsIf1FHDcBwqP8gObpNLGQvvAsvy6HuJHdd8FTXgT9ZP
fbFwMSitmUq4ACIaGoQSqnfRtAVzsDz6k3hSPcUr+izMY7e03QVbxqw6hTvJpw2Euk0uAEsYkV4/
MvjwZmBI5qr777guN0bDkvKAC7DNmOqsd1+iVwaMF37HpCcgtCpGXR0P/XJkI0jEZXy0NtOa8gd8
/bPGRXbdCoFAyACfI+kUnE302acvudXGLETQVGH6iq0KbLTFr1AouWdqgKLdV3G8UJWaWbOPzpD/
/ZBlRbYhEFzSoKvZgmVT0daTJMxCcipHFV7xuijJj01+qhJalGxcQGBexuTV9qKuMCeCyqp0qXFt
sekrkWn2cyl/eNpdEIgsNlnuzvBhnW126sZYFN7geCkcEd1vqmxyQGdyY+7OI5CZ9BNz6trfixlZ
z6qnWtbMYk6JGy2WYbSWcyZr4CuCj14IBMmtCtffYO8cT/aRavfb0Q+6HgOoj3DIuH6m5xsKqfCa
oz7lXUKcI7YwVDWV6CQY9TUQeXV+9C8XsPTRbDCIOtjf7bqbfS43Felp2uy2t+0ueS96+TGtfg2Q
QM2P5EU9skKl5oeblYXnzkayG1DYXBmhMgBd4ns9FPuiQ/5T3gkWjKhP2QyUlV2CPp7FAIIs/pQ8
qsg0fOdR+amPOT/2IbuCpn4jD1Kil/Gl0XZkU2vUeJ5gYnDS12YflP3lPdf1m10flbfqcSTBA35u
Zw3d2RrffWgtarBUniREUGB5O89GXnW5ZPwtoFuHhgtym6b4zF77A7niIN/brMbw0Lw/XoAxgMqv
RSlv8VKeeFbRTHlY+Yq9/eu0i82V+S1IBm0TqhrL2CcdXZZX2yYSOMRBWWm6wShUZCl2+9VULBvN
Y8lWfxD7Lai/+pNb2N91UjgJ+gO4GywsKRpai1I46oOi22wjnvQF3As8xpbzGYE8K4Vo1xS3EOUe
zn5Xt2aMkZatsE0604Hj7Lg82RJOmEoPv+8Wx8l0Exj/5dvXvSUGBRKhRHWoO96w5hpq2hcjeZFh
Cdc+UIXja8JRq1kcXFUXTAlCJu/I8ZIbzLNalZ+9JivYWSApJS4qvLLLVIclfD96JSZjL5RHUqnd
X2kbHvc7uIBsHXleAmEJD2GRuaSxWioR+82LtC1wvzthyVfj10Qk3LPcikhxh8gnsgaU14Oa8x12
nXQZcgLytRtOl6cdRsNMYocBKpN7Hkw0Ss9f9SjUmCnLgOGmIRB6EZ6xu9/qkG/JOUjUrMw60jsS
w+dkgrC37Ayw5Nm/JwTQfWSn2KWN9wm4wawsa0mTbkPNyzzl9H49kFkoZoq59mfVwlYGduL/amC/
5tKAx/97F/8UsqXGnVjWO7mlqJEzcWXhEi25/TwHKyvk0Fx7w7pgvaAm5TOGQ91n45eDhUGfedSu
Pi6grBBykT9/V9AJqDsn1/+df993+RsWS4r125BPmW9XUkaWzK2150ozkcugwFVzL6OcAaySj6IW
rVu2b0o58pkNpPfjaFuUIgtUrCPfdu4gbKz1/e7zYvQpLN63NbRduZc09hfW+P1ZwSHLZm+JLDyP
3kYEgT317oGq8OMmylySmgTVdz4Iezz2oTUW7u1G/imSIsoldUjfLz8kiokXYS8y+kWiC7vaxxE0
jQYuBH1K6pQU/t01hs2baAIyBmjF/F6zUTTY8EjILpTAcR/TwqxKO/rUsYXUGYQAvHYEWp4Q/yvE
nmwA0Eilp4XeswLRjzhCjirPBUo9HmWT0G43WSSljLcc1HGe2p1dQecZVQcR0oGeAuMiTxwUKVo9
FKifRZP27qNx9Njwusi20XkSDlAH1LDGeQRoz7JU8I1XwRG6PDBMyZoy8ZUlY0WsAZMjha78Ikfj
suYRJrT+WJkMNZPR9Ls/kmSO+95teVyiIH2N8MvfOiOtJNv//BbYjnLwdY4FJRvIq44T4N/Az8zT
V3iNRXj3KOcJTiBAGBDvbmGv8+Xc9q6IGPPYFFKtQW66RdsAtKwE99mDf6YI9xpbfTXNRUwx+k2P
ixl+yfe+jLeF0nQESn5+8eIjVhaMyOIcwuBDLlifoEWiSLkOStBCOCnNa+JcPRnwyRpzc2Tf3+DJ
K+7K3afK6/AGhLg53cl+epig92YlkXi5h1I9RxDZU9KtnyugZbOirUITcuGuRsjxviQV0NiVyDVW
O55juk866tMO2D/rRkZ+Y44HErWfKByIqqwJDlv3oAiwePf6OyrqRWM1U8rhbGnkUMkYFiG61qtB
kh51D2ZKkV2n0LByqpFthX+lRVEtnocVE41EqhP0c31BQK/kYnDqLwtj7xQdjjSMm3yqX+cRzwKx
WuJcCRyTdNeE8/zKAHQ1g2brxcm3mW25pGTRFzi8v6IW/QLpOTSwtXI2lkPt3aQzR9nXHhOu8dkY
nMyoMkJhzYQ7GOSV8GPqpXVmb61vu3ANLM8BgUdOZzWh78JSUaIVy25I8aZ8mkUkONCzaeooy5nB
I0F7F829DH219U6tougalxN6SF4g+LbWqKrl5nJuCUYq6j85DnnUxB6VfKa260PryYiEgIP33ldZ
tsSmIh4QkYvqhwak5uLywsvWN/HQ851lFotCgsjxqS7EAVCjy+KjJug9rjFqmY9Op3xzPz3Wzzel
+GHxJAeuBpb0JmyHi4JsEp+Fr+Csdl4QskbFh0faOJ+xGuL+uWI7k+BDAVeHAyfWV+4GWPETb/78
vj1U+fOfEtCSquIw4iViOusq6aJSQPoL6X2+tRpyVmn3clJg9R2leYXF3Wg9LGcfcTYyHNf4ze/C
bfto0PB/CqDmPpaYlxC5LFdevLfOgwZC9s2lfUVYgCmFLdNYFoJ2IeyxiOWPTB+LRweaPIj4XxhM
l2R2udkt6dAaS/j2uoIy6DqO+L2H3HEgTg0CyWQV0gJ07wYeenkSpxxDybhb5lRV2X6gJCdhF4Hz
GixIl2Ub4pwTHxBSSiVeqEdYMnDeeqSfKV4DIbs3+Ei1/5jYu1FB7NVuhOUxhGSPXxGhHmnMRw+0
PA7chvaMWe3BgQnFxBVsm+4IQBs2rlYlVwpdPQnI+XHDWPreS7sMN+uDWOj6kGyjfvqpHuVMe6mW
sxgF7JwE+ZehTFiyPZLZygk4ctoi9K7IcW3sbgep++dufEXoMW2YhVwG2EQiqAzxapuMJXfIvYik
UsYEMZHRxGBqXJJRA112PfaWINWziS2z+zV/Hsth/Xj5C+Lg1ftNBYRXuybUSbISu9vUboLPEVh3
toLCm6zpMkSTqbjx46SwVgfvovoVJUfGFnHA+VwBo0s+j19nFsPvTOuRtcsrwC1sILaR7wNdY4g8
DXOE2hI3SEY/8q6yy10D5+Mx4miVqjQMiiGWnIHohkqKhKvdc9DShscOmd9UFk8k6sBOjjAot7Z8
rUg9p9zvn0ZyIhhho9bsj2Fn05fyp8MNwvMgQPcDdVgBjfTcRrQK4w/vSC29PqpcjEDQV9EEsHLP
dS4FuAGe/mgIRlM9ejAiew/oiM9NEz5TRtQaESW92hOdKwQRp/e7SNWUXr6zRSg4H1Ta5CvX2d1m
pi54LS83vRrWuU1vtsKhYS5ZH4mM0nZ75OFYD8V8CnKqOzgwKKGxU/dFDAptUw4fNgbdkYHEqL+F
bhG3m3urRmgRH+BSjIRzWVWgKvI+LDhxobRq/ewwMmf5uM1PMMYScPe5jxD7uiLLwHIelFWH3MHN
al3KnnSA5EtQAwPMsf9lhNP1EiSZvmT1cDrOiid14dSFxPBcg2EgAobdk9YNxNDdfAUwiEOs1AnZ
aMF/mGYisXLFIBqIrstVrXG7Nrt0ic5R5IG1iGWIHg4djCNveTeyzYSIYkibrQi+uw/dGLWdeUBF
aLKbYpQGm9hgI7dstPLM4x9klyPRLJkml+xXOZ/PZVGOy1khgcSDgVDrYAUgIUTh16OOpdOcXEDH
XFyW2/SfkNm4J0q/8wFAYzyNP69GteyGqMa5D4EB6FLvv320qOduiWzuYTt91r/OnrtrdPcoMA9g
71te+DO2vul6LE0hXy56oVImEz6FPNmdacz0BmHHR5u8mzQRWK2QPP796JNNjlF30/8k5VFmNAdm
r+gFXJX+Mwwof5d3FiapSkDmldolLsGjPl6NE5wu+zaVmGM8fTDJFtAWJYgYA8fFn7PEGqHUS2zz
4zjVGRmAOJEVzxQMwe8J2f9+RtgQXawEZ/r+9rrOmqqxLOPt874FEbf3r7b+XF78OAMppD9GLaLQ
NIQSjQNtnRcHUdW/n7Px83amBoccN7z7c1CF2artA9sLpzpdBUD3OHJHxIgCwmL4aCtFJn5x329N
B90owY0lEC0VrqD5oVmW6CpseEn2fUbjjYcMdefrxtIES2vrmim5k1S4G5swW51qiQL2WT4WeJNN
vjHBeCYbEazv5edQo7zq+OVPger07eln2Ep3cg6f+FT75QWKCtePOxBen+XunaY24RG+r3HhlSpM
qalb00Vup0UxTz0l1uOOSzOEdZWgfFhHC9otevcUdyFs+30PJtko/tkS1UW+4VGThuY1Gh4VY21d
PR7NQ2QUnLRK9O7snIHxbAnj/6KTv+U72HhO6ZN6RBpbdwsiLdp2zDX68JF1zHgDTAvVZ0OHtRUy
SqVJtgxLUk35kgcyj+D5dHb6aEBR7TlOSXPiC/rhmgK0S8qWsDK5US+SZXlRR1vfQwxDzci9CN0n
dXSlMqOd9+NCrGi88+k1ik2yRODyaZW+LIyN+zqsBdBPqCyCWZiR/d4lqbWD6u/Six3sBjPnsd1b
kq8M/53T5DMH4DWG2jNBeZaAytUrSKZ1UhtjubMbxUpsdojcqVn/gszlvaD5JRqRKXLtsJHR1YJ8
c/on1zcR03ct5Lnm8V/tLBVTKhNctFSEuIHrCvmJQptfzlKRYt1nBG09EuBGP0vgo/FVx1+hNKDT
//bE+X02g9KjlSUjCH3QVlKkxLK2awTg5GT1lMmwYfXqwGzhTm4/roc9kfZJqsykVveUNMk0uObX
aqdvAJbhqMyPK6w2p2KdKBGLtwHQNm5KyQTVCYGPYY/m2jeCFOK9AlN5QFi/a5Cl2dLoemOE3N9z
xPxfAxoRTyQmen0EMGzWFQsJpQ1cvXWb7YQOe/TEn/uXMe4drjT3G1gdFGsRYjTKxy7A8RyR+RX5
YdUJ6jqiVFc3GJLfrQv2ezYR4CiCymeYHxkDHQ/wSSCfUzppZsxURvCuOmcBiFA8zkGuYNzb3Dnl
w0MTW2lcfjQlknHQyU0X4K0L50M+m1UQT3nUmNWA7o3jnMzNEav7lVb8c5orDFYiLZ6SxwLCkmww
48idb5st5wTdN/vO7Kt502LX8yj7HY+O+E9IwBUFqDxR7JxsEgKfboisDAexp9bOaQdVHArkbK+F
A4qOP1pTScQ029vGx6BqwuM+ouTUsusGXAbpqZO5Ylyppqc7effmprYlEL/6YcqLKbL+8E7wYEyJ
PA8+dhsLV7FcoOtul2YpaDpWZjJ1WAuJvr470CZebknZPGEkb70KtLbUqFQACBLP8av/KhvBe6FE
UPM/G1G/DpRfmFS7DGFyQDskw2rUMbc3a+7slRL5ylaLjQowAsH81c18VKF3kxgp1BYo5HfEB5E7
7rWMmHRu+qQ4+M6hsdawYdjRrGuXSYRD2VEYQDMNq9XH4nJdPoINFCqWMp9aQ+nL8X3IVJWeEBsy
Pf5nD2rwrxOUuSMkXt8QZDSptf/RoM8Rf0/sC7Dw8OWCS2jyc+efnmG6aGvqniejit1IctsGSn8O
0L5mrzaAM+PvHhFfbZ2xFUKaXH+PSMAQ91EuIXEmzxAzi/wsKner93JN9M6Ci+EbT6noiq4ADrRm
2AoWuiL03FxalDrKKhd9i1H2Rab6BcApOdT5gokamJEM+zPxUKI3T3S7F3H6drY+8pDOsPeg4MTZ
h+vwjzyLLp7CDzxECvpbqYOkdrp54cND1KecSfjUrrZr8Ub2oQWBuG81mFM6ZzvbRp659i3c+Wx4
IwpsmU0EFuZC8hx7TOhWzsjf7V3Mf1g+C2qls3fDY/SGoJPeikKaQxXnK3HDsPe+qhpq+b2Afqkv
y9JE/jlir1FjXVBfihv6GzyPfhWI5V8WWC31K46IyjQaYYZtnaFdJ/mcVNDxeiD36OuIWwYsyeYp
JfLJGn8yhZUJTD3lxhvMB60SyRAz4omyOnirwjU8mVrJtN3IKebOyMqj7Lz9vQMon+Ja/a3tU5p2
qSY23eJ1yQKllzTlsGUXvm38uE0fix1YPXYpu6md+oDpYAZCcIW4mFG6FpkG87tiap3te4BhVuRo
wPs9Cz9ikVdf1rIStiaoHlC4+MQiYnHA2n5ijwFgbS8WStdt6MMoEmXspuo2XvSzLMvGgWvoCMGG
M3afA1/UeVglNKJM4UyjSiDPao0lD25d2T4S3+QNUsUaGZ0TyIJfUWCLbadPcvdaNn/gDQTFDYyP
+gX8nIXEgPoDGvtc103Sid5jB2g/b4981wxqmXmGXVMKkfz2OMDmjoxoX6ZTPeH+fOqzsVqtExFm
A916UyoEJ9JN2AwGTTv76YnJ71rHvrroswJ8g6nGeYNR9Ea5MsSsjEc16m4Fz4qAKoct8oqecFor
eBjH64P/rmCJGgz6skQLEPIcRR53XusTIrcnfUIEgda7fBxxnHXTQ6MkjQLwQDIQgU/EvPioIvLu
HCulZDA1OP98LRpWyhEUwWyOJXeCWa+ZhhBL93mzcZ3fAQOFFgdJ5w8xzWRwbMnS6UIxE/3rOjQt
Z5C5MGkBwrvHNOwEY0ZX5j3Wd8x+HSujFovnD7j56p39ha+5hoE762j56w+MQ5CvgJQCgqv+z1/U
yMWJPw//pGUTH7BtcwRiQyIqUXgZb0pPGUU1a8g+QPx619km85HjsPCqujVk5FJ6b/hJjBP9wg9p
LH/1OA8dR3r+t1ipUAXjpuaGbi0+PRian0CoDVFq/ZPm4etm194CMAV6qs7Sk7zGvQ+lYeqCKV0k
H/fBFvM5toTOYQZGlgxLtfpcLsqcn+ZdDErmnFkaVCFCEUmsiGKVLdmhDvZQbmOd9pMLWGx8Rm4U
z9SKcsssbwKkQTsCMkMb0HeOZMSZINpjFJQ15dMG1AZgyz2aEeWhhGxejWyzGJIvg8XFwahr/RDf
FAighlF3Zf8+DtAeNzeftx+x7d7YWgDqXkWTPX34uiTfXuUht/n1wcInMzTzZzuBZq3tiYHKc/7k
aS8v6PlMNy9T8Vm5Tpgok0HFFRSFl478QFC604IbJ+Z/jn53pMCOJD0rNGH6MH/AfFRohEHve0yF
zSoqIwz6+dggZaydPlDoRshuu6H5ISBPI67lisD6toydylQpymFn2sslSjPqq3HS3c9t9hlwviOv
RyEWFuz61OO6KNrwe91e4en3Mhfc3MGpzEr+OokrhxZYYINaHxp+aF2vkJpOBwr+2ouTXjxwNQc6
Rrzdtnqd4A3Uv5dbShsr2gGjngIQcXiFVvyuRdmcD4LGMYz5h6+HcBKh0faUzrTcMF4yhmIK0Su0
BBG/mSGWVbc8Mt2KdnLqM+mrYmG8cZloB3WybxvpOsVUe8wLR0usAiRMEasc6zcpJhA7/qT+POhk
M4ce8xHfOSDBbzISLvwwA7zI08/a7HtU9w3a+mKWwQQ5y3gQliieI4kb9U/U0o4jiEMbSiJkKiRb
QXAWTIbBVHKIJNUgkcc66bk2r+fU48mVQSooPkbL1CVGBB+rM2KMTu1LlcutbCjCwA3S1+uUViy3
f9WFTUAJOZz+5wUD727u56W2YLrrHQCFhiJX3fQjlW+fzrShx84TkmwHaUSlEl2kUyM2fgWT1dXl
LnZWskf3XIXkgbsgF8/2AAqzUtqfTpWYhUbQmflKHi/mARcxbe2jNpqNQVp+/G5dIr4B+sWq8xCU
qMWfDDxcBwT3RpNNC+CdNaQIQ9WmgAiEleIjd697zbskvatomnowhPxuNSXJf2cW3+HA257I0RJ9
dvE+6jWV/d9Is9LvhLfv97i5k6m9WccjbotFmCR00P2SxjmPskyDY/HelKb14B0IsMyvWd9DZoSC
tn2+T604a2G2H8IxVPoDF9IITqUvMhgtHsNcJy+VKsVrTEskyQloml6j8XfnLwCFqcOBdYrhRywX
tXynhQldk59X30IOfTXC9ZJ0YV9I7WtzmlY+FfHtvSbfofKXdvNt0XWCS4k3AiRozoL1XeMehpj1
mbo7Y14dW6hyVnUjVk76XLsR8Y0SnEA8+MalrZXrLYIs4JjGQ/Ch2PlhbkUXQOdw3EPhg0u8Bi8c
3g9QOD1iJ2ogk9V6PCAA7hIvmdlipADYdyk07PN7anIa+dOliRazby28KDClESBuudvQqsIc3tHf
Ba1crpFU4BgXQn0j9Toa+IF+BOX/jR0jRSTyUWMEiZBqu/8K3vNA8npDUoD3PELeI3qMmD0HM3Nv
n3ZXRsZJ8Z2z6k5IOQvgwi9jo7rt0oG3oUt856Qx547oLIXKJl3Z3BzfUQIkTHTtB5nlNQyJkJTP
LnS3MP7wkVT3tTeM/enA/mmURrUQdOmG+fwUGOV8W2j1rFWeYYC4mjfd7/29MXlJzk7RQJq7VaTp
5qAPg37kNcvRqAApaDhTeWVHD9LlZiRzW8oOi/Gr8bL+a+CX0qi1tpcyUr+Uxo0lU5imomjpA6XS
XjdXJiSwd1QG23FArXDK2oB7Sy3PrejfrXq4kFG/DGA3IED6jRlOkLus1tHlnzOF0rdngma/2fNd
8b9LV6j2IAm99Ddo07yeZbuD+Ot3DHs/0YS8h2u5rHHyHDbrhHPEWK4ZBooHd5uirXlmGPr7ghS2
dghmy9FugSN4FWBODDEAs/1GuknchkjdeNHHApbBJFH6MxJirJH/y/RW3QvJvQr+BJcRoj7FDtum
SLSe2BarykjGl2pmWQ/VOR2xVXJ3df2YyZsxQKZrWUELT0Q7kaxIWAolmjPubsfr3wLPdT8mjfOZ
z/BY5qx1J2lGJ5KFsp4SaRhxiOINm8ESheJNQpMUhxdV3MALe3tVnKVDrGjweYx5wIxUuKlVO82w
V/S22/cYLkPkigS/Bb9KMM6gkO/8jC69trqFeeQ8rlukC1mmGc00IQnjgiEbWq8O3Ysl81ocF1ZD
lkXJ1lAUf0FpqMoxw/FqIXI7NKctvt2gW32PUrBt+gi3uLAMivXC89wliuSYeze6US0p84SWBq9G
ag+fUHwYOq7pfP5qMueJozvr+xRNvGzG3MgHbvoTHVXPVSkv1Quv8tKet0jqnoyJfxcFAU12/xRs
Bd+blogXdG5Gp1KXGeM/cVpcypoTUCdK812MCdZF4CNQ8p1lvAlimaTHovAwqFTPGBIas1DRMeKp
7+ieHtvEc8lvBcEEW9eTropBk9vX7MgoARytjANFBlU4LNVUoHwZ+xjZPsxlZAETQDMrfAh5ySjg
96qG6GCt5y3wIr8r780prkerPGEJuL7FyCTNgCMnorl++d3FI7eDg5dXTVHXnznyY55BTrY8w/ZQ
Rd90JgkFEzprmDLPPEyJyNNiksnvtYc0XBBtaXWOGB3vK3Iuia+e+2wInZoWFdVogwy2lQy6fZ/p
KUvFtq5mKR6fsgAD8WXq4/McqzymWEO12kmxK+xJA8/Jn/LDY5YxMJT/SdiLFn+0t2AbMgvz+eRo
aCKasfdx5EJ1nhJVK/50j2CRZQardXLyaJTs8urBz96CpBAICdFVCZ67F+3G8jwDsexu5CGS0GAr
+6xIj+heDnApf3N/cwXVOMal2pef3sLs1wPCxQBTawefAJvMvf9gHqFx2ex2iKVAKkdEipUabN5F
YvjxQ4jQqfiQnZC/4gnCRsmADQAzGiGo+EKUNNVBK6YgJsvqw2Cb+9frDb57QPvTPqa6e2DS5rYL
/tEY7MNN3nl3NGv/yV5/QQHvHZg62xG8hlYfl3fXQO9aDJTX4vWei3vIrqaHxkFUCjOcPDcOuhLy
MUHlHSFsRUe+NEQzSO+HVTog7tWkWUeqWYcVH3N0Z3G7RiH6PaJRHzJoJrwAhpRVmn3HP1x8DnWr
bIfeJ2O7dSgEs5UJadk/DVrxgI6ZGHZpe70qvZx4BeZOBLuXip3VframSiJKhngXGJXADorH7FoR
q7naaUxSRd+zzQ7DAewo0l7X2umr+iZieMZMShC3LYiTugGrSOgClgaJnCiBc35qTxV9kfkQf7o/
/AhPQRpBKmwj/U0tXe1ynkbqE3b5rsFfXOH7a1A/mPlw/N742ZpwfAQxwwWk2yyMkrU1+Pnkx62H
wEJEIo9YR3G4ZWpOB6lfm7vGhWIYdQDY0aeAZLwOiMZbEIMXlFqoHI07GjxE+sJEvUyND/+vvilK
vNvrKPuSjhvToWmMP38P00j0intGeF4JmuNESKKbvZSpU9dYsR6lV11CoAa5iZmVE0ElE7PtxBrN
8WVaPE+mQNSQGxVEn3C91+JG18Vg82AdfEp07xP5dZiC8EFrsYwqFle+WSVFOl4xo2SSo1STxX1W
me+qOKTSRuOMsTxz5jBORX1Clq2Un/gxHlepHWjhO4K1A76XE5vTV5evLuZOKhrwkNYQczfDIfMd
geMxiEoHOqateG0dLWcK4SxtvJ5oA2aOffE6CMZ7lEv5kuN5tspKmyauwKGnHD8tIZi75YiPjzf3
GMM8Gv0YJEhJpUFcxL0lv1TPiOhm250u1aNfmlX4C1K3etiZtGbzB8tS4kk9SZsiZZPrGcd9ptMT
EH4VcPaa7JBncaTplUkxE78g40VoBs1T37nllThZucj3qgjRwjYaRZIB5nEtsMqUS0tHtpUQBXx+
edQTai8UmWVnZcyt87mYCW6oN8X/4RjCt3BD+Te+VrO9bfqvdkjSBQozsHm1ZSBOdTpOLeWEysQp
imktslFa65PxRz1JfiCwdRb0p0FFU5nimo+DplOLDILrswEbdx48lD6N6ppBUY1L0AoSWn/dJIdp
Hs0GstET5a9UIP0GMP57Em/TVkGnQT95jOPD7mmp1KLOUsDTeX80fH6Azw10EwJamIkWU808/QoA
qOjRTwK0M5LQaR2hhK+xL8XCXpATZ8H66WDa5YJnhOFXf0Bxf3GNvmtWidOjsiaq6Nr93P7IM81w
Rf6NHjT5BIL01zg4wItHHnxex+3ZIp31V1ywWgPhMMGJiYhuwkhfFjsXeu4r5cYACKZdAOkM2OQc
0QqoQRMOYWoyeFCLd9Dnn8NOY8Rm0x0tSNWhBFl5GHgNcr7mMoB/5sgyFH8JRdc7es5MbGPcAgcZ
jsdp93thXJS3l8r3y7Iph1NLwbhFeM1qZdWIgBlZzkS7Vfi37w9v0N0qFmg3ziaMVEq5q7p4hcIL
2NMxMj3dcHVaFHsLSaNwE57PyWKnE0Aq3clAHhth0HgYY5j83xerJEcE78FErDFUX9Zasabyt5Mw
nGjfJS4aM3WJFFMtTWollc4jbeVHhgDLAEJRPuVlNHM7Y8W94uI6WzpXrEdHs8m1q+izLaLk5TW9
0/7nWzxk5t7p3OVyKwhSXgQBu/oW7Zjvub1ioD3lRpRNr4gPpfPPIfrVCbrq9G7Fg7DWMZ6d0RMu
goZbecrpv/SNPKRkuhRmdx5zsDMYfgwMBmLC/zngvmbj71unyIh6pALYzq/0gb/J1mfrIj80dj7A
NCVI3HePiLAzAJllKALMPRZUEadqgcFfKa40D6+nPNoEGDk1it0oLmtynU7DMHEeQe1es3jWZPpm
bEiImB9e3NJ+e8IM0OWZdP7JCf0WyMCY2WMaytGtTNdsYv2ftl1dquYR4gEBPSQORz9ZBnVp/K0d
+s09tkY21V8vjzXwx7Fgn19jXbALOheiXxso+U8PQ1sitpebw8NjFzIaX9Xzjc8LBP3iRoY5bomo
6RN2eeaQuYfbis8h+Sptab+w16CHqFmFxd/iJLBIy0NTKEXv14ddwjJ8ZPrPeF6mkddDfcHP2Owc
sQC0v+DR0h3chTT2p8GprG16TQysgbmO3zHj7Uujqw1WyMWDAaeesizAkrwtA4Jvwe+I+7bgys+l
/Xu19CUWZa5XJMQSAbYvZ6DZ+IkSoWHiiQEaqLF7r4CM3M/imboL17EoyTbnZM2z88Slqx2VdtSE
sjgXU02/bEZBq4ojWSCx2/u04gUdNuwWzPbDJKYfjLOWh8+qsZD6BS0Lo+Q+RrK1M088iYUxkMX8
6DSrmRP7lIXIDJfgAeGJiaEnsMBSBUFq/Trpj7u9bvammLcUtP1e0y8b7Rzk3FMFsZqueS1xjVN8
htrvwnsyOeHCjUstVeV0aMRHrG6PjOwsEeDae3+jHkKrT2ybj3Ywo82sjA5sEOTg8kAvdjA30hgf
YwzZa3f8MDsug7k9pFdcRUkt3V27YeVaE4ggeN197MF+ccbiyjWoInMXqQkXrz4ztErshdNK6zJU
wo3TVm3xyti8pqcHR+dmNaBMdfgw6Rxd6LOxo1IeZ31/Zbsrp/DbyvAV6SVaP2dfKhBIcaEyaxIK
50tteKe1Xjrkb5SSGUuvdtssahSGeqwrHgDGSOFMbME6+kahT5KCohtPAE86bROif/zIR1kRjXfb
ozOSFuMdrrU4NeA/gqGcSWzyK21L/aHbPDdninfJD6gycgyRGX+5Vd2gScarRMe8ZsIBW0FgfmXa
+K2oJRf+I3hNLbIlm0nFuOvZWh38YjNlfiN6mSurEBMzSjkcWanh8woGGgdlq9SGjlyDlQFgeTfX
/ykDjzs5M128vURgYoD8PJfWyKjdHK0a48spq5+PfBtCKqnwm9Bj1PisiWp274ZEs9MRTOsL7aP9
r1CKh84d5HI4TcFYBxp7cGwPLc5coO1YRshznQ4TwZyH4gGKlDKhIMaovZvV0/CTigJhOXy0TBcU
LEKFwTVnp6JTpYnTdHu7MXQUKhTrczy+rEwPUwKzeuoyNvu9Ims0JvfPEoteIVznDXZbFd6oswI0
gueyZmxtDG30xvkcfmFi3cIhaa13IQa9oQghnyt3HP9OVhHvvUJTSQY1uzBKgCdaOGIdXOkaISKi
owZqIn+m/vkyhL+UqpoAjvm9D47v+VLWsOWARQNSjHthKKNu1J+3jLZplxd62HNypdsajqbrFxEt
C+WyYEyqrAAGovep9AGfqN4BhF5DUmkwrPs855cLRMVOUKt68KBlbjmAoSNxgQGDSuRBXEI4Z0ua
U/B9owdBC9GZVLsUX2iI9zxuMVbAjTouRgOM9fAY7YLf4JherTAHiuLIRkzrxwbxg9fk7XXYaSYx
rsJaCFIu4hxW7usCr4bDYQuLrVouqDtnro8ourGSX5CfJXDomrRruKAykuUReH5J3VLN750DU4s1
g19o4CbV/Fb0PmB+s4Txhi1PMrySwkBz4mjGWXvo4JiOfr5Ld91tWGCec2CrlkQnvEgDvf63bWRo
7djKiesYElt0P3BoeGSV1qTMJ3RpxhuW4PhEY0LbT37/Wapdht3VGQBqGe22DP9JKEG+aEwno0sh
+OUT5EtMQvKhgzZVxPyXjq277psJx69gJEAHSTGHXaskJ/NqzwKV5YbcRQ9PhYWjja+IasEVgSRw
z8GUli6ZfT5oSU0JNOXnaxRiFhiBnP/MGDE3JkI7CgYkggSSfMJQYsxNNJPCBzsq0ZmbBddhQwwA
rQkALDjjEyJ3WozZ/LWOLNFtJSOy2m38JP1IB7VVidsXCtZcZ5YDRw+M2Hyr0FXE3GyI3ZdD1m6/
3igDddDJAWqg3d0/e4EL6fTmnj/eTgoGNXLtu3AmEPKLVlZJVKg5zJQ4C6hun49NlBNo0cx2TJh7
SAd11zZBn6VzCaddRJSraVVASOf06nSa51M8ZlXFePzeOR7aS2hMvIbNt/7dJfmUGj3oxAMa6l0I
MShzqfXny0ex+pveC3RBT5r2O1hJnx9hesXIVsk0RnW4MqZ+cFFlyvapvTHfOt/Sl7H1u+GLh0OP
xwbK6ixImlGJ+gYcUFG7Z1GfD62+fD2FVDxnOn/fGkgy/drm3oLyfXVHIkgRk4HYEPDCDh02Y9oW
77941oAR/+EgaCel0i0BvVjWyOQXmdhyuoRUhh0apN8pTEehxG7wrC2Ub2v7fXEhq/N4x9KPfzoh
Kqkl9x0b/+zvsWczu3b23NAzegiEuvIcmAoDCxhggacBBlgnfPC97XNdd8wHuMRbWJZtOjP6EVHq
GlzQhC3flEfNQiEBBERgzQqvbaQrO5rprT+ho6gcMHb6FDliJg/x3XavOvb9oBpqXGB4mvZ3lnBE
ZeDYvbm3miXDFMAGj7gdw0yNG9LjNhS02OSVB6dG2TDjyOGKoYy85sfIw/fs8A0ZVEzHUpbXi+7T
Ez7BEKt5srd7j6iovHRskCFH4LOuNJ3rrW/YmNgYT1xdy0dx/3YEQhgByqk7pd5Ey4YTy874FNFa
76SxM2lonVJW966GjhIQPa7EkVUfa+QM+Gc09mlK4ZW7EaLXmQdj0mp//eoXL9zGwsxiGx0QBooZ
ZYrko4brjNSw3MV+Y64rWbncgoRMGr0F1KaMgF9CxOOkS64BbTp7uLF/GOJ9cSHIBb7T7jWrmbyv
jPqwosmj/wIQjjh5+mLY+M+QKXwrKOaxZ5p05WrELaY5BRoSeZPhWRGjBTfpsVBvb4kvzqmmhoRC
qfvAvo+EdHfVT6jE8IJZ+rMvN9xgRoDSR/QUbpTwpj/PnPGu/IbUceYX+1Mx0WW3Hdr0wub/UZEL
GM8iTN/j+l3lbLHkvIpl+6X6/4lk4lVRYl9dPShR2vKQXExvxzL029adg1WWwm6+dfEVvj0dM25m
UEmNB+ycqfgErRplY4Lski5Zw/IOJ/EQ/l4wS6cGmCVBspIwq7X+seLuS64Ccl34W+2sAKzN0EwL
bvjuNiFUXLjpHAsZT5ivJekqmuoJ1YUZvg+AiEOaJsYZA3LXg+F9cRC76IzSypyU3dZwZDy55Yxr
LUtgEeI/lTBKWLHjjoKu9Laq/yIcGQZ8v0XxzRWFVo7Y+hzNHIDfPNbSFf1BGDTdpzgDT1daw2Vr
ZK5pTP8zTJYrvL752j2l11G5o6+D2FUula1hzXsnaYrp0kr2lD1gSJmeEw+wgBeq7f6HtMpbJUmW
ry6OcfydTlFc+2QwtEDHVhiHCd04hOatK74sx2iYUTnKhUeJKd+sUB7hLanUB9lTu90MIXDn4Sdz
NnGzyoqa3Ur3kc339B2YT8b13cdo8BWZ8xG2VPz4WbuGJPro2rRMdeBpqgA0tmrAdMEcVda6qhFg
MGnAVFPJ7Y7CzO9Ry2f0gPE7K44o912zRZrjGZF5mJgwLHuP/5onvAQ9nniu3T3hnX3B/JnYw8l7
xG7bmNQ5bYTVQNvYQaAdrGeV6VE7gKBAXU3Fzu4gtQX9bDYpDT8aX1gF4Qh1V6YvhJAB9JEiljHO
APnvXRhC3Jk9v1NyghT8Y/1ztjZo3mcPu62vRRnP61qKgxtzTu3c19vHc7TyqFo+d+4sxKdcFcYs
yBJRVAPF1BdJALbo88kqI93aXXmU5gzbFXKILE76BmiDn52OotF3J0ciOMR/fBiZBUdE8gW9BK5J
+eLLwPpEPu2dWVOKQ8wWT19Nn/vhSYwTDhrr6SSOm3cLzN3PN/DhRQolQz+I/ELohCplig0ZHcXg
dx96F4633ZQP8CGTDOgl+PBZQq/RlM6PbKkKAyxRGoDW2VB7htvUd3spUKQAik28ABnqGzRjotog
E3juSuKmLZAaF351lEsmxfFzBHizheY/q/xoljYa/nDc6SfoFiRgn0DIWyFxyiiUGvkSXGfeSoJh
I2tSx020TVO8euVZiIi51rN9fIcF3sj1JetKONOn8Zbwu1mDdQNrDrup0eTpwyK3QUXIqvzufdrr
a+K4AE2RzVAS43sX7mp52hMVRXIwX69FKEYZYlGpqK9xHs9mu2NeQkP33o9JxjOxsshXtO3IKElT
FltMG0MrdMp1AM+VGKSRIzx30y8S1rwx2sXGoQDt+Q1k3pOqF6kpROmhnovbEH36VMCJHhv8VeMU
YAJ6HR2+rMOQT1z4dloz7cZuoHXiJ5d0M90qlTry7dGjv32r2Rlcd64GXfMLSUbOVnyZgrn9RvQY
PqYfEZ13kYyz5PAhWeglSzrcXhGzBSGYbxRNTO8JnjJDM4nB2UvtuyBQyQLUMd12PPc7eo8/XDFH
SrOHC/v1gka2l4pjum0HSqIuEVYajd1F5qygEFxc7ojwsxRGgx6lARkZJ0SKNJ+iAlwgh4W5TYTg
UJlR56k87YKJbdc2T2PcsA6nZQSwp9kGH0lm2qVcg/pev5TFlmrS3+6UgxhGkljuf+fljX4Ie5aa
ueVKjHQgqZ9NwRZW8HlhW5Oc4PEjEVFRSJIDZdbU0VRMS2g5dPjZcSzkh3U8lnI9HSFlhpXjYCm5
TgQZ8tJ5TQRXpuBjOgrCbYJ1gxkQsKqIkc977d/INEnlB9TlR+IPM+fxx7cNIszdTcXoe1GdwMwU
L8Ezql1VQ2+S0g2+ltp8PE7fDojUOOyz5UY9lSY/45TOMig/GmrngY4R0PrAECvxIUxg0u05yOzC
Rnfvbe5rTEXpsjIfoKMj41GhIIAeP8ByQvgaJ28B8o+8ljF9oU0/jShsqxqNzxQ1qTPpc43OVKUW
gZoatmT4D0WITvDCsTuUrxQaT0f3qzTkbdkbJTZrz06MY+Z1BSvsWOGOznUy9PCkp8vpg91EjS7Z
m+cFOmVuJrdQXWQgVAgxmmtJoajJMm3FQCOi8T148Hm4AO9GGBSEUs5kbaWWuAC0HHOSrePktoXZ
unsnDFVD7kdIPFp4pgDvY1imHHmK0iIDf9B2gRLsuYYwycrIV3CqxnlIoyONxhGlxoO/zlhnMeEJ
uM+KFszZyXzXRFPorLsP5uWUcHEwdLNfNdai3TczKGrpFdd/0KT26pw01gIb6AQU5MiCIzxErnix
/FCFtCjejfId5GhtkfRjVqF/DyKXRsBDn26KPXwy+ocufbQQpej5O6pJSAYt+2EHxMaAAdKCVo1M
gfqmFHtpcTVfsvpPc1/TfNa7k8xHeQsLskx2ItKiYdmCRsh2uv4xiShicznYytxVhFpr7MDz78PA
mEzZuzVrGoyGKNJliG28q0av0MnqbGBYXWKFrADP9bMFh/y6ff0LjiyxxVNVtjNJVYkxuVN9qYAR
1dcUpWnQOGznPAMIsgKlV8/Pl9jQfAWIv/sGqnFy/ch87f9ALXCSLnksmeMj25orhg7aDnNNzxDx
lfO695Cj8Ys6nf4WbeDl37mB65dGTrlD4K0357HOxRbOA09lILNX/rWj1pA3bngOalFmc3EXBDHL
zQccl4pwmAb5f4JhEJsXbkxk7gZXjQKXPfUH2SVcxP9dd//lDfs4B/eS/4psy1oy/ITLlILOUbsG
l7/f5WBbKAbURYWABUKYELBCqysbmokqOM+wdUh2+2nryISlBvaE0SK5MHf/rLFI6x43tnQ/IUvE
xcoeht00QHHWEddjPaFVqbLpo6YPW5+giJhX2kk8syt4rThvp0oHNvfh3LEQxn+74b+qBnt1X9oA
2pA8iHxsdj5Cqw0NaW6jkGcwqbKzR4JPETLTARRktx7i+5wSgONDF8SGrJuH8Qp7ApM8LRAa3426
VDZPicZ20ketcgZ3OyZhhknbLt6bbCCqojv1qihPDenttFHlaj/vGHg3/FOQ3MzBLY3LTessa1vp
FmVZcOz9FfLnTaNAVsVMFLJpwJO0qyvwWu2v05Ql5peKjOPDLX/6YlbtfI5jRGMg/1nls4IDJKHs
+pGA4zvKcNdfceiYSE0uHziQmwK1kG93uJWOaRnGdYYLvwlg5JdOJPEVrFYL7EnYqRBtvBGTw9r2
R//2hE9c17CBO9MxZhhh2PBZooBFEbkLZeP5+Wap6aIkd5gttEhLDlugUKqRrexlzgq5/dGtm8LQ
Hx18U9Fq6UeTyKJge84APUJjIbxkrSq9z8rEerfnMRxA46M88sO/9p/aafAk0dftCxBPhpFCRVpr
/l2YpSE3AWQ2HqBLgbijdABuPvmoYMCDN8U/T/Kw2rGH0RlJxuHG6uvvOl2wBFpB7qidHJlf5L9E
jnOv7vV2JZkcpPXoxQOiOZRnbYr1WQnXwtvzlts/sUhqn5Ic0+70ZNYqPlCa4JomJRs1i9zFr+5g
lKqVYpgj3C2RN/6S6wNAttOw5h8XyK6fJRqs+sse7BEafK7nsgzqcJaHE0G2CpcbjluaYXs3G4xb
Vvdy3LdZcQODngy+X8gTBaINcCRpK/kDoM1kHD01Wo5k/RdTWoOuu1ariBTeDLxAVSSaTNzzw5G/
aOG9Q2fMNWWcXP9pOt0TRFEdWwAg+4VjRb8GYG1YPP/EJy6YNoQT88U+jtUcVQM1Ymor3t+s7JaG
cK8T+4C0nAG9E6Sbv+qAD0Y9S0gCA56fOTYFy3jq/Ll1HIpyFwr+GxXdBNnsWwykPPM52ZU9C478
6bq7PjoL82tqJOQvZZFer5fiLLy0LY/t2NBZNszqaZOJ5KBdfss+er1PCI/vfs59pL5GWGPlCgQo
4xr2fz+la3Bi+DAj/ANapdSUoNaMGTJI0kSSOLRCZutqcOWPGBzaa2YwOlpIq+AAwH+iSUQHsywE
3IdYTR+owlN63fsMwwReW54nfAP+jWdq9bdCSGL+i7mjgTWZGUXWTiqAjPbriMycdZh7cxxIrqHN
vSQE51h5X+4OExy0EZfjXN5KKFfz1QWQxlUCmDLwTaYi11zONfU8k1A05vVj3rY9a9XOoW4Cgrdk
yXVaANEBlDmPt8AsdTO+Mkm/TzxeVmIa/UnTgrQ3v9iFVa2LhPzBDeSlFtWeRWxP8nXdMZbpwd4B
8x5z8yPypwAbmYYOLiHVsB5MdwtWHtWncs0NZ5qTG6JMlnVCfhYc0/qZmRJHqchhY1iQtEX2OgQw
M20QYZ8gmVzw+R6IMw76KC7g1BK/kPyedYjBeAfMJ3qafUh7QLs70pyW5lRPQgSaLGCujADeydG4
Y8AF1mx00598f4dg/607X7tjYBne3SFnjSOOgfWBiSIStNOyXV3R6FReHe5BEYUiFfTYWNIn4Eci
Y+dfdDkLU3YSVQrTls2veBp56zoiccMiy6d1QiSTEzQ/ts4BzUgz1TwPjCyLZj9taSIYwYEI7/iE
wkFOqE0Qwfyu0xnUareNjKgkvFSLYWXBMzJuHYKZsg/Ah7g6bB1Pmxcgk8XjAQR1Y5cfJJVZuhSu
riVRAm1Mer9U+c8K1CuHCUzlHgO9StcdKRN4mp/C+TNXJfINeZOi770NVyTYYKTyddXtAm9iWLp/
XT61JBvnqfUlTOJXEStKmiD8NKPMzXvY1jBpjuMLJ7M/gGXow/Pn7iBKQ/d8ZGnjXLr3JY9D4C/C
9cRlqVjbUHnuVY6e3lwg/4K+bihpBADPIiyfX2N+VTYPAZM7MpBSHB9tMAQSaIh8e0fjWAj11WwK
fBqswZvKJRmxmcv5nDmODmOC6ViYC/ZioXm8N4nOF3p52RKXxriknT4x2OkyxnWUBeXAJwBEXc2u
y53HTAm+Qe8zmQGI1QUgSn446h/6Lg5pQhu1xlSDbhbpUASpYSjFzx/w2ewCacTlPHsFMx+JfgFc
vfRQHpTNtffHFFTyZbyts3mZItJT/6L31b9a0QWMlE5FCLcvpb6FLA903sYAYN8wHwrn0PjvAEsu
kyf4IQKS4Guc5JQONZRSlqcxCs+b+WuNKs5niI0K1UXaAR5E3L+qxI7JbUVpe8ntm8I6tbFVhy5a
yXywYXjVCYvCoGuPtD+lh0w/HtPfBeMGaSlO0XiF2BUWeM13hgCH2F1zmjgMNGpaWXUZ38Wag1zQ
BNi5kedcgCng5lxqwWtivcCXi7p+WzXBdyVBUMzenhdbskwP98aXN/RwLU9fpREHHK4ZQnrw+Sav
MjlJ329bQlMVCbzNI4VGHHFsMlxDGw1KxrLINfg4NSW4WGJSddSxDa4ak7g87jqNiCgbKyjw/FHI
ObUADT1If8M5hHBdEh6QXq7BDNAvdb2nYIUxl2xF386xVx0qQuH1QqWujuvsgbn/4sX5mL+BWyWF
jPYWxN/BJO3E3tOyaojBEaClU3XJXc7fMn+dWMz/TuN4+LMMv9r9Hk5uVGlMM+QbUkgrfcOHsGNw
/i8iUMZuezGwGqfFejhbUZadnYcdDBeuGqc1PuhjsrKZMnlznyz46d9iEb3u/QmHKuu4U7WpvDZN
kEUHbC0DTRerG+2IEMUDr/tBotAzZVTkvuIYwk7h/DYjpVpp+18Ocqyul6p1SDJUVVDrJP04jlOv
qHiwGk+IFJfCURvesY98GFt1Au1ThAj/bO+2QdhZL3dT4RUMPSvVS3ZbBRhyQVTsk8kgjm0OLpac
RQnBF6BIAnZupJNEjgiqcWljKgrTXh5ESyK83arKZ2iXKdA3Fkhr/DL7PUdXE6Z8fAivl0iUqc+J
O1mIbNZ30cW/O1y/c8txH9OWWex+iPR+apc8ZkTsQ/Q2FPuBW1/XhoTBY1fkgOSrs2VCQu96G43Z
taN+3DfcIVyLaVeEHiOdKCwf2gWwY/Tewt+ZRjYdm6XsNy9Hm6GDChnKATQHCeBBvqiBb6M+Xgqn
1+owbuaXFSNVVbISnOn6Uo1ZVrBEBoOiY86S9VcT2V3OF9QUcx1QrWQMPcHPQMDQ61nYN3MSbkzF
v+ppRWElBY0HdrqvJqwTH2kahfN/sT4yLqf7fNVlwMOmoLNUov+IKRUsMsG7ubbCJyhLofCho+Jd
yK3jWF/9Tlci4hk7nJblJ8t0BhugoPCWWeh5UI24KEXRGY0MLrObKf44fgBBUb6FX5hCsSI43pDa
eCX3HavWQrJupOH68/w0CuDjLrxVRUZ8i1CqI9fotfAzbnUiRFSR0oJ0T8dfIMSSioEX7Vo0tpHF
svIZU9dcK6pvlIm4tZwPae5WzQPgvuQattTSqrnZ0YKwgc2vqJRGI69pbvQWkPhWyINUZc3TArK5
m3rKbuemO/myndAmHs0oQ3FzR3pipIxtqxavl4GwCODLVch8jGlUHLzlViNrtiXBwNB5pAaUIaaY
y8eiiGU5t11Truy2nVXYC6v3+Gl24QqZKGxqXI4P2sXYfzu0PAUSdA+NfUAkYbSz+/CBqvodrO3i
4DceKKJyslNx8yxN6lCrxLyNrFkV2GMpUkmCxqTO4L3eM3v10r1vd59kKKuCAF3VUSozvLDeqIcu
CtFC8epMDKV4bInwvMcTKaEt3QcdIWmXslC5QKjhUMuoWFnh1NCgwqMwKDBt7Qrj3JCMARKUsmcv
b6cwjAYAXvwt2C78+sadSj3Hq4VTTn97RSOn23AI3zRK6fJpgILW2NOY9c9fMp7+eaEHieciYzZj
NK48TQh2+2RS5WsnYKghsAyXODKyD4kSujQKnoTbTrHxmURVDHAeckvPn6feaiVrfAoaDg8DaPpE
TnQxg4qstXhAAh4p+tMYm4IdY4ctx5ArIMsHZ5FQ9HUvcJlzQtLmFE4b6ANTvM9372I55Zg7oL9x
x4JnF2GtBpzzbDELNQ1ZPrbgdjPtO52M6xhvMGFAgn6HxKZd204eo2uV1/237IDVAlAf4lRZk0Vn
Dr86VUq8pb2OjEkK6QoOGxLwWPtO69y+OuN0cPH2MvAhnqHP/Xwb+BZ4PTbd1bIFxLVCkKGNtANE
FLQCVuJF/Bd2VYG8ofI33JeIijlItGObXc61BKZeebH4S2e3Y+DzMqSBbAeRXjvKjw7qybCg08Dt
M19DqnF60S8m6P2aJn0WODkm99vggCV+whuiQ3XHXSjxpvg9DSAPEg6tbADSOJwHX14B35X7fDNC
gHMndU9U9VQrxjy1jNqbjqyTxYSaoikI5hQshH7arVRokkvYiSdfgoBoX1exO77GLDs0A1x6xh0d
/89HaVgVHSK6NBp2+5qhXLn0QQ8Xbt2o7vQV4i9c4+407VXY0sZTVVNe+EvuZZtXH1nG8hIOFmbX
9t+GNukiwtriEgd9C1TislmLhvqXDL2BAc50sgmObg3cGbwWWncwUbNXyzIOs/qzTDEhajUJHfhN
qdWiiJvne9DsqkpXfFRnXMDnRq9g7SK0nyCoUPN1pP5YTdKOfFtR5WVztjvbUMLZzQv0NzkEPqRk
zlUA8HpdcC9woNbP/dHv/mv7RPWNwfctaYBsHC+pItbV+SVq6KmCre7s3U61puBXnxnMLIp+7iAg
FmeKd7kPtggP0QI+la/4GR2FAC7iWR2wquwtyIIy5TZT/ea9Qq0JYG6ni8A31pgpZTXoD0AoJrhg
Hq24HWq2YlAzWXrUQ/sokYk3ZfLD+DMOg4DqIfqj4IFu5IKelXxxCoaLsAz76JXKWxAooMiQ320t
rsjM8sC6TUUgNgdYRfNxw9IcseihCPU3l+I29Wr47xYfTpxcv0Sq6fQQajrQ0YGPFXF748uahk67
pUzQQCLvnLD5Acw138i8dO1LZNb5esPDgeGYUCJbbAgyi2n2NebhudKXxW0hIDqwwYsHBBufgfYi
eqzhxJm7iyh8okez3ZaJqiMiFQs4kMpMYBlQJZ6e459o86iYi1CIrKxpoioRiBUsiJG62HvbjzEu
rtjoh2a/t9q5l7/ZVQL+RVhqUoVH0RVhbDeXyhQ5A1125wLF5Awwqe5FiqBM40DRMAmhaz6u6ino
7+fWTvhufNS497wdHutDs96kM4V6TG779+tCTLovABLp8Z8fN3QMh8fYENzesc9We68el+gtWkCM
kGOTpRFNhhsp0DfHugrk2PzNJwrbO1/ZwKHsfwlg/jIXTUfLfQFeqV3roA2fXuE6x3HeOQzimHOn
oLTS554gmITcevX4ddGpVDIvzxtUATfYyDUb3ahDyEuzr8mKSXdz096munSb7IxyAYTJqkBeTk0L
0m4ni4iPpaZkSxFZ3uE7MPJmeifq+AVFW2/+9wE5LzSdtZhxIj8r0pdrmej2AiaipXyVzZM7tWIN
3bk1NNacSBSyjGfmpzId9ML6GRFOKSdFHt8MQQgoH7Y0befh8TxHrWMxVHT1pQ1s3eIGX4I4OJNi
dylTS4OY8zKaOdBMStekM92zYgFrxyol9Kr0TJq/ddBcE4zb4ZIWKs6XOkAq+aXn5P8kyWKSymvV
w3L89r2PWWwp0FsM+nGR7WQq7D2bRAqd2Gjw6uxKeiK3WI/xMxtGr2knyQHBsDfOmP51MQL3mpsX
qFyzh9fMpa4itRdCrSl/WUM8YIX1kSIm25G5E8rOJoOqo1KsyYVgQKDF29ycctlLKmTYoe3xfyG5
1WESGJe/755Ti6G3q6tLKv9lGju0OObdzTG0y9B0tK1YNHhIQJ6bv2DbxIiIRBqzi0jd1jvv1GAz
l2W2OEDfyefmKhqpkqB7SqOecl9aIIPv+WzDOefMJeGqH3zCXuVEW2i9XZ8Pz3PZ22wytSb6s+Ya
efHt4yhj/rrupFD0kdaHP96eVVS6IzaO54fRReCdOlC3DJ7J0wqqGmQ4/JBFP32Qxl9ykyaVVHE9
zFKCixoSU/x+dtXMd8owERJcRSLdnSfpB6ebwcG7T1+eETgqbaQM1UBtqV+KqAME89tF7Pja8B0g
7u0jpuvkNNx+HATbpCHVDW32J+rkWjg2DoBdxcrFCiuS5xD/a3DgVD/ddLztvNtT3Sasll29AwEJ
z3lhh5DJYDX5IVB3SoWQv8HtYtSV026Zz1SSu9mDWzmCc7PK0LS0p3u7t9SoHFZ6XEcLKObt40W0
ufr8ZEh5IA8KrlCmpdeRKyVCadwq8G7w1erJlS77ccf0RbqdxPTkzkZuJ1F2zbWb3FavdV9Iy9H2
4RAGCgXBq4KD6XOb9qZ01F9loXSVfmImmzXorxEt5c9N/zkDyA7REOBxf9wkFV5Zvl93oqZ2I2z+
OpicULpexG+09jN+foeuyHunf42fCIqc6oKjbyLadJBZc/yDNeA94I3dPBzx7jdfU4uX1pNt4Uwo
CTXtp/fULrZwQ2YQB2Jlz1zuL8qugxskB47DITCvyhtVf5dBvG4/y0PWS5AkPZcu424rVqJJNHTE
BAjR5MtoLuA7xzOKJXzhN7bd38ox3dDlJLgJsW9Ccbal2wI7Jt8ADusvjKl0cAD6KpZFpjzVOp+F
s4ErkBOOz922Nq568E+tUV6Lbv7kA6enY2r7voO+nSuvYK41kMBK8+gSLDkRgo/XhicQOhCnKGWj
ERzMwvjaHLVF5eZwo6C3E3Te1tV5cttbPGOeeoQoUnXkhWNrmNIJWm7p+fEQvdjeKfWVcn5PRq2/
M3WFM8VHrbNW2m4d6hVYCxc7WjBdQC3Kd3woH4ZJBoTDtzNv4FGSJjgEw+OS/lBr928Z3N5oWopr
MAfnnYEmcpWJMymScLK6AiA0wucc2GTUrGxcy+Z6lI/QNly4L701fobHIa9EcCqVgOCGgsfE9KOx
8zQ8UZ9sO/kmMQbCspDQhpYsqwvXllGkiiWgmADMpI90zfMPiAnvs4D1w1owSnCGcQcYqwi8nNIs
jhFA9Tq9PZApM0nyLpQl1nDMagF6DMAAiB2aZxsZRzBQPrGrWlPmNs5/fPmZuYRvcsNvaPtlCYjP
9NwBhM+0AXekruqFWf+7yA1GGca7xWBUXQNvSM9LbN1q9xNO4om7mEUf00NQTuZWto49ahQ9qacO
UpXz5bq+Ut7dly6bfituZwKvVjevzfcqY8U2xOc3qlEvAyzlil0DBHAJJkjNDQL+qtNpMXtryqkH
jk6T8zZbRJDaSWlvuOpJ+kKl8gUdfkBKV1OCoPKlRbRKBrfeVt7K+DzOUm7FIVCJbt9Fbh1Em4Wv
y39Jq6yTXRxbpo+SmqreYy+SKD7++GAWTb0E64KX0GulZKDtf0plpi6mcafO/MZjzHr4GxrYcLDF
bz9deFN10cyY4RnIfGhshdVwsAWqo4w2VlIWBNcwDuNd3mYhOnxfShVEOoK9xUzZDFIdZWz4v6T1
NhMW8CRw/KmWtooJ0eEZc+JBP4rYvzmu70H/dDMPaqekmENETmG58FfwCCXmCWUWEIn1+CNrJF4w
9A9X7XGOwcc8s7oiWPfrUT6e/vYxnZc2MbEQL3ZPylRkn87mYppLoyE/J6bBzxXXIpjkTHYQXjOg
YyTDfwprTi7yQwERWK8Vl52qdvClgb69XAakK2HHNWOECENG4KJDUetWTT2xbIwEH4GL/vRYejfA
XO38lRXcGZacY32O2/y/ceCgHbxR8fZrMi5QQh8O4a+glLhS8TTQAGDHc9MZT3C0nOKyBXWHjLN0
3xfeQ+VDNRwUBRbonSJt8J3VjVDCCCHZBNBmdNSvRIopJg6edzwCOlstTjZ4jlccWD9sk2CJk3oX
tGQ3G5rWxY6fgsmbdHvdkm5KR7goxAARZGWCtrHxaGaPipwWSyRVaJIbXEg24i1RVNsUzDErh0ZU
27Mmk+H6ogm9NpSOQYKRZb7+gIaCEaS9v6Gxh0m0ue1y7pqZWpSDMGOiOBHOXNP41rn1fwRjP+Ss
5kPiYDixXqwbraPaIVXDK8tJFnzR+eYtUW4Abibsqim48SCDPqprKzb0d0JRxWWFmpRUYhvfMWBY
9UxetH8xGVOZf1dp5Y/s9ru8Ull+0ooJ8syLK52R0xUa3g5BtfZtcbRTWzrLu81XRN6JWGhMGP5u
IJLz+pUZ2mvoeVhCR9zQnhVaUyAq70m8aoUfg2cV+OpQrOT95KAPR+aOOtOoL/jOjHPI1W++nNY1
mP5hgCDx4HCVVtYUU7rD8OSzOsdRj0jOpVyZoC+oBOmRJNaOkpUIIg8I3LsD+2v6QOjAjrR1DCrE
nJoHXTNoZLqyGyJZcIKc4xgkVHBobb0ugSZdHqwWjIe2eMc7J/JauHnJdFB3mEMSRnBwnEh9x1mh
MjPceQ1UFauhTGApraRrieBvY1O+gu5cTFMfFaIW3/pGouowIwKZdavTchjySNyYQ2UmomXg0y9M
KQicIMzcwcqZ7KxIw1I0iHI0G95n1EGyaTefLlk3iGUDLsZgeFFLj4M4kekJ99IdMSc7RT/wYhI1
PMj2bI1UbcT3KkW8NOAdEEAdv4IAIoOIP/CH7jssqUg7vL2ySmVcVLWuxxPzoXNNDeURfsG0l9JX
uXfsX+9AhlfeON6qccXxeTL3ThjuYfl8TqoZC8Q5S5O6S8FZxg57/iGJy4852sgFxhvREeIVRKwV
Ll7jzUFoNGeouWaxVRRkwDyb2PMK3wmvXRYMlZ7BGze2I4Eh+rtmqfoH+NoJ5FDrFLHWWiDwOE+y
XzFcRxk84fLq5Z9644CEMDBNgBGYO/NtswNcugb0M6H9flUYH0nqszf0+41qANifOII/RG3vHCIw
p4vyAsqK+GJit++jo+WIQWvry11ajsrz1jLPt+0TMc4K5YNs5pfT10A+YoGoJ1ixUr8oEm8hsTLt
MAGY671RKcNJCitUeRdlkVg4495YZpOK6Zkbv+wiOjThqriTuGqWKtJEnfie5bxSr+XfusJn467S
boecUyL5qQ+YSJBiMfGfISYo58ZqWWhBHh3UIrZJF9LkTR1g53enTMzKEvUlCI1YYxpyynzB/tHe
x9Mgr2XOjNXeBKaIf5dgbQsED8djjJ85tRqoKUco8DXt1lNApUDRNHaEBJkZsKDsD/5hFatdW0Xc
fqYakyF3Fj/jNCDvuwHrWmjZ3rhCDGP4PJagfi4cZvJYeV1RTH+PTcjF+N3hLnOSHroBQMv3hSz1
/IUqp9BjZuKzZdfUKegRGlI8sdFa+vJU3XxFy92c9zO4XMVoorc4rb77rN2GbljfECqOCPP4iHuq
YYI/HIWtjPmnxFfM6+0A69MGmjpNT+VUlgF7FXu5LzmRx7hjhZ85wFO0pUNQGLGyQ56WpFD+rU4t
2+s/vBX93WpxKBGflqODjzwPX1HS8CRDE614sZ5jUaPt9Jr+AuZNV8FHjgc76dYl13bu5Xo3YR78
6gERPY1EtwzRd72bEeDoPiNJDdzmf82sRmS9q9DxdrarXcOYmuKkCoidyLVO2Kr1iAV5bhqs9l+z
fxr+zIrDiGzeRciaxH6D16mPFJK5wakX+/5j1zSaQBqv845dSpxnff4q7AssQFf5TdkTOLaE7zFc
WrFbqPdzRqnbRV4A+A2/lzRq/uLLP0Z32A31N5qUntxlmsK2JewzIhcMzuXK4rQQcR8XaFyaGe6a
z469ckz2jtpDJOvxYAy3XufZFa2RNI5pI2CN/H1ALHmaqdjYDPnqrFYYjyp0LZ78HHWjxF11rhbf
asRDBwH3ouiS/AAJoStiqpaYEED+h5QdYs5An9e2VMXrTNo46N+Ko7fk03mGvIKzxvxRaPMa30Xe
1290rKT/xDbrVcBD2IhbvyKON6vhhOmrUUJO9zAMNp7qQ8k5MT5SpRHAnlL6wSJHsj4qkm6gJYSg
T0cj1+dBrt62LFsKj7Qq/OVu6q63H7YzMFCz8MEUjQZ6G5yn6hQ8dpvTYE0Qu5ok0tfBzRh+6mE2
ueSHrYCBHM2/0Pcay8IDoK1REh3YnucTOtu5uh7VxxwI4tgZXBTej6hxCyh4OMEKgD98UEvJo140
Axpsvqu4s8fbXfUVa38JFYwHds/lTWfXufxYaiSoFxU9qFwHCzbCrUbC6vcZ+wwhyl1++ht0ChEw
M4BZbmnjdUNczY7h1GPL/m9oqrgNHlQ2RXEk2wXCfwuhT8YH5Y7xiXL9Wwy+TCoogq88ATy6j/PF
yXkh759PUw4RM14bio6YDgcsEsrmQiFsKS2g+PBke04YhPM2rRsKrErd/gmaQk9MuF0mjEUZBD5K
cqR3yXPjGISqmKtNs+mVtr7wnRJdtH1A1c00qwhDxClNYSSIQwLeoXMWt4e8+8GeTKVG6uJEH6gd
nBlneFsFqGtXIAmxi5aSBTvdpMhPwrkm23Bm53tsU6tA6fpeH5Jx45rKOwaWhBlyCj/PyTJzhd6h
x8SDMCfS3oOSgJ2g/yVa1vN1+YMF+DMIcSJV6H0Y3GG49XwEX1EBOW+3rKtyvxomHy/3wwTv8dHJ
s0hIvN9nLeHmzEOMO/W3klyIxt7f3EnO0F09bhkzvDEWkN4+ConVKlPruXI0JzWZB5b7eB45Ew5K
QyxSiA5OqA89aA59hEG+xl+sBzI6LUwxgjWwAyR0b4DH0rNt/LZztbxb51sRsI0JTIfOWwS89MJZ
DJHha3aZ6dVkc+ItB78JpAJJ8Clpd3gR13g44lUtuAqNW+vQwAu2BVL6fAhAjUZOTwWPcjVKfaiM
A/6QPCW0/pVMVSooTPXVRmmhY6Lug3X1JvNEU0/vAt2onUZitPfz+UJYkl2nO64XRywu6BK2G4vm
vqJk2A8gV7pnKdMo021zHMigRAW5heFIwfxod1q6UuSsoeUKVFLg7TwARu2eteASiB7jBsi+3LD+
aWJRJg6w9gb/ahJCiTC98ajyGcMFTBvju2YDAKErrVUDjBF4lSoujxC/MeJfDz1CbEyQQ/vGPbla
8L23sRjiej9eI4AK3g+nVN54IrHR3OOdHRtOa++n1HQ2ltk66OXQqq3O4Lq0vB9cZD5yFRPMgwn/
ua+djbvor/AP8TGAp1+4nc4rGhQLFFP+Cm1YhI0PXzpGCX+qgtPTVUnL+UBZAMyG3OBJEGfP9VYl
fokBcS3SX5nsoBXSATsx8tsmrZyvCoypU7DGVWED544Q+XOjjSPvM7XfblnblNc1jjHh8wAxu9Zu
GHH+Y7McnRj3DrvRdjMZUhDo0nu0qRBe2ZgOel4BYY5aJlfstNVCQaRb9eSPVnqv6d99nqbj8rq7
JNTaYtmTCp+hQMoktgy69q7b1Jj7pOrGGbzKw+BpGKBB5oSKc11kql+P9PFeOXuE5VOa9kyjZb1t
jgvS4xup5A/eZycpX/jpobLUM/KEtm/lTqASh+n5Et5+MeIoN8Ch6x4gqSTb57v5RJcP2RzVnZil
b8iaDf0Dsyj4ebaf9xP2tmcyRsZ6y2AtGjws+NUhMa0SFtuDYAdRIWcW7KIYEnhkg1xHJnex3H2E
N5l43aI7GgRbOAw+u7v13+KJCVvUpyaTLJ4xN8sbnhUpkd70iA9qg+rnELdIw92391wJq+A6aAzZ
oll+8gQVpRqvPh1e3sLjjV7TM/iWrBXoMZ5p761Z3sMIqRxzULslK5B1VmM0WZOpLV6pT3SCotw4
4op2iON774BCLaXFrY0z7tI+8egGf2xu+2myW07jVu6jDAx7OskG0TOwmqe5ocRAO2m2qDFhk3Yh
+O9ozEi1k0+yd/pxgoSOpg95x9YOfaQLByBawCOhgcp/+bPl4loSLQYOftKM0bSFe9NfVNvntm1D
s7eptITx2N4DgIyp+IJHLm394QofMIkV4Z3AZDxus2bBLRyQx1VAp6Lvqk3/LEduDbtkvaRlRQKf
5rRVQl1y8SFw8wRF6gB53OLPtQRPiOsDAHVD/XhCvvInhaKXtgWApNp2SjizOTFHQ72XNG9uwO81
gmwzVJk51/TNd0bx55x7WtdzB6p48V0kNJhUCCux8wXloHeP6BFGPPskNQ17uqgyO7HlOgvWlfqh
H0IfKn76+L/h7xtoTC6s+1C5Km2gte0pJUIY19UgoBv57XSCUoR6KeC+bR5b3BGnTCSx5L/CVh54
Yrem0d7RbWqrWn+RX+dl9M847ZbgwWcyyiWmQhKGyN6xff4Uul9EhQ7BMzw0FQteVA3/NTBwOxCK
OahqZc3xyZL1aCCXXkCtQELvQjmmhQA2z/HZ6sZctw24elrVXiK7AVKm85aN1xIUnQR5+FPw9Nuq
UQyzaGIwFt5+sddyTGjROSXOJIZXEJU00utJruCzMNQJH/fmooQKo1lImxie20YYLRcEyfOudThg
mYWIXn7ZZENmVcIxKKb9QyqjFnKRM8YUV6FqX2FQP8VJW8vp4qtdTbitY9bYw2tPoscDzgRn60+C
AVU9Z5ZpD1+IXfceEQd6RU+B7jZmLjsehAy0oA/o6e8+MuF+CcrH1umYlpBKy06ogsnhxEF/VILZ
//yhaV/y4fnK070P+ryDQiTvUcAsUp7lw2asNmG5SbXVrezWKygoRepINoYnWSKVdnr0IdE1K3da
xuK5qiYUMHBrApZPh7a5EybNtqKrg4zFW6KtwF+A+P4Q1KkRTlP2urtmOvkJTe6EGgT2a2dt0iHa
DeC6Hukpe1zgMSvlJcHNyQH+CaI3pW2taYNPusIYV5fD2FPo9ozghu3vL5/q+pYzr9ZTXEDfO8yq
9DgAx0nDEP2Cmc/WAQ4FzM492Cg0YpKyi34vlSqwAuq9f/g0Ckn8cCRX2ExJUfItRc7JAUjZzh8P
xE8q2NmGltQyCkvaSAJTH2DtOu8GVq6xLGl75/KywYWkxV+LxqAKcIqhkIi/figxMTvJPA5otgb7
GZFJtzyYyJeL+YkOb0MWF/Gm789uBDlW6SYLNkE2F8QVOrFRfAki8gMSxkS4cKe7Uf55d3gKmmbc
fMZ06hJ8fz3rctXEVXcG8MqggwR8biYEdV1xqCPPBDnZ9SeWSzPjKFpK3kdsGqJTYv2zjULZorea
NQoGMCJtteiaYmwAVVlwmHty2hrJ5gDRGVN/bJj92BziDtZFDeLnbfqtzakr8JmVYBj2YmVctdfF
D+MQFjdxF/5ftAvI/4Ic8OkJrCqzdnyCodyuJfoWHqsoqhx/x1uy+yFtNNnOssoh21rGNTzOxOE9
woaRA0B9pL4K/0bLkH2Ro37lXgJIy4PJuwhtSJZz9UMDtGnivmKJtFPpZvv/Z4/fa5YKcz2m/Uvs
hfoVv5XKB8DWvMOpPrLN41N4QlGes8VWjDRPiYXtboy8alvOUaKAHPtYL+aSoI3+5OvD9mMz7GHk
Ttl6Evbo51QRB/t9jB+lNmOEPAJZKLrM8gHl/rZGYYxCfTBmVub0PV5xZq9nweB+k1qgLNNnlDke
kfNHW/sHNMFEevV+SMfJAbCzskKoBrm/pkPqSvLTG+H5/eox4yuNwQKOPJz67mq2II6XO7wzBUdL
rHYND/8F9Y1mjx74ikFyEr2vDZCBIRYOy15laCY91+lHN/PHv4defawPeR+yzxscG6tyRKzTi/+J
kTa5DO+zlAdOHcV0aT0IaR7CuPKAsbRU63NKDN9ObsyUKokX6xKOA8DL4RilFpnfKlghscPXgmk+
zpUvMxx8EuV2NzIVdKyfudcoxXVcDAOqLM/a9FtfOcxw1NejJeMUu2kQww8/hbV2HqajEPMBEFtm
3TyW5WMTXeMbHclieRVEXzmyKqsDZ7vgczVV2/JCUFSsMtQQABaIx4pLUKnmUGzgO0owX1CV7yQm
TocGA2gw8L+GQTppTRjFW/yJbZKLOiOqVGQe7G1pJwFMVSs7x/h2M3KGG/3b5p2nqSJeeH4tEZv3
cKkPkEwV65y4vW+dbd+PKj92dF3M3+gGhYLl8Vswtd4Dx3XqjANtv0jn2y13jIbIjCticbSPvNaQ
z6vY8QPP/I4vembtwanIHE9pCYGyMijSg+pJBA8HDXd6Q334UnLt157zIrNAflnzpf09cc8tVC9I
bimG75DfSO0Rkjo5RM4IKYvUuCXBoEYDBEs3ZT7zoQxPS2hoFmC1ucIbZc6+qpRAMbKX0CvUTk3q
YDqoC6jXOcpZQ6wVA/fDRE/qRsMvlmKPEl8n/S08TsLZCSKk0pWxY7BJCR6rep76tqNGzvUi9Crf
FY3dekJHBYcLe60bjpO6zMzB5zqz7rNcDH5XySeb+gUlh3DOBhK9bwQOT4g1yPJiAevJx9TDVBoS
ky1uPBSfi8WYPTbhXM2pFNoIsWpcqipgIMZIYF2QdMTLAsa9WfTiMdtKSewfGXLdHWaVulST48Ze
0nW/zI3GHSyFbJ1KpmqkPNF2zP9ewkkzVNaYITe1ShvVGSydXfL7usvMMsQkh2KD5Z8K4gTFGHvd
etcjUeQ0WZEB9xcNvydR70BSbmxrYaok5gNyT3junZQCQm/hps2jXQZXYvtIyDErK13CfebJdqHt
FtEQuvLRkHjwqpf415S8ys5DAI0XN8tw0uUPFamNQuoFMH1Co8jWqLHitbtsZ2lNvVzTFJnRTq9a
hF1nhZtnEcdSwGiwFHY/R+2YsV5/0Z7Ypc6C/emhlcbZqmkts8ON2HAzGJ9f5PH4aqBNOx9kcKVc
sWbXp0x+0x+FYge9ulkoef57un5tEI/vx9qy/XjxpVFsyo/i5nbRdWs97QdKrQOvj+coWI6C+ZZl
lEzTLlDNZcct+Pjto7d8AJe6CgBfnQ3ffOdiQoeDlR9FQlSLR5HC/bFBIgobpLOVdFtOdydoBpsu
f05tIVzi83WwXMGUVCa7/BhGL1mdKe0Dyk+Y4fx6/L2ziDNg0FJf+U1CcmecjW8TZKFN4b23KLUY
p2hCjMb5SAJOWO12XJ1wnBYpKUBl/Y9L1RwXJuZ8vZz2Uxchj7Pqf+jybPjLSZUpk4m615gKHMh5
eWczshi+IYT7wzoZjDJlg7XoVV3/t/AnJcDsR32dTPuPl9GW0hGBjIDa1wyYSQZ/9QFzCMYjDXCH
vQfm1up2QUDOlfYMUYcsF9WNt+aht66jvblBhLfo40yG3TG/i0osIuHCdYyaP5woq0gZCv1y6SU9
VGXOvPld80ZVmjWU7nw5mDJx4aGm+djPr5GR4t7ESFeJ4zY2r5ttd7sAFCoA8DtVPZk9BkrwprPy
QOamF/kgbLuN/vWOn7rG9A4Ls8KPpg5aTeQ/59BLBmZM01BWl/NZiJoqW9A5u14I55rOw8SP2+mS
zR/lsR9l6pcQvFDV84MsahCcioxZ2PcUz4o3YUirsbBaqYhywWZtcDtvYsiYdlTGRsOGcmqKCu9r
5nmtg9V7Vf0F38yMaSaqyCr7YUs+PwsXn+jpLPaCptB4IxWGXJaITeOJAs1Pr9aMEoyuxKLQKfz9
KCe/4R2SQWL05Bo7whEEnbheJuwTA8Ra0v1ZV6HP0vXVg7UZVmOTRbUxnLMoutO7EBi6pDxDABmG
Dt2v0RBl6wgNcYMO9SAKuUYdbANsybDpar1Gzu8mRg+oa9ngNu2n1MxT6vx9tIUaWmhswe95OCec
P0rrles9sKIiWdRY+hKqNY6OY55EdtoFEbpVRaHZ0qeUXOEs6xlMqR76XigrjpA3FHwp3tegfcMh
RJ42awIP0sVbmAL3xVz8xBr/iuSSXD0tp1dcoXUpkx050JAzk9BeWniC3LJSV6zUePW9zLMXJmNP
Tk/cor0TorMr7ZHo0mFsMvWq0GSlfvWaURVUnXUxhOKt3ki80hrX8w7fu2koBn80wljTY3ncAS7N
rp9alH9uDG/VxyKLUWF5r6lqXUWqs8PxF/wxr0oRvMovTXwBJABdPx3vnOrrr9RYupsLKmnk8S4j
WzEFM1lzcefNEg/TVKku+eiP6xJi4ZNko9KYvAIs0/BUQ9tiPPAXuobJ8BK/OWxzJmYw9P8TUPLH
3yb+H5hq3hl6gTZsC0evUYLeskqdOrXpIm8q0VPSMZ+8JAH5LOJE9hfCtx+BzR4FH28k8WnfyabY
C1WfrVQH3/OacOrvyftC7Afy7W91P9XXXpzI/TLYKlTPKWno96YUO+kpiuIhNb8MMI5Gk3zPBjAT
SLFRIrZvDDU6UJYmv2EgIImWheW0zKZ2zowwNaiG5rX/UZmiUMt+O9KiMr+pF/rVOJ1YT66VhQ6I
Xt5Fpw+Axgdh3XJ9moNB13TQAR+/gLXuODPk3uYcOf8Uy5k8MX2fNXldB6ayyfh1hQ+sip9lbtOg
gJEKl9z7dV5EtthU7ZgHBl2/gAVa+I2cZ9j8/sSDwjOP49TEBCdCQthyvQPt/knaAVtAK9YgUN74
6xjTO3GtTt4qpvQdiCY77lvhFvJ9nvFutfZoBW1tTtyoyuBQK9IA0ed2XYAKb/+ndYpzXvgUToHY
iqjRdAvBLMiP16O+tzhoZRdEU1yhWHfEPFPg/HX3CWgbp9feKDCcjMuV0WfGbOVgsQoTitmcPeHK
nCnpdhTk/gbUNcQ+hvH4PBJU8rH5gCxoLa4GosCSY7Oum0748jpFEs0eiMF2fLcHTtydOsN/M4Np
0lj2ix4keqt6Hc7Q+IQcxgRl9ORJdOwMeJ98EWtEH9ldjUNk/yi/oTQj1BOTOdpt/17fy4qK05nz
En5QDXyDGU9pXXnbcT25GAugVWuYPOoK5OA0TO84XE0iD2XLkSa4jgikqCCVpGtgQmPwkTObmlFc
0lc12TmnjexfQQISb9NadqQLu/MaEG+M78cJhdZ53Zw6nt4I7CsA4XKfho//5+r6/kZRiD+pUfLt
w+NcR5Vzsnr7T2/HG3kRkM3WrXViocK6Q/DBiBdd3bEGwq/PHgvscu4UpAPyLxZto3ix/INRttaH
HE//jroEAq6h1L735bufZBWyh5nJaqgHil50KUdWMsEpDZCn1jcQxAisU7Ba6TIl7rvN/ePf5VRG
N0KH4YIkHwgqHgS1RUUPEZ2WwGM/Z5oKqNM2QOIfRayCis8/O0rWahNZvG/bquXFvrHeJgokEAAk
eYk7UYimu32UIcCSHWpG1RGElea2iwtvEZ10Vdmlrxapbary4ZCH0Vv9wo6CZZq4phYOZ1iePUUJ
1pvfn8heHKSOdexGEIXVIc8KNx/z0uezPWdHD0sJ5xXOyGG8UJxlNTkYDfOMTL8OGDGBCFxSJkxe
C2tLOGQuBbSNy4kSDc3o9N/HvRP+5MYPPj5mXfJQhT1z7FqmfmIdAeFFTKz4yuHLxAuTnz39TLpp
txiQenUB7fxEhvF6ydWP8TeuWgbe+nMV0eOse7SaRfUbTIm+kniAMoykZdAB0cSrWuxrQ121AiOn
fiLP1RiSderLD2jtj7Ly6i42t8PXF0xz6LBzWdzHIIwE/5bTlzPE7ksCuZN4Y/ZqRVPfJxuuCkun
LWRnHQ+0rt5jXdJJJLO3+AIfhqkUX8zZusMjr/Gns/BaKqrkwNJmzHeQDeFKSYrw9g3AdUgfn/Cb
Mu6k395ESJI+5mOmeBRVP27/8oI8l4oQYdUDQ7Djor8L1E6zhiWP8AnJzmlM/QgnCFREBQWKC6uD
5ZdtC+42dYQMCUHwFhQxTBDY7A9CAcakrOebNsiaANHqp8h7eWloAFSs2xZXFucsfFCcpzHbUPj9
QO+uTm6G269g+5Wxumx2u7FC/ZSvX7wRM/458k/eup0btYiKfX/Pn8LpIHsbkp3PyhU1o2uK8xdC
DEGnsHKMnXyb4gC1pQ/rCfU5jNjscnBmjEFVjRzs2XVk6dKGBg7fGhJaLDh39abIa0GrS2f7muyO
tM1at537HzMnpjX0sRAHrlfx79UFO1EAnjMEMbYYA10Kt+TVLG4GR85BSZryZ32Oe1AaxipwNPqO
Ur6qakFUwOlEV5ez2zTazbB3uA9sJCr9ikHz46Fb7ib6nB71jL4CPEaUxDefVeTAdORzhNzszyK3
pyqViO8YPiKTr0ItBpFoA74vGe2vR+YH1c+X33+melP50Nlft6NF2GQJmt9XNXlXd1xWeVFKTgGZ
+YYLKS7F5ugJG8hQf9rb06kyYDU3UznqxhQO4ICCaamIaqqFiyEodmdMsn0KpjNPNj+oddWrt09H
YscHn1L1//gqJShqYbUVahfbBXoYvAuvtYqHUbdiTm9paljLBEM7AtpTe7w0mcyVyWEmbg38BGVB
+z4MMdFYBu9oLWnjEYQfHntuoyt9j5eX3CvtGitzjjY/Z2UbkxUbeJ7fIJMArGh5jVHqQed/TM+O
erPO+0ajeYLq+8+0nu/Kk0MalnDN3jLZhFCHChzAykdhcN/yDaKtqHLOh3rQXVN+uZY5G7CFvBUl
yF4CnbBx4Qw8Q3n+DEbwsQ8NAGqLbNStV8xP9pG4ammdC9MT/4Ts7xdtoopMBRPVDEv3NkpF1hIT
crgUBPFETzeYaQ0FKsqztjyL802n74IG6MzUVdOKqCnvKhvKFIXfEr3Dx+IVjnZwHHKtUz1vHB/2
saNnnA0NwSWfquKG1oHekEyL0shbbnedygIQpiwwMTN6OZo2aF2wR2ZJp8wu5yVScEQN/Qkocu8x
2jnpR1FLE3JloA0ww+LUbhHXpdAOCr5m4Gme1ZghqDmAbWaeE9zvspMC8FDErkzaHsYYKzA3Oi3V
xsHqxqkB5R3j5zE0o7Q8ddnIp5OFTZ6oy8nRSMGY5YH3pOju5no6vm0XDfJPM/WPDyU8jKtIMngf
vODjj0xFgcNZagqhfxu4u88O4XPObPXIBHfHbuNjx3Y1ezDhpCXZKUwuyep/J2Thcpn3HX8NOmtU
014PXH/dqdS2lqmMxXAJ0WpA5iUVxA4vNBt0AsCN7Kze5B5qLrx4tq0DputeTyDkyNFD7FxQH+Qs
SSjxP9jfbWuZ1PLSu82Zif2IZGKhDa9/LRDuV2Mek20PKo/pzx66FZ8VTUNWGnMOWFIObyt9UkFN
uo3BMuocJg82e7VfRSh6WReI37sFLqwF3BG/NFuKzK5Jr5cV3WpoNITIpRPZXLiiflaqeuoSj3Xr
S4DoKDW3PQMZhSHLVMpKfxGasq7GPbZOgj+AyBEgXE+3/FYKF9CGelv8VMQjLN/ljG3bIFpNXJnh
2Uw538MntxOYZUnozO9XrtFvoBuYh2tBQ4wD/ya83ZsAxOBkzAPBg95iqPqjL2cx02+Zy/vbt2cR
ZxnPpI6lRuukuwMHP91fkWbLn2ipuKn6sLLF9qnHoaScAjS2tHM8pnCLRduZ7xALR/ckZermJEbb
XA1htzwCQ0UnduZ5v3+jMu7rAt95lFgw7ZKMibDwaPtNtBar/aURhfXI8j4Le+jt2rxwQHZ9yOKx
/ecPbeaqXxcGOPwTZBoZ8uz6HH4wJJ41zeDU9yyfl2u9cek0QEfRqA8/hFSMZ+nXIhOUO40MrBre
aGsr2Ok2trcRbBcP1KRlFn3oPvf2uu0ZH349Vm9b0Fd+wI0/fsYXek0TvYJcCde7wRYsL8QoY6BJ
pQsN46xWD0BjBQMoJQonOrIIA2QgCk/43lKomtEQqkYkcq9hLcWXoF0mKXMGkXDOS4EZTuVP712F
FYZz1h2Y1sldy5eKocYRG0ecTcqDBGa4lOudAzZ5Q5dhkSZuERrfr/qDqHPMoLyuL4qVRxmH1Ubl
MAWWIndGZ+oxXvXqEWvUn3LaMJ8R45DdOgFv7pgDq3EhARSKzwmZT+Drgj1hAEui13ergvcyNAXI
ABHLdYwYdlfAc61IQcpjmtQuTZuO+NwwCb+MwAk928u2JNtJhYrQ6Zm+A/is9mPtAqdWIWgKVAfu
JJfAAd01ln74aaCmjAqW4ZzF3ygRu8FpUppbtxd4kF47nvet10KRvaY4aSCft27JHA76TwgTbLQt
8vI0LGwcz5fEXUDnCMjJ9N7E6EXF9e3poVnNxT1uEdu4vrwB1eErRaB1E8xsysE6rrSIEoc9Ud8e
g25Ud+ochXgxFNJAS4pxFpnmmzT7ab3RFzEV38jQt23rcYiJfBoxonZ0QVb1PB05DRAh6dXP4MFx
K9vu/QGpiDIPzNjDOuvX51DpdUms5lYo8CZEX3752bI353ITBEwnFDWEc2/TmZlNqakT4TGNJQJs
UWkIvKdQkcQjHfgGFEKD7BsQPtSvAsH+fTC9eM3CAQYDBhT+UMdHii7CQP00y9iBv593xsQr4+WL
Ce96cFDeOVCbyoxUXnV6c7dw2ciSyqMweAqHBJ3o6Zivec6R8Ir9jL1T/oWd+ZIeSa+jEx2+RVcq
VxKfjcLbdlfCt3pW5GfVP5042PSAVDqvaHc7mjpl8t6OvuihgN1F5Ovj2mlL7iD6bPxaPU0HopSV
k8PQdDu3i5l2YbWJZjxtBN1K0WEtCD5EWFN9rghCHwxAFkl9Dd6B3Eq9H2oAijdnMe510p/tQYUX
ms7i6vmNNEGfKNRyEOSOjz1TmckH+3Dt5mZU38fghQVZp4+Z30d66rupzfX0ot0/Mor3NLjfm0uI
MAXtWJ7/SDxlAQFCVxbpklxKRQ0os7nrKFlyX9GkhYkviqKkleQdELN4DQ3t6RbWWX7LLKiHDET3
XVkEmao1Q6LsBmA4ix9olpukJ89my8+ehpa+/9CuoR/liPvM5M9Ak0eynySRzOQSKgJZmnlkbgyt
/tixIoe5/FKrX6qzSxzDad/BKrl62dDKOeCuLTR7LkouvibJL4+I2hHAsaHVng1R4rAw1rr2oiVp
MQ9KNmOfbDpKPjxSmZhDlYLXYzXU7oZuVnzbx6CGcoKOiHa6UuY3g4Nt1/hiTOEOvllS1A56nV/H
LcBBc8AJxm3uciEndaW2dGVHFfXxxg32kbUrBKya0yd8bOPlT+8Iav1Wy8ZVQT5dA05vbtw/rcn0
NUufB6JOUpGvHwpLfb0fC0KTj9aoEHkptGyr0Mpni9FUHplCo11Z9wgr+auI2Rppd25e3RBNdsif
HM0SGHQEMhGsiy8BRYEHLu9wpXrQj2ykN1VkMamiYIgdneX3jBZH0dadjG+Dc8pol4qVf69mF/P0
crXdy0O9ds7v7jDXknPsPHcH8viWUI/wNqESLtnVeE1Ak19tlEdhzR3xM7M82QYH1igXwbiCWRu1
rRSolw0VF8xaoROW+1IEOdMN+S10tAvIkUSjSOkv0paj0WmTxymv8KQiX5TTDt8QozJTDvRMVAYI
2I8EfLhVF102WiWE0dwcxpuawYyM67+lys8dEeZKNCvmPFMwz4YY9EQK++vc0pUqAjzZ5JZKmEfs
+ruebvVzTZ8FZhOv0NiGRzSChuDeMlytxswIgpJABv5XkwDRTWqPCm20ghLpsf0uKqFY0rApWoTg
6JNbyUgoQijUa0wicPTYH/m2ZsdraJ9kjDuK10BTuvPJ876p3WlC4RvRXm6jqzNvLP7mWL5+1BE6
ItVxedOLp1kG5O5awG8W5SBt8plKDxikJ9ISx5NvpSWBa0VcCJZjgGIFZ4K/cxaSvJxoOzIU3OKj
6NPIkh8cFsOlYz5pvFhSsODjXof/70ey/wI8ynjXJG+t2K4M15siFji9LWxP+Ui23fREX38fsQ6/
HfHCBSmDlIuwC5FZSolKjP7l2o29qeZUv5S6H+LAOTQyKxSKkM6wUucWM6+bdMdUJQ9WNA1NbNPm
TMm6IUOm+8G6A0FOYSbs7KZohV6HtpXMnx5yVgqAYxo1iWG54/SPd6pKwHk1DINqpF8NLaf5MJ5Y
HBHLJj/GX8OuC+6qZozzW1Bnu3fX80m6TVkvmqDa1ulKWTVb8zD9mEwG3etXPrLnL6aqMQ2qpQWt
Fw01+SNSwMf8TokjAY3EIy1VXeUv8MjYURqf5Jrs+B+nnOyrss4/DulxAcySSnvSmeCKwC26MB1p
lckyW5uocfbG/GcvDzMvlz3ChFRHhphudZiPnVxuu/d1acCg8bB1eZ/lMewFNuM7BQD8kMbhuQP/
1AM8B5tbjQMQHLNmU4BtNvxRomp1ZUE43R2FB81Fy68iUw3BkvuGQ8715nSJB5OQVf6os95omsiB
/xqKtQmjD7hDi6om15NLqsM2n+z0Un67rmc5L7SH9aPiNgwlSNhg0to9E+9uCbrBpVMsrWunVavJ
8VJpwqKtBHLyQMSyjYZ3Nh/ZUlfBbHcfrkTSGz2lt0XPHhcv4I6QkuRx+T4mMCTKiuMuJvTW/vvM
PC7bBh7x8qpAeiApwPvqUdofhH29FqTem+cAuX7eP7IrGPqd455M7OOgKCKfMKlaZk4ao/c2KSjE
WTUavDhD8IpuRBVygoUEIOeUaO7/q5HSUIqnvOiCUD1P7d0nNGE3DeGGb1lRTLhJ7DqptrWwL8lt
RghByUB89X+7W0rWxWXECpqM9FPWv0IiBSwKRwOV1ybQjeBCqHGvS514HMHMtKfsCxcib0s3vxOI
XeaRE14ssR4NZLzXVHW856Zed2u9GAKKVvQV8mIHNbVAh8xllEZsHbzKNzYMQcF/7MXHb1MKZ/5/
H+4Xy9aRdZjIoqYa9WBUZx7RotEiyBOjLUgmbnmWbcO0nhVuq9z0xDrgItM0LgQ0b7awa42C/QSk
E4GpeTscXEBwdBFjYxbvHwwnnpnnUCQK3ksAv30Jc8R7Sx8yyJ9SKo9yWA/mQSIbBWW2SKsVNTgZ
L8UGZzK6a1Jp8KTnIg7eTy2uDMHST1xb1gB10P3BUISzVoFvPBZsYOm2wIxeJ/mnSxCWFwG9VFxz
sQGIQJlgKMH+FZG4txU9MoqjV5g+8OCPvV+nOBAo5JRyquTiKESsvcTe7WKGw3M+ya7SIFJZhlyd
Jdv1BxBnsgHCXmOT4egmcro+YYW3kpuLytFkfA4V6/mH/7WK9hCTxc/9GnfEkdIB+0joQE7Qocjr
32xMnf+UHpuGx56XzqMAik82eoUTYt9VTTVUXglkghUOADNnloA1QIfr9Y9gv5LJdypic8RUUrny
nh+lREFDHKO5Wva3IKseDJkfPiKm+YVfi/lo2zJi/mcTc/eeA06F8xvauC1XOXSqNv+++r1Hy5Bt
qD4eahKv3Uw1Ktf7AdCGWeb+kliAmSmyB5II4XH9u3pJ+7X63vGgzkKo1q/Ts4AAvPVbaH+Tt748
Id53m+tI8c6Cz1ARqvfZkEmQqW5GCiIBIwxCcTNfpiNG7ZmeH+cjrwfcLuY2sgxYieFxZyLwhNBZ
wwl0yzHiDKLcmjZTZoMdqhbzVLIkUZiiBy0E76X0bpylnyiKPcujBf0jzyj5V38ENBCnk4a/jDva
VJ17sn88t/lAeOM30zuIk/7mKiobcFIfNb+oU9IpK6jczjqLzacujree/iB0MG4a4j1E7s14Bm02
o2P6hJDIaZE70vx4bmtdsjCzeQmivtsxXiarC/daQm3AsxlexUXHGAGtQE/4ugX8Ts0pMECCWCIG
X5C6hZF6aLuyVMGb4RXZ+HaWcPMkDJppUI/Al7UEK7PbZShPJvzvjnGz4SswMmJP2mGFe7Zk6BQ1
5ZnBq/cPHgdo0DZKzLFSCRydcJ18vOsyzn9rnDzWaHewJuzvAlNLpJL287jqvSN6aoyg/1hg/uOA
PdBkaIDNHZV76VA14Ie/PzbsMU9kkVXxG2PzMJEqR5VFBufTT6x0g+Ch3oB/aw9vu5/oRhlAENY/
igph8/oEwO1zM8a44DJA6x+QakMpK4OFHaB1Rat2x0wBrMCYu3UMMHhPV5TTrx0+jW9Oj5xGiljj
mioCR8T5sKc7KwGbxAIshXs2Lf58MceD7uOSIFlwY48HdCoVGe56u1Hd4xtt+MycDHrjJx4DP8JJ
U09X9H4hQWV5cbIg8FEyBHcFJnuTOSnm+XWxcGgkEluehIiimxNr0wEEkkLmE0asF5u+LHjE6WYX
jHGXmXULaUBeE8OZ0omIitooM97Jw4aHbIUlRRenZgP6djjVLpaMc8vSfY/xtBgbv/9bcqDQSqUW
aZtLz4+F903jafd+Xl8OMpcq5O3mdJR2rGM8kZZliVImJPqMs1434xnKd9JFyFl5hCTWXnXwFciT
qbBI3iBCQuqxsz/jJ9oOMWe2QFJFYUM4EHRX1sSPUwZJB8EyfY2m9GARL0+r3iqdfCLmU/fJVdRU
WQsZ2xSCfgrU6QvOoaARH0c6LAgGhe2OQBD6nfg95jZsyqr3nlMmLGcXeoePS1aYGcKRnXN1/ul7
pegPkViUdg/FCX4+K/byNOLVwALfrK5jwB9C17kbHN9Hy+JxwYU6c4GdBI81Fd6BP4Qd30nOanbG
J097mVEsLrqPcRxP+VaVYm6pvyH/xZh3qSBMf5Jl5MsPSKRwoTI46A6Ljv9+TfYRUMMzMyuxssGO
IdUeT7hwZ6xcQ9Jfc+lQt9HK3HH2B6rUkBiBRmAS2g/Hv+x6N0e4UijWn4OqCq2jDtKBXuJg59Dw
Vo4KsF+ES6IpT0SgD7eK/bcBuko16QLUSl9iQgmmmlVHjFcrZkpCLDLgvAgapKuQN0JI3TJiZMD7
VI8zHLc17O31ChHNSPrQIHJMDKYs/35eCdNUqoNfagkNMyxJXJiLFZeDU/JPaKkGErtmJTMepvOM
glI2Rjr9P4EjuxHTMX8bYjiPaY5jHsILlPC98oykauKZp0JeES6g8eEoGg6OHfwWue2Tbuqk3njA
QF8S6vY5X17Lu0nPCgIDtcGnLZpMeEm1yQqlDkJk/6fN31i2uw2O+kB+TDbZ1u9ukwGpCBTOvcTt
c3H+b4tg8cBweJ2LRbbelbSJi2sl/ignLks98o5lqfiTGADo04j1eNsga4Vb2qSfKCvg+IMSUzJ8
KnJ56mnC/5BVdppQjHC5J/2yJ5gmDP9d7A7fPuy4S7euef1hvYI04CfU/uvLGzN5DQmuhZ6Ez7D2
Nuw7aupYU4MPSL39mLSqfflprxvuTTAsLZ9i26gmob0sKTIKhys4TjKl81AFbs9+MiNR4SbzhPId
MmNSdGQGgD5rHTsBe6WiItkLdSq1dcALtwpLa5hiB9KUh1dDJfS7KcYtAJTTQCG4UJRyVTTgZDxR
6i6cO2mzBzhdVuBSFKrRv+CE2b7cuNvr1tR4EbsfRElJXRCM2lXXe7DDuEFJ6+OZnvE+dZfaB4YG
QNjRVUVFLeec0bz79y98prjdkVCFaMga2vPblh4ZJ/IqSAZDrw3dyTugGwRc5uSw2kDuz4pktuoa
w0tIUd5Ia6EimffhROe8zIUpq2JH1nhD99QGEKrMvO/faABM1XJO5y5YAj/0F1jsVBslv0IDBx9S
nmOXskalTa762MDdHAd8wA3n+OonO2oKQ/zLV95zc8cugLkXhNjZNVLYtA43MVjUjNP5MgKYfVm1
M7IddHsvCTIoVYtNP5+ykI1QTHllpKrJ1j0eSOITQL3riWzTAKGjz3Yuxb+J+ikpRDcppkIhLmji
t8XxBPEzIP52LrvnPmTP+Q71YdBycgHdjNm2QulV4CENwfJNvn/BUamr4N0vHPZidqm9cXn4z9Ou
LKNEncTIGBuMyoqHhyQOSy8gqGeoc9dGZvu+TEFfhTWzfXHmy1R5VOBHEfddf/rdJFEbWJHJACfL
GyDN3WTrMEho/Tkm1wkpRG0etCUKI77LnPtjGT3FC2eLcAvDxOTUaV3qagJ6hDGn/P5mQQicHBRK
zx6iauI3oXqLLs4Lm7MEOCmedv8WXyXUn5FgmtrnAi8fUKuMKR6Qx6ZcwS9J4Y68u48+/P9I0jTC
duPg7wbzpwMsy6wb/UjPlohJ9XaaVf+NjxtzXWuaO76SPc6D8dxzW7PmBWRqpCZDmQvi7WVTal9J
XQAwXwDt7Euiz0FGqfOBR/WBX1JFTIwcYPxeESfNSV7Qehrom7HS29VhCAO6aNrUW1rWdjh/BBw8
Dcud3l5zk8Cdy3FOthA1BtMuBtHn3lTBAfD6eABwtg3fjIi9EBXt/02vGkZpNU4xlJh1w8AxYsRT
K7AAZofRbjwJWBk1xJB8+AF77AVY4eEIKIEsfd+jR4K7MaL2FdgKsGfA1qhrtIHb3cOPs4VlH846
XfGqv8tTIPwAfK95QkL08Az9k0NJ0G4evEp06cik9m0IEamf/SRm0OgxjrWW73/wWYQM2evubEif
AyUIdkuBNiKXrTvWkFJz+imn4vMz1fXZVC6WmD2wzi4Glft4SfXnmeApDHZNn6LlknXSaqsGuW2q
hjlp95yphSro9JEOldmTZ/GM5n+fxCrwh41ZiC1JlvXFt8TbHMA/7sJZS2XNgl14NMS3UEcpg8zA
3a7ixATAOwFRlL+BZra6F+NIwbAAeuBN/sn23u2Y7HUWkJJ7D6q2x5QHAkEkRQoGaPuy0AgzG9Jb
mokieJo4yzW7Jddd4x5yJhl1spb/LZDZc41UUNSthdv1RhrTK707w4XHSuQuvA/gAffXdi97Eyoy
Kl/bwTJcE3g4boTBRov36fwUSznBOh+uxu3bkilqz1NF8TsRJ7B55HuRtQCXSNBB06ZPttqLVC7x
i9OAkyXFgKAQESNci3V1Ef5WLzoeZEBZwcRiRuqMSinFf5pfO3e5V1eG9tiZPRwf/EMijncoEJao
oaBYLGMsIYYCGPZ9LXYarZA91s/He+bK44//cMI6Wsi3RXPAjkwge97vPT7usHLjK0FzqtkFvjDd
pYSoES5uWkvToF7fRuTvgBsMNl1RkMwCDTCCarbuETfUHa0kcs9qAZvb846T29WRYgKO3C/Rzn7j
Bh0pHPeOUdPMYeEW0oCjgq+0SfDpmtHbi88UUSwxrCOBRaMKaB7AUCy2hF1lT8zrCr4BfpTNRVEc
8H7RwTXccLhHtvFQMFdu/DEGY3WeZ7l0tddXAtH87zy4+wmaQ7Qhvt7Vrsu6odSASV82I0aK0xXO
NUG+vkKo4xxncGT8C+x3XOelsERFKEoRMSttsMK5LyvYu1AAm/4dx4h0kDsJ8RKo0Zz2d8hnahOU
ULicVI5o23TUv6UjyiWAbQk7kwwz9UrlemrvrCGQJZMtFOYROD6kgoHG20fcZmMAmQguUi3sKtgq
QLcd330u6bgLq3/EL5bil1ufihE8msR9nUq+tlqkcNKGes6zS17RAfSEqD7s+dfy4b8c9qOU6mHO
FGDtLLLC0AS/UM9oW5WBvUyPLQ+qMSqPCI7a+nVMGBHhs8ozS1V2C3wfv7f1voGZQ6NpaJwDcp/t
5pdzJ1qoV/BxXlgTuQzmO/Xw4pzL+zQpjTBJoWr6enYP+/xNOblOndeenw5cXZHKwSv/DFpQ7UDj
y8NCqkrMqreJsLJtjcUFasTWKUQWC3okSOUcGQKrYUiTev/zKGtmYeETEU0R3k41zwb36DacMiMO
3zirvZK3mzDqJMjyOB5WSryt+sdb3+rUoo1nmVyd9qC1XySH9D/tTktoJ4QZVi2Qrk19FhrYJw+H
kPr+OnCclQj0KZX6edqekF+xssnXwW8U0rYV069KlynlXaRv+igldlDOWO3MOtHODFv4auMM2M1+
fLmhDcicf1knkfClU0rHgbAiJOrLvpOdF6Ou2boeiXaAcfqSpnpwkri8vQGhAVgtL13h4RhktYRw
G5iDr7YXnpHlBD2P67FPYrOgKUvaaKfBDlSGzGAB1HAL29LlkQCRfNwRxuUKEOLinPwVa4v6b9jM
iUyZpJL5EGjORUjg44pX0YrJlX6M+U5jjh1Sk075FkIy0Y7zmeNpwa4iNcBcrgn2nGTnWcnMnJcl
XKEFA4I/2xIS0cu9zhBdpZvuCYsznOV6ZfnEoeijEKGRALvbDQGeykUU/WqMMtojpxw+k+62zsOk
CpVeo5yH+rR+BbUlgBE/2HBxs2JkWFQUmpMzR9CyvU79IqJh4TGJvFG6rcES0Ibnnh3BwKRs3DAu
S1Y2xJQioDYcO4j0UqrSbBhtYi+FQSo9do6TE9cJGYh48JrPT4GFXES9OUiv4g8OYKZqbcMtjbm2
vZyr+U1ga8eTN762bysWD+e/EbTGZ/BvUxBPCXDFjdRxtuDxczZFG61M7P3+wiRQh6QVgK4COQf9
4E1hL596v4XJb6fg8/h3X8Af1cKPQzu1ZzexwsSeWxKdpKrHqw4x5CiESK6dW8zxphKv4s0puII1
emBvq1XXCwLksdR6bVuy7tlXic8DwS5EQ/lB3DoLbClG66H2HHQQnANKpPjLPVlsJ9kc26vIxWfX
9fAhAJ2NLGxjXg+QsaGmTJFAzfuR4G9yExCdoJWPGg5iu/H4DxR+ZdgohOk9k6FIHYhvy9+BG6XZ
eSxPbPM77iWqnqRn9inAtwWG5Uw4RL4A33j9qi4nnDIwacdbCO0OYqEO70IiLKTymo9OH6EUJvEH
LMRW++rLuNkQPz6fs/kvsNuhKlWp4DEw+jHUTVM9909r+aizXrgP3gz3QGWg7hatKFLF6SvOAPM8
qHRJVUYc4Lcp8r/5HGUFGJVg84K4p0dXKRbzcXaiKe7Zdqjhjqndx3IBQQPAXNzFx9yHx3eTk22W
pXwX4nTZbNsKUEEXWufZuKlzKySr09a1kLA/G5SGVS/AFHIIde7BqaySkQNETGO/gINyBCCwzrZs
zpZIdcgKZlcwRmTH+Y5F9sNSkSONSyFRn+oKXg5sOFunrMRX7D3HULOXBAJn9/dijzHgGMX46S7R
kjP/Sp0xQbxgZhyRVCuTo75YQMsG2eoFiP4jNin2O9y8PyqU82u2E1LmoJc3lc8QY6BZUU0OFKBN
CyHJOKWQ7O159T4/Pt+ReiojznknFOS4sstfn5MRsy8eKc6WL4sdfyJsz507Pm+xxS7GyiAiJCYw
VdgRn20wL33lQmVDHAuzv9GiqTW3l6wc0ZAqPpR60rfLNNfBnv4eSxyN+xWeiT9eC2ZRwNBRmzHM
nCiCrF7pRGDl+84jJkN/Ny3L1d5CcKfTegKeNrs9/k/AZ3o+sFJosWnYWOvDjKrynEBP1fNfIeID
F/4d9GAl9ntVZhg9ldDNeQjIENjXhFHrj8KNKt2++V/zWBzFzLnKWrKBGlPeDjMiIQHC62rYakGy
5cxxzdOfl+Usk6bq3VY37VVat2vHjEm2N98o+muMIez6uxD4l64YZh5qx3aNM+V98yFZFzlv3e9x
Hl6TUVJV+X4K1Xc1XSFUlBBStfdwNoyAe6yzZ0uJa1xHFJrXVcZteGZO8oK/ZMzq2G3o3kCP08zb
fxegDvKboYd/gkFMt7dYpIttp23diShdwea1pUHBMhuHwW+M+UH/Q3VKoWTqMBNejwoy8g5tfTIh
FArqh2L9giqktPDtOcljbgHHV1THZvGRkaMo1Efz6ow3OAMid/YFgwbDhFeMYvbfrOIJ6U8376Ux
/NqXsvIZNsBd4Sf133a1FOkxfd4jlZe8D7fd3QwkwuZflrG+JGtBenCeNRNMTlTN2dFM4qwqE45U
V5IWFZjPP0v/xVx7sP6nHIITjIAn1Blz7NQKGlWeTf9Y+gpTkb0Yl6xcL94kWukeIqT3NkhJ8NRs
IiKPQO64Y2fjfjla1DgY7Ii48yxgRf9rswnBxgqFjH3TnkdYqwKupwWO4iyqhH25IqE6SzeJYLs0
nnb8n/xZOAloY1TU2gdfnkX453MLH/E7hLVP86BiKxISFH0qGOKiVySrDTI6gKQ2IyvKuik3SIXI
i4Uj9vnKMopX1NmgZPiUq/4QARpmR+vcEFhVGEgsi5HPr+ijn79b+hcVUwBwbJmfat2Fq7hzj6v3
9ZAPhrG3cGAl90b23MaWsGWG4wZTzMyiXvwcJNjIRsVgtpB1h3hirGeSuJiPJbGMx8RX3XYPSRDd
GfK2A7+vOhU+Xss2jFXlEeStTYMI0O1tyMsxJsaC31th1v6WFVgjJQlQpTm+cRQMIFNKFLc3Qm4v
hFnPBSZdWFMqQpdopfFVJHXQRPiUeyq5pH4XlbRTR1vzfD/t5TUjStsJPOxy0fSZrd8gu8f8yrA6
YqT9GPM//+qkU18WeGp4oARxID5/JkVFsom+7l5AfSp7Cm7He/GTtllUE2bH0xLZ5q4w33AHaHkh
W1erEl/NBsmrt266ErMPGmnc2iVYXHrL9Z0x9sBOQ7RV2xS/qakkf0+DDHM6YrOZWPvUtpuD53wv
4MET2CUgmZ9iuzHcrotdGm26fyBUGXURH4UHhAO2GbY4p9G53ibdnCowDI0WAHXMgWgRAr695FWC
6P/ADYWGZ3GKKcJ4X5pnySpj6T+JFlBH9Qm6VhRYIszd7zjZJkfcmyysl1RqN/DZzXEi7rb05x9H
4JrCX02IW5XUWSm5Qb6eyli29JrHO+/xjKiTAhoobihvH/PRu6OEJo5xIGqsJJBqhvLGOb/r8jw4
/8WfebVV78/MnApHllgsAjzyCzC2bbEKZI+6EEsRvWGSmKBsQ/8J/ioO4ZZdhvJNzQW2Ycrfe4YN
lnMk5qOI+BQqy9mM8rDFG5puOuD2Yi8XceGkfPMJ1mvmTOnIEtLnnH+gXpzwPAoI5ZHs7P1Mxlvu
ugeuEIGode7xdz6tFIIEAnhgVlq+YuA20aD/I3g42iE0SQCjnpO6ikWdA3D6O3Cq1QrXHvHwxMBm
JHXNCc1cvs/GtYBaRTknpZJZJ33PiuoNYCzt/8wHtGmPCL4fAndzE4hl5ZLdOD8aGug8HoJcx7Zq
QAZKcZNjVxqqO0y1sfNtnFQEfiFRaALwGXrmjgPKjxMGBqpezqOuZdKpMNAdqqOahTBACdLRcTR/
OVTzmzV+sJ2Qd8f5ND3m2eg/z4ksI6TzkTopcagPHusEd4OZwBzqO6qSHyP4qhvn6yMiNXD1eK38
ySHVBfuL9ioQwMMmDE44OBdlX+Qo4JU8ptqNHU3r+vy1PlJdyZWn+WhDJLArjTG+4qIDGKvkbRTR
pCLAjQHz+H85ywDXB3PmwyC2kfbAuiBvxXD1In6aion7bbzkmq+jf37Y5eBAdAGAUraGRsvHopIy
G2bBoA9P82qO639m2JpR03d+xmocZ4Z5bWgoZH5xruBmvdYMgo4xUqodvdYO50rbr3qdCu60sZgM
Kv5imn4EUJY/zBHrtAfmikn0JkVoHhlCsh2R+LNFfWBpNM7mxZdwbK5DFEVOqMLImVA89xo5wR+q
o/j8QSLq7pAceptUYZkWUTcFbWfafOS7Tk821V9SGmVJe9d9JHkm++CJwF9pdJpUcBgZGBrdFF/3
dxERRKjmNs9Bjju16pEb1cQi33Jll+7qasL8+/0tMCfKU//BTvWBFGM6JCpMbfo9Tvbis/wO/ESI
Ard9m/i21Ey+rTn5g3QGTsxA4J/gfdpLp45D+6KFoJBIz7rRCnvGrEi11aCc8eb2YTjPYyXA3wgZ
eFFgEg5SsS0YrNS2uQSUt5UrIEwbZe6jeFvJsqrswH/4aw00CguS14aXTZna0yi1US/cyKuDLHLP
r8/5/P1lSuOTW9iP7TtOdKv8z7wjIf04m8evQH8mxvJCjR0WiPf+1pcmFg+jtUonjVA5osvzTdMS
UNgV0Pf8A198S/fHUKeD9Mfjwxc6EFVDA383Dc19QnzNk6E1cZgl/UBjC5ZVYoMfHn80ZTDpHvbw
zw+PdpGnSfdr3n5o7lHsLj/3Gp4nATSyl9NP9dd1+jq3CCXIc0UhkbHQ0vWMc5GFplFwL6dhpmEK
zc/KtC35TytPDIoOmtThd1ZaEd0DylZqY1kStqNpJIOZKOUEG1HQ96JbafqiZLMq/xlnGZd6MnAo
M1gLHbFUeR+qJx9rN+UnkxK8Bq7c7Cj/KReXv2kQK+gXSEd86QnNIt/9KkkjfaMvT4qIzUdKNt8u
cpuYkL00MNwzV9OO4OVD7xSSp4KbFSDqP510FggHptr6kxaKURCSKUqG+1QGTB06Nz35datTw+wm
A6g6a/S7yk1NDAzoq8amJrxMlXWQTZa59Tr2gCPlzaLZTWFgSi153q6URdo3CLuQ2ipd+LDDaZZ2
iBI2dZgbiy9sCv6CG8a8tuuFpUSdVTnWT0rUu75BkBKdXgNSdqTc2qCBt0gkePSSpJdeNvDzaBnX
pj8TgdeeKNY6+zs+GHfCi8bhXgf4v0tqTFwzgJdu+st+5k+bFDNxGgEvfL1tkfqqHWfFbZEL2+gl
RJ6EeMpGcj02U0RGDp9CoPwAlO7T1MmqTYkCt6vwDswrKJVhdcjdy2BqPwawvGV46AawqaGcdVO2
gjwFEtlp5BpY4AdMDsJzmzul3B6Za+/CNnmTqLtb41xtFIxDk29PE8hyjzNx+XGhKJDl3XR3db4D
XXDapuEgI4f4U9sWqGmjKe6zbUvHN24dmMeE8yQXnMbqAf68alTxi3C3XS4s4pNdWjXWCWTxI+Xj
JWShL+Cfv48VWfa5mR3P/f7ePFSPCe2V3iAllKRd+aGHK9sXI9nDNebfWg+mVXkVw3RLHIcXmwA5
nnuKvMbky8uKO13bjRjDp+Oak/al7UevSZtdhQGuVhCgj986sPh9I27fh1WMhulGAWGW+Q2qyS4F
aNiMoNWceqEocHE1x41xKQLJ0FYEgMNLaRhmfy3Zt17qbOjmysQVrZWyogF4ZsoTx0YzAIC7+IY6
PQFT5RUNlgMITCWrpyoZadZ4gR2LqBqe10CYgCBm+4M8Bq9K8UNW8mez4aDF31jDtXP3LsIEyyt3
dAyTq9GORSy3JvYJbQ0+aSjP1mZY4JvCjrDNWWaUCIgoCY7RMFfZira3uePSj9ALyTnaa3UPYjdc
qv3czWGVD9ZfeD01sRTyNGRHqV8aLH+F3C5dwwGiwdki2msTb3JOYFc8Y6rYYBpYI4CU3652mnR/
4fghf3+dR6pBw+2b46BRbOgRTKUsbOoTGVYdz4blQ6aLWjZBeO+aIJfU3AtM0Cs7qWDZRn5Q7Apr
D+xYSrl4jsnGlaJG+NTc3La06wQvmZH6YUsEtjFmtqaXfgGUlWGh4BfCE3KPmsr8ShxYBjQ8WC83
1m5rDxqDtQDwQ2ne8N/5ErLyloA3OUl7Ew8eVzVALzVEfZ9EmSiAljiw/DE0JGVWTqDwc4qQUvZK
K61CX5YEpdoYUDejQ92P510i/8Oy8+W62CG5k4brXADTHkn237KsldPqIYIIq3koJvWllFwHOd/S
yAvP5EM7C/H572SKyE5QVsfUvj2pTr5PwSTENk5ei3+n4NAiBCWXshn8hD2fr0cDLayJwuIBc8bk
M3V1zU0rMlw9PC4lKLa3lOj6qbpghxucYfdJ2LZjppJyss/1hDnD+uiQsmYlbABarG256sao8ZX3
+gAU8mM4R3qrXl0jxN07nsYza2G+KxHPlJPb5bB5gOXxwI0NLoiRcDqEWiEGSDLx7FTF7lZa6sNd
f8F+STY0f2g7nLQAjPSuITSAeDrGLKCx8UJz8Q4bXGkYkwktKCt7utb2d4rddPhpIGVpVKs8C/Rg
vJ4ZBN4e56WO7t9ja49128Icv/Wd7miXZy1e+1ZZWgWPkxmcUjZec/6ETurBuhnuEbP7ZXZzn6gk
Jt337ZpTK0lYh8kSfWMiSPRouO3KOfGpzYy9X4E/9AziRDLzh8Wi55rN22J/rxx1ujAtfI6BMfan
woL7wp22rkjOvNTxCOPGDUf8v1bTlm3R/CM4RAH8wKi+lhq3YBS+yT4P5LqwI9tR13/nnA9tatQK
wuphbC96LBEjOPc6g/nTVK62XzDd08ekS+jHx3RXa+Y1VHhZ5ehf+3Y3HHN2wkl1r29eHXXAYWK5
+qGIiAAsKl5OdGtgKmEO7tLK/Hts60uQMZQunghWirMTXzONO6qY7DvfjPLZZ1Cb4P7+ICXi1Uea
8AV4kCqDA6yG73LOR70bc6/a+wk+rWMHdgTgHjXhB0yRiabXvNAQvi41KZs3b7pBYTJE7Ldt1Owj
GNIAg5d9SX+GHsRgZ+zhMF1pQB7J87LJ/e1biZACoyLeVUpDlbFq0iMYsFWgPdrM1O6uB6etao/X
nB76rUA9mXnqRybzADsAtBy6JhoHgLw6AOQanpUT7T++Xm6G3OQqtvWmNdh7UhxUKD8dJWmzdOvu
WKxgvfUZfgn3kxhIrvj0/AAfCYBOIbpiyROimnIAa+VUuIP5baGAvwuEsjYy3KQzNJWICdJr9b7N
XEdweulOY0XVtOOQu2AQR5BRNaWcUkLm2VNbF4nMq4mxjfiDpCm8GL6wfKrOUIZo9ZVcAo8JsQER
g0SSUXHIzErI4+yDufpatXC0JUNPA4Um4VDf7/qEK96Wlr5OZDdDIB4vgTtNtAXTfcNyb94+Mbny
PA5mwSV+teHp2CxB1ilGrQQzhzwgVxGa1lWwCWxxEwlf9v6d0Ao1S+MUD1D/bU249uZth4e7lnhG
AnXBiPQDqiSp6pKmaar933lJTtLu69bcnpWsJ+X8pX+8D6H5CRQkFecm6wf7ulR+jiMp8kscT07P
lPXCWYwftuG060njnzUyqIp0X2Sf5d3my81aHj7ENNiUzylG3tkTjcW/8WW2XDBv79zBSzBQvfW+
OoG21uyrn/vrVh2rh2nuBnYoi1vi+miGJ3TQdgncIhk2ketMQ3SMVqqqADs0slH2W+2L2Qvdw7br
qkrIWopvkVxWXvn0fr3sM59EWe16N8Iz7MQGCQ75Ir0ytXar+GYdq6nhH3hkZyQF8oq3JD0ASWMR
Ah81uOKzXoPN4Jbul41G7bWsB0/y5GaN482RcdkXc8J0y0ZYRt9OtetUSscTgwZxKcDRF0jgqZA+
wEfwZqwTSfmbZB8VsT22Qjytp30Q6XYSdJRr8YKisDRhoUTunyvDyPqfbUpa2pGfhaXJ6mpJEntw
CQ98tCFfykbe5r8zr0eAJqcmU426rP/4oBno+xjARTTZqt8ohVdjmjmbFb5O3+Vej9v49WZjmIyc
/cK03kw943cntGWv62s4Iq6MtERVeLlZ2mAZPr5F1N+vzLcBx3GgFLzqcUtZETc8l3yhHWwCk6Kq
xUUsTWYKxCDQ2Ku1k9Ic4MZAJ5LrMC6KPJ+Sm775Y/A6xa2ydeJRfEFotdd5Luh4oSDYQ4Fezf9o
qYy5Lok3m/fTJczjJc5uN8qddB/8GVyj5BAHw6mqjrAzWu8gact0Q/7d80phAv7bza12BdJEpoio
4CsiZMMl7MRAzscUkZbZQA1LTDpfeFNoL59EvzmbUfYMi6F8QwrFL4/kciO9NYKnMuTV5RHTbkBN
6E4uLf5aR5ckfiV03H8Ou0DdA4y2uppjwZtpioYt0u9hKHxyUD0ctydg0wftktvFkLF61QYuoaAS
40p25pwqJkk1ki9MzSRDy0wqOZoUVUc//EovpwFJPPcPUGncSnX3hEFjZnZWuJCfLksH0SekmmlW
s+SH1X6qwuItm+58GIBLGh1iUw0BT1qF9CLJQGyxlNqQGVbcQgRuMf7tTdnh9kDIQemLbG03/WYE
i7LWw3UGk3L9J9aEmmjfrZiOiEF6oFCHdWOSMtgQWraVdRrXqYxC7pngxon5GoDw3l5gfiGwDyNo
xWh0HhZc7LJtYxLREbGvMQhzvlc6aIkUV0s2idCpURulTwaDlxo94758OOwzxFGaWPb9pzN4y3T5
/+djdwTl1HPVhqoutzwUUo1UqPhjacMpUACw08NksaQ1WqJiSdfkov3dEVgFQi5DeJb0ArYalQfH
b2bacvmKe/9Vr5Ef6GnMYrvL+LUkWqgULXPhlvtCDh8c2B1G40aEgwbWk7y8+2Rq4Ba9TDlhnuVj
PLIHhfLjHOh64yDD6n+3rSUzUj4BFAbm10q+HVTXGNK0Wn0mRu2AvFt8XFaHOiHlsy30mU7rXDbg
+44lwhD8ls8nm6pVjla1iWBmBillwMAUWf15M1ryLG8MsWM7iKyV60Q4tylwKywyRvCGbJgq5KaY
U7/PLeFmblJ5qcTUeAG5tjAnzrHAypmZc0PKNh+bdrXnyNi9pJskvy18ighzRfv53g6M+hNOJen5
DW/DwULjqxteJc4JU+1uEGdhA+TZF9TKqd/sK/Bo4iYC/ocw8kOQa8C9bXrx565jeutpWPy7u76Y
93ztKewux4ZorD6mF4PkH8KeSMWzAg9DUo3u03v9IqNe6Nwz4wjePl3cTdbKtC4Z2pmKoqhozq7r
dKIlEvXiVnBbd/0Xw2iIeBCUZqpInaxEzDZ9WQNiYnAjhgNShJLuTtreFhnLDZW6jStOdzqZU3vC
OZ27z1T0JyJnFPJN7+CR7CM86XOCqCbWvjdplcxRr+ZqP/Bu/BQlHLcU66/qWt7DFnxJX44GFyd5
nDz5JBj9WH/WJobGulwCns197H71sthrverfZVbLG87MmtG92YOLRv7NZvHNqCvbAlNSdN6bq2Dw
mY38ACi55WC1KCdLHp4FIQUsd48AMdlexhKnb7xXqugcZuD2L4tkp2B2qe+cOTflFpbHdgEJ0bHD
jmosZqUzi/Di+ydjzhsZYMRWFNnK+K8HCFsMXfvKUmE+gc+zrtYxRJCuX+SiTCjHRiIZx38fjlri
fwzmghcZ3QY/Pqt6FU+Jf+G96SYW8e2ZOyLPmsZq1ZnWWKqs9eo5O1A2vzdEj+5P6n8KftgBHAD/
3b4v7dDEeRNdqPW+fz0DczU3qbCCA9gI2H0B6yxVypf2+6xHPzz5BGuO5nfZAj0H0DIAFkDhjr9J
ewJQBBqKqGgeR/GXQyIze9in0h+yK/WPWjmtGHViFCiLJmJVoQSReN6C3Ig4hkgCpgwT1nQyl+7o
QVse+D9YEwjGjeuXBamyZ0kfXNxVyOmTnusb7i5+PgpIt2J8A/YEVIHB2mv5HIV1+TxlPd+jZQ7b
HOiifebRwSf7iPF0YFi+Q7uQxT/Fe1ETuKy8RwH3dGLK02nWDZF9xu2i+DONn+yIivfAv8licGVE
corZuSNFVIvTJ2Zbb2W82dCXxzqGdOWxbpU+ScyOlYezbfngPafoCDtnjOkJJ6jiNIdyY91DWSaJ
IZwpoUdk757PEiAiFKhpuSdqjFyjl5IOVk/0i9Kg46+IZILlqLrdmcU0ECL38DBOSt5Cxxm0mbJV
x69WcmvurnzwkoyhK1jUzotFO75J+nfInvVfD/zQdWETrKF4fTf3le7anTBETMnjXzSVkmLq0zmC
Wfb3UK/j/6PXo4o2Jf+DwiF/fxjjX1zlexL84i1g2gLXuGf5zAWU2nlN15eEBUI7iyTbavU4danL
mxPCQAfCazEFyIdtJQjg4uVXYuoVaS0XQx8nHRNp+hvvJ8hvaJWmKW/+WntGuqW5lJdh60uCGWTQ
0nazvaOErzLfJbrYlIiChosFeS7VHqF0a/NDafvohh7JGtEGKaNSjVRPiz1UEercNNMvD2zkK1H/
sh8ljtEPg9Q6HsnnSt5L3d0OwkI2S2i8MCJaZViwqG1DMJRhKdOz69fZ6sK2/uh/o0RajThAnMly
hbEpgfml5ZvVw60fSvplFeg2RMnYPMkusTTyedkrisUvKNh8qbaTTfPrI1EwHuUgt1h9Lo3EvFh2
H45WGsVh9fzl0xEd7J/FAaCTF+LEuhYLKXTzbXSyK3i6mvtC5wax6OSdrsBTBN1EkCe2HfVfsYty
hFPJMyA1lAXsq7m7AGeDu8Pix2HntOTwwuVl/lNmBB/TEek9+9vB+wp6dwzYLD1k7yeAJkCEJTyv
W6/4KxbQURpDfPUnrBSlPpeuFd2nCeS/DXTZbE7LjNTj5FEbD+LB8o5SyMMWwPNhbUWieNE6FHuz
KkjkmoOq4l4ocgT8WpQVo3kWwUINT6sRaSgyYF6PJwwWJp3iMRQQ6rwj34DWmBgYem6rOA+1jEFR
wtKNtFtVzi1L2btwaYv6QvhDIWYgrlSEv8JpbAtzRz6/S+OYNHqVT1wcgfLvDGtqVg3tWl6m3irs
Yzbstn+aaESRidauJZFL3wxz91G7gf/OUJeHdQZhqjiwlcemHr+YxGrX7wcPMXYPFuhrZcPXAKQS
rsD7qJPiOqAtPvY8U9bzyNFEoyv5ZY62y1NgwThfRiyRPUNpsRvAzgyrwJlNsK5nqDFtmM/IzOZB
KtRes+X3zQK/dhT3+rvy0DcFFEGoZp10LxHkSljIAAFfQ/AjOb4J2w53Y4lpIKfMb3C+a7JA9lF9
LKjKqn9VceCvfl79iKAFPwxMbarFFnzM9mATE586YKhLlSO22225VQcYxOtPmd+zLadpL4j8Hoof
ACy4M+rw+fGPONjQOUEsmI12DLJ1AYZBgwhQpH5uZ3LD63Nb2paGCDw0YLDUHYmGqaI2zrPftvZv
4Yi8q4tgmanWT1Vkr5whRX2jBmZGOEhMFzmjwW78LqM04d0DzNieWeobcP3nZBDK7iB0sh3yA9k+
W0NxAImBOLCVGUD7hCygsAV5nBoCWt7Xr/n1c+1ggAWoTyOKx9kaIIUydLJal4n3prok9t6YzJnz
qcdApv8Ce5OUap/mHm1z/VN7eCcvcrKEZNNFffMYJL9xuy4IyvEvmfA2bmuPAjF/kRtykFHoulgz
PODpUPXPyDXAiIKz9nWLHngcUJ2Stn0JT8jocfRglGmUxgbXxY7xg1qIKDxh5iEe657EWYwArxTP
9tJnTK/ibjdTpTan8nYijhgUaahSS/n/WbGE3YE6INQAgBri21MEmLQnCtMv1cIfYbAGgbplk95m
MyfbIfgP4hb4XmzLnEqFVJ66hgstxcrVPnK0fv9GBVFvWKPARV1dxWMfQ4IHGshaoT13yviwmCpX
DvrPq9RmeOXy14dIu12h+7UrC+jc848v+Of3ta2sKNHKqzyyqSSEs3nS4sf6uJY38ClDP2V1D9GB
QkBo2PdbcB+C86k4/+cEM+bn+xLlXPbw71375RA3V2Ept6kNp0l8fYx6VuoAX0QDpX6fD/7F1092
j5whwpV0CCWsAbxjyLHnM7w1ratYOQSihGqupRAv6btsAsrsGpUF1syxSj+xc4EHjyAuskf1AeAU
Ve2Ad4IbhLguMQtinrLjIuko/HIjI1ut91rvdoiwtPPmEFTZpLhje2kpnbHAMptFPOcq+22Vq/kW
38BT2TC9qJT4QAdB65X8cLm5gug4VgiSErDWyTOxcYrFzvx9zbgjKXJMCaZCzJxGqLynstz1bJ3i
oo3i+VFRT61k3JEjzS/Y7rQNm1QmTBfhWjy0SlBBfcKY7fvdtHkRIbHAK+BoD+lPdhlWrzk/vDfO
1G1Tz1XCiK0GqL7rFXbyTWb86A4gsBmA7alij+z38AFjrD2tQGHGE8vNTZ6EwH2bMZIhBNpwz2vI
EPz9qi5ehDW5haXQ5ucNx4Q5vdNd6BeysdnbtnqOn53bwVaMea+3N8Z9c2UcYzFrhyL1zzd3na29
oiL9yqsh7JDgjY+EaIllTlpiFLBi9iYiZI+QW0qP4zgwCmyyP5QRS+bDYB9p+BhSF4UYsWa6a4V2
nTQFFnvcS52aPCfZdPONmDwdgqHGLmzCiZ9PtPPYKG+YHGwLlv/GjCa1kcmNIF5hif7XfPmHopNl
402hbpiWAg2MFK4soSYnJiywXJ1ZlhFgJd9cZ8fN6+KpLK1rAMG2sZI8d9UAJvi8i5ftQ5i7IIbW
iVLMU6brxh5AOIjVNqzXMKuECuTNDudAvxSIqQ9nlX0/ZVNMIEjja4Gtqw9ZsZj+jyzsYcU2VYBO
aWiOnd2P05/lyi+mck+TdE5I0lP6nlplb+difZt6y6Hkoqu7T1WLXINndaAHQaK1LgjgiA1s2IGW
cvqfz46HwNc4+2hM0BWfhAFx5d+n6N/mYYe9xwl2y9MdOilUAzFTvX3Lhq2vnig/wAoQjNiiRaAV
i+vxdsJDnEN8CAg85ShTdkve33tDUVS+DxxonHoUuxaleT1zK1PEVB3ka8O2mb+iZYI76TzYyTAj
FWLyVpMvS8y5MRJmUamKmL39oDpG3oKzQGzPcpLWwFSh8bizbojbWtBehpt7cdxgsbtqMRMPnvBa
3ob40Tf1Ts9ZVwrLhJ2qvn8KBokhcxvzW3FGl9ebJfqZbdqopZoRSJAm35lcE+M2SpEWL54N7r3B
rRL6gTxB2EPnqBj+HyAbc8CYRZWSsSb0TLw8vZiMZJZ3gTuKopsYrne4zf65p9msCZb/yPTLrqTv
8df4KTjH7mokJAfKVVuppgwLbjWZk6nAvkIxqSMRIVaDaIxLpkkpYO5m99yOJFu4RsMuXzXYN5KG
C/7t8ZU/ID+jutqyN479ve8CVlqLGMTTCKT8qa3UsL3VeEhSgt9wIhcZL35gArDxoGns3dn7H3Xd
BPhW0ISjoXlA4d0HB5pHsG0mTrBAgLOzJFSwZnVosI4t1kH5ceGpLCTstff5YdWjzMY9SzFvIsTC
G7zTA5E0gYsfui/z9qhYW56esfca1mDpUlRqIxrKeS2yRQiL4fcxUFnqVxgOy/blFUNkK2vyHCe1
tr8KqWd4Ih1t62sH4grE1Z0MRv8fsGceVCH237OdEtnsPqSlUMAV9KQEirC6KWtomIASLPYqyXP1
sdKhLWdqcjJi73ecPA7mUeiNXFxHqFiTDAJd/MzNVUnhOChb7fLzE61vtNomEJ3SfRhGhjAzwscr
4JNx/XvQULHmzSA1Bj3yIPtBvGlbuzmTbFBeduUdyChtVIoTa/1XslWHJEKb62SDEC/7I36RA+W2
MkjAuob1O98Y91DafDzQSDC4eu9pu7skhFv99GfpC21/HoyYxfQFtGB/sVPOhDs0d/PmrKTwy2u9
/4+W/D2HtS+jIQX/Tj++Ky+oeZXENJzyd2eis1kgn3YXhTuLhFKuaQjupwY086VIH+mBsqaFo2tI
i4uecBYs3n/S06LY68UH0e8MvoD7mGeJWXRQEl0tIuTi6vfyK4o6F5DZ1V02Ao0gFH0KAXD3Fv3x
w+RrUtVH0JWzvPvmvNRAtjqUqUMhbXDqNJL7Zb4ajrdUMN+AVariOGlBNIcNWpvZAj7eKyJfun9V
iNng715SgW0FvsmffDxmsLGODfy3yfJqZMLwcbBT3uULMPq/8dffAjMqwwDDJipGfXzn632lXcNT
zeTqHMKWHMQZU7JUBnrPI4mbpHTT6j2GSglCE4+Pb1uiFjv8p+VrnYndR462HdvUZGZYCGTzeu/U
Ufxc1Ft2T7XP1wv0qehmBz63KZg6q0b5qlQhdKfLZmvBzFmDTj2IvzZ8+ti5XdrUIIs+5rs3WXtK
9RV7tBdKcke+8EhJf6l9g6g4ohxV3VCtDZUP2DxZwf1zgqbic6P7wiT98VwfdLibGv8aD0Zjc630
4i+HlKmwxkgffJZxoCVve2ORV3fyh0rfftt/1OKtujt11eOhF/uJ5RTLTPCMHOBHoX03FBi4JmJs
Nkgk7sta+Hzb4lMrSITheRXfKkP0uaYMiuFxQfenU6CPDYvEbUryHeK8zUorvq0DjZ5zkpEHKuYN
zP1uekUqGZafD810/0/VyMq9tFzEDw0nnuB9TGt9sFKhCoibEVyN9UiWPPoExBOaAAJPwbJr53v/
turG+6zzz37EWOrp9+XGjok7ESD5SZeYMPwpYjc4HtlbmDhIx8ce8Whu5ofpTask1k/KHo4z6EUz
hue1K0FXMghq8bhrouS6iMx8G36Eieq0SoMERitf7e/8it/VERYEXzS3L+TCGTrZ6dsSCt5SwTLV
7PK5dsRrO+/mCqh4JlzYsDrlQXq9ylQdP+k1NAvYH+6nioGrkPDxwY3BywfKnw3J+5Fn7mzyE40O
mI4LBW4Qe/tKT/CPfaYKEotx5tPCjI2gI+Ym4fK20NzePTtdPLLqsPcSJpJTtoMp9qR77/iVWqIS
6JhjXXV6DVti6VmeJwWxlW7rcKqeEHkk3TUcFdW5iFRiw/fhsIi94c0RG0gxxcC/A/s+d2QD7CQG
qXlcK0ey7yOU+UuTzCDNjqe8YNaSCnc98JJxfCtEm8zvB1HNcYNLXYRp7gXhaKCdXhZO4yGCh6VE
IteJgmBTdBakV7uCKT8EragzsJzoZDsZas/D5ZAnyBRTl2UD2rRNNrUtuJfX8PLd1NB2lqOE8ljh
tw0CRrCofRidrjtHggUkc6A8UiQwjXauBxBGfbev6kxXYE5B3L9HL5yZubR9TP3iQNOT7MaRUpXa
1dNyBbZSzbiAkzq/FxLvSSt6efzV8AWhdginML1ITpoLwc3ThNFPGyZ9SQJfBr/52oOqz/5Uy8aG
9Zyq4/TUuQPQKJNY0ZZuYU3xF1JpsxsoePv4GY1vA45Jzlxbl7dpwGFy9kPaQafE9KZuq3I+f+r+
GiTEYQ6vph7dyPoHj/Mso/JYuotlPDh6nqMbtipIiW0dsbbfMVpctbTJD4BhPXGQaE24/lts6lhE
9Jhx8oKi3XOcGafRrIOjpGSJGnp2PS4UlKmjT5yPwDt5Ps21Y1ytmCokMTQ8Q8KvJ5eNJhgBGSYd
/ubxj2vDCBta1xJKr033EP5Vlhk9dmt6teu909TNkE65+Mygxe0cwwNHyYyNMgQZYaKOdMsQQdBy
Wpfjw5A0Bho6WqWv4FIy3uAGL+icpZfinBL9yICX9rnAba/AOs2v7L5U10cg+04PBLgSDp35JsVv
pneQREVD9dMVj+qUciEwFGW4M2ZNrt6mw0dvT3tdiSbsjN7ykQ8cH5LUnAvy3nQ/ZY8+yf7mnBjO
MgjirBrrNmQD4EqYWxlE1wSC4zyxqebCNR8gUMxvDpQRQGKzE3zl4u+Mi6cZQCNCxnLUuuNkhfR9
QkFwO9h5ux91/FZRF8Bh1YUFTUNM3EYot8+KY+yW15uAe9CuP7ZRvJ811hkmTA3+/FY5aCmnVBND
ApFp2Grx4x3p4DTF/eF9LL3GUBBaASsawHeJpIMaOytMh6N8FWG4OO/noQVLG7MsM/qCx4fYrHHM
FIVdXLM9uOY2AOZPwtWAI5LpUonLjowK+y0PZeS8zKYr3zmuoyxMXrvb3QZ62Np7KICAPgR4HVhl
y8xaW/Mp84NkDXvL+h6oL+03z9M8BUMqojEZYS5TagfZoePTmZm3teDie3A+hfm8MIo8/63tAAlQ
HW0JZdQmt4QuYF4nJBNsJnQCEDWx11jV5Esvr09WYK7KDEsIcL0bQL5emy7kOY8CMKmr2gjllFDR
HzxtxkPi4uaspNy+f1ZFk9ELj10I/RM8rnd+HgY6mnVLLF9ovLiw+28vzPyyrnhE0ifmsRQvOQ4v
pZYJrYQxEksPbOAtsKGXPw0Ekhud4KVbZFxPVwJk5ZTocz8FmIM+13U64gm0bjeWxr6Ld9O/YWCb
JKx989dR8KDB0sSldTEobb+iKqP7K6W/cC/+52AqSuAbZ2LXKMtqx66iMw62aZFawtDf1EnHGTdj
REFnLbkqV0O05uP2RkOWEvv4azrvM1txSxkkSNRNBeGbYE3RPf7KN8FSQ2DL1PJFg8CCjYWSvsH7
RzqEu+MjZBrl60i23SWmJ61No9hNkfW5TK77H6mbRgzYHeaS2885WqOMcqkjfdf0ExQl2VnYkyu8
ZrGUrVixLDaa1yvyoZWRlL9GeXpo8TyLnwAhSh3bJiNSXQe9kCwdAA4hyPijQhZVCbLBw/N3vwLG
YBmqJUNyoJk6s90c7BCNWbvYMBAvxfACLGHeq4FKjDiYfhAyfVs1dwjzoTgSfrIonX6aZ1v/JCED
U34CoZUgLee2Gp0CPAE1FdbgVHrF4vDaKWesluFK9FhUsly4eP9jeD/uXO4s5z7F2JOAiyn+XDql
y6dGaZUQrsNrRYj8nGgO3zswGvuQxHi4fM8UwvCxjfBiy7xvrcNSL6wjc3MUCAwz7YCXIPusDERc
/A6kd/Lw32pTwPpzS5iteaUM3rau8R4vckiL7MaMxTWBPz1AWfKza/pIV/PovjtTwrXSAQpgZUFv
7/ZvhHrzozHHkPeRzO54u6i2oCEAEwL87LcBOtYdk15onNLcF/Gi9S/V0udPQNfI4yhhNEEJudl0
Nl9Z3w25qoAvgPZZm96GREUQvrxN3oGE//0O3Aqaxy/Sh+L/BLrpnkCfs2lfwP6bn8NFsW3qtXnq
FDxeaMTq6/m7Th38NtCU4QKHE3vBdrl8dvY6mE3VpYSx3zQEB2Pw02pRnHJIXNKtYb+rJd0OvFPn
9ophpggVtQJnMpkXfRn7EpVfVpd159vxvqOEglvcCR2jN5hQ/dJVIUmIPhnJJrVe6dl0fZlXpP/0
wqM0oDAd1qddPSC2PHv+4ZnkzjgRVR2N6kP4slEqfUVFJpa1/JJeyH2svwEYEuLaF0kiY6g/5+Qd
KqTxSYu+L3QuDxmjNatXUdZ3auBEaBoXQxfapkGn5PDVZQ01E3vQJ3rlhaz8Igc7AVuJp2WPKRXH
NIIgLUeNEThohIaC/epSoIJZXly41Eu/7yo9F9rUEO1navu30JwD0Wc0a4ttZzojaW/YNnIRZS9d
1lKekxtALawlP5svV3hitVqEEZqb4ECWqurM6qIuPab8p0V92ZVRj8y0suM1aYkD8swkPDI+7jJ2
+pk6iG1gRb578D/P+jso5rw209KpwF+0eAt40BvdDQvpR1xuq2UPTzRxWvz+J7wVTTMVuGcC6uOz
xpeq6r8Hnx+r08bVNnH7OX+g2HeAw6upp9ARsZzBjsooTfPBa2Xgkn3ECOZShWsOQt2XlYkAon1M
O60MG0EWYVgEtXKJfQv6FW16CIwVBJicZKhFQg52bQr28vmoPUPZ8ApDei3Kgn2hWMZMN/r/eB1R
B7yIm5759NXwrg6TyfIc+4qK02cOFRlRAWE3cj6/uOqfEiNkK/kbrPMBkqWRErUL0RCI/Ug33WEf
c1aDSX0VO5B4gnl9VmV6Wxdu919y2ThxDzQHp6OMYkzm3Kv9kaGaVq2CODRHWAgqc1q53RgDvsLs
9RyOa6bXbNo0lF/Hh4ESdZd4BUvKB9H1yLGUP5KFDLnN+O/oiTP9Zovk8DAtpK8lcVoXOwwKDo1h
1ytCrkdqnegTt5ALdp04Ne8i2paM1IOmjNgXdz5U+STzAIJXKnmsBlkhCjF3Rq2XDDXyyUZ72e0B
rIKW3NZ6m5pj+2Umhb/7xU3GgWV+SX6htTqs/yJc1HYWcFK6CjaaWGPHYGxF07IJqHg0479WBEsv
W0gkdApNvCsjlsvVzgksMigfO2Bb04M+8KtKjAC3IZjSvRU92I1N7aO4rG55eO67vequmbGpQo9t
ZOYmMZnXHoz2k4IpeVArA2TteDNH+F4o47Vpu9yOS8CftZJduClW2XRY10QsqUDIj4+lIDc04XLX
MRLU4xM0hlPInol76A7y6Ztzgn1da3GDlMOINyOfTj49zQu3tWLqu+yB9SwA95xEIZOYfEMD1en5
xhfvErs/c4kr1F74DlsdelymiDynXC/CuTBiCO/HTcyZ97g2WElnPc2UsH4Z1DAGnAjo7RKWRclo
MJYPxol1pCQDOor3ufecFozskPZ/UhJ5siT/UeazwMX32Py2OaG24TcEvmMIa5JRg7Y4w+2T6grQ
90DE2fU8+3UpUVK7XdXe1QXpHNeEnMl4NV5WEMyGWtCs8iyF6rneZGYqxDnY6vbLZwWXw3+l6PTv
e3E/mGVIIOH9VcYx/yUiPYKWXcqXDIXg8UZSpA2aKcEK3iwAq1DvyhIdNJg33tnlpQxdel8u9HaQ
g/pQCSHoM3KLoJIsq7HgKrOrbaXRhKbn0LqCnHw8nl2y89ipRT7TWBilEZbS5K8i6/GqG7qgLEt/
B65z2S3sNvCuNGzvlwnX9WX6xp8angPplsZUrEXpr4RTZ6VVTOML4PEw4gb2G0HIXeLBZMFP//On
NNAHZAoCZOqzNEGKhMjvpGswK2pOzZMPJSuKxRlgUQZLtBn+LIQzixOqtu6N+yQSasfvvXMXSzGW
0ZPeA+zh+cqVg4iI/QEFJYYSzYJs0b6Ed2AWs5hdAjpaPlLCEAQdAmVr8rjVRifh5G+hCKs9ITqP
ABxhNvCm/lavHzM3eCuEVVO/aox1a3pnNPWTsV7rv51/a2e2mkzLB85pf5tG5c5WKAZXbXen+9Ea
spk2qsIHyiAdRNu/KFd/2794KoFu0QYcjI8Z49wL1344V3sMjSXuKgyc3IpETtRsLJyBqpQ7Vthn
Wz4tj5hQploRdDklLtHFbbnsk0DzMatXFFqK6GPX20FokeT1aSj5ei27RYwiIlRuzc2PyBh8ofsy
HnP9uIcXYxd5u9cFaY5NNYrZ2IR6YMgW9vZxOT2Edmxxg+oHQgir2zjHTaw5iA5H+XTTtQXSJ4Vv
qH8xkRkMXL9p6uXrfPXFpZx0irETc219JyOPid0KGF2NrTQtwhFY/GW5skm2grK9llJRcQjAAxcb
YArqAkUd7N7+ykwRggyWsAQoFmSQ6G9JDTgIuGFySz+0JA7Tp3JL/FZzOFr0tQXH4BMjH1JWifJS
LmVsofZycCnty71ZenHLIDc348FMU4q1K5PkX1SO73Hqq05B2yP9xLYNeV7K40b7MeGFEW3zBPwP
nKzs6K1y2TR4pboudhhvHBXT9urRn2CDmZ+0Zs3fw3Kzl3YRbwr5CHRAT+Q/rBkPusSBo2C15Idx
hT6Nf4XPHN6e/th8sgXU8CG0H9S4DxfYYCRgQb+hUZ7+DMWkiJI35hy7mKcdN6XD/OprZD2ObFRv
nRWknBHRuVHgpNnBhJ0EGZl4IjCqONdeeTm8p2pV6Mg5IYIxpMdx57DlBMxKhXNhrLq6izw+QsmF
N57+LMUqRRsv/LSbyInJ34MeBDVzM08YMUrkYQ1j1wQJk7zmnKB/ED5z8nMm3tA4A58uRsSGLhKP
5zcxVoou6PE6SbpouAR85xJCjOvDvLgy1TQw1AhLAarROO8aEncjnfcObN5HBbCGkEsLQGc7EgNY
f1JMOa84aIwK1lWoy/VcCWqMRQNLBu6G99h2yr2QUWrG2N/6+LRGaE7sVNeo+b28MIX1kwGg9Crz
6goaUx7i6/7glA2+wJzc8VVyLh4aR7UQSWmedmIrmz+WiBysBTFx6VasGWvvkOLE+IrtPLzr4L3v
/ypvOAJJkyxZHDovwO4U9xKUzL1qOdEBJAlN7baaBt3GRz7Q+LjoQ4ZDFQNm/TiPyU7PxUePJ6bd
MtRSoHiP6psZ8VwybpjpixcTkMGtgGNrGb3APmNy5jdvtKg4sd0JuHTf9scktLtbnp8m4R3K6rLO
Kdm09cEISHv//zWl0eUcMt8AF6K+V4c8tAGb1ZZ7PNzxanFOC8vzUageQVeiqrRFabcqHnmYSSWe
bgH62q6v5L7HsOyy+7bUbWFJ7sjKTq3f8QcdCWMfPpXp/CmOFqM+3sHpiCUdLPmeonZ9PE+xCnMv
mugw5/seA+HOjKWy+aSJt7yX2SLWvRSiydyb6T4FJssRlBK5r9n8IEe/EYxI/cdJMYXce20MfJUr
dBvvrHHkh0+QPegeAbTPXXq4ZCCBfau7Ks3Zgrhi81v/04kcY/uSSJ1onHAhoaF8edCLRP8onGZk
JDCX18026e6BaNb4DiLbgXkmIQvvGGlE7zvWqTqXtylPuzWkLoHph4mdhn+NYp7APRuQi8E4jcIg
BqVtIoo/MfIIm5FK83vmngKEjwumGU6WmL6IdUv2tsG8+w1Mucc3mrf4tvBP4mxmX5SaMoleI+vj
cpu1fnWAPC6U8DfqiEKZM7LMoBZhaM4jBVQ146bhmxf6/qeGedfG8oUDgXoswWes340KwE9swwPD
pvI8lKIeEYKtOKX76+erd+h0zDlXVTeW0me0il/GIO5R2vP21rinDCKiESBwGgTv7NFzGoVzgjb8
cdJzWsJWk5oIN391+UkAsxGdWqsNYFDyGWMG6WevrORoi2LVx6o9+GR2U8Sd1ZUOR4WayGByUfIi
PKXcgMG95aVE9e+I4AH1u3zbunbqZiQsxVc8LlJOfyLf+xFr5ro7hf9tCJluHz2oZk7j1m5EmOlP
lGT2TSEE6bBnObxZhC+Wp68bTgJbXkbdYisI3I78sk19ubtRR+Bd5LinulifhwJEa5V/6GTb6TzM
yqPPOZGPDdFJ33rvp0HtNURw3lIjMMqWouVs8FOmXg20AqNCsGcDFhoKF6FOAwhK0HxXvISe3uNE
/yqiyP0Ak2hJHer6/DiJTzNwye1+1Qu1E9lmcfYW4nTQDa0uiM2mkRJSKRbzwsLGF5+kDoQJ7woA
71AEBMEd0NXwuGNgFVmkpgm97rt94KdBbHhOz5/g2MWsv3VstEwJxHdV4Mh3DbGT6jBeXDHhhJoR
IaqSn3vbV5loLrZnO3iKEof5yiFJA3Q6fMWMdtozLV/NAaoGt4JJKDaJ+JG+JdDCSiWaluQXmtns
7OyD9hTL/hUp51w2Ea5y6YX/fSLKV9tAMlr49RPV/5u+ttbNr6iKOaZcSk84Rena3QT1f1AnDPc5
o6HI6S6Yoee3qcaSUOTVh95UTGeOqPGms6GqgXTN931y6sGGgFxuEQ4R/4Xovng3328li8rllI3V
Taw7TVKEKM14MuhbCYFDYiFFkm7Xg9t36U6S85afQEbRmoCnzqXmw625ro0Uu+CixbZwxIPpMI35
GqYS+GN3vCIqhYE0nFuDOauhXCde8ALCd0wCQOJHDD8IswBY4RL+wDc8WPdeF4PHvTx6kEO7a2ws
vXnAfLEQcToo+pppdeA3WBG961SJpWq7aVEcungf+hfoJk6t65Xn87GTBm1aShHGkdfUH2JNv2zR
cCcsndWhandEp2VJx4pOITvYjbt694ulLQy+gUP6T1iFzS8Irl1i2Bf1MvZCZRzOsqXDQjHOOBiV
X8OdXQ/4KAtO3LzgoC2IZlyNQvnQV3PGkggCMH+lUH04t/Y7w0GqKqgGZ26oqdNxHyPTC/rGnfxx
X7bB9Hvu/5ImHAu/1oTAKWHpXRjbL4+cjO0FMYpyd7Ll3f9rUoY3VCEgwpbRFFEAqH1kASj/tmsa
5alpHK1z/PHJ0t1QXXZ01AHwCeVTrJ17AIPb73v/ZFm2EaoU0tnfwkLcfU20wNwh0nNRvl3am9jx
c/VGe8zVzzU/sE9F7QLYFDBaC4grtjSt3PTe6i73j/eQBqR46CcoYnbZGIozwUcCQjmKVvPQ8xm4
GcVt2TxZFh1yTr4eAMsDxkqsDk/hRZAFIS8cYnTi27Everr/OG63rrEcNO+zJy3j9snC/ZSXTvKR
dh5fKV6abkcE7d6NWDQQVO9cxBtdBzSxLwrZJ9+YDZRu++7O9ium5VRxqaSgBlW7JXu9aV45g2HW
zntxVnLDPvgLkeANqe29FExr3FLtpcg74w1fzH2MS3Zc0H56tVPEQfL1eNluqR3onuVUiefYl43h
nSpreK7UHXO9mM3g5quKiRPpkEuhg+eByp3cNXi4rrFTQaJmTrVMqVX8CrYbHBT0HF/fx5akfP5+
sYsviW8A/koSoaCLHqV8c2mjABEIevDD+AAud34FQysHXYNITwm7JIJhOIwPj0Reh242zhRVRNGN
iKD/EhP/WFYwk56JozcOldr0kZbVBnG2123WhhpslC2Nmjd3dRrXBDaWHAxHprgHnaapYkn81OIp
9zxLvWf+VYDGq0ap1VJmAVmd22ln0jYd1MmaGNynO9fjMi/cAbHfGxnA+TtkWCWW+hNV+JCmardo
wYMYPxXbVk5wYJZAbNo8h62vr0FPHfgbpGt+lGcLXNmULveJS3Bi20kgZeSoJafu7I/NcdYPChAJ
Ptw3IOrHt8QZXYp8l5zyD8pb9Re4ANg5BGdYXx6Cmg8eYDLzVVe+sV6FlPCMXHmN0ADLQQPN5AbT
vIJINRUU6iZEH4UPGzi7wcd2G7/u7InH2vcFt9myt4X/aNo5V/q/2IYe9HhyK+gYfkCTc8B57XD2
ZzY8uLLqn330vhMMfgWQvQpvqnvclCmUMW5aACSEeXXHtOJPb9ZmLPCJe6JQSqDp0zky6PeIbeo0
xNV8GuFH/SNEDnn5jFEOQyLmUKKtdGPZa/BFxb4hrsYtSsb0vFvDtTzpZg0vweQZ0HeT2bfwCNnh
GBeZSa1Ipv6pskrlhom8POP/tpn9Fr+ZLJpb1Ge7EihQyWWJxBJlP1bRK9DPCDNDeDVlzfLNYxgz
Seu+VKFyqda4Gizjl2BlrzvLXMQIBE+2TYIB/Sf/CDmUpim8qctoGWGvjKjLAFT/6Sfqc6eyW71x
4PDLeu0kARpEVW6J1szTmOC/i+ym3o4iM9IgXimzNGSSgSctQAE75U5xpUjx10yn3Tixk/G8V+Ve
mykSd+zmGYiPWxrAV9lpIhF+MoRwR0IQ8c4wmm0fq/zOILi4GdPpRp8ZsEt2oLIX2vQoc+dEPS/U
3RaJPNzQvxDLpyq5/XS+Y720xaInZ0uyg96bfJA7OZBF9NvsnyQxbZL1Vka61M0Shgae5vGCkRvl
Yw3w7kV9WXnjXZB70OK1GOCZsBcYUaFdtQOgd5a6ESlFTRs8Tc8U1D6Q2buObzH6dPxA0cnlEskZ
CxtrBTBXQLiLY7bd78xGHP5WcoRZyOQvq7YbMyFXB4daY+3XuQCGbux7WFK1FqUgKncrLF3gSyLD
BMSsm+OXIjuXCegNCyEtoEBnsfuDxO1sd3g5b3LCjJtG+YtLFJdxlTzKefI5Ob7XJrzYJ0zXXhxI
fvV6GaMyxYrfW8Ywl8Svn7g20rVeNlLHw185Isxp6/7061cHgsSXHkBpuzKeO7wm5hZh0SQOoof1
BwSHtKS2302dVWzodidjbahNWz6WGJ6pvfHBU/Uytv4HJSErNWVglNEgeHhfZKCfUs/XaTmyOgin
cb9mombUf90Q9gJGfqtfzzlqPSl52FOPm6iox7lbbrKcVC2REhUX49WKO04Nv7l3l579rEurp3Ph
LsVzZfktTlvaIJuInxaFAyiMm1amj5iTU5cVqHfgrIuUQvWL7l7eXgSCit8fCTAegpT5Vwtx0ce4
7DzIuDqryHhvblXR0YoGAnzBgUWoqlMwiEsw+pNp4ZTwKjUutZ0ftndbCIY0QPoXZ4/HEpVwX635
RaSXoR0vclKSKVF3ogRDPXUTcVcRzC3m25nG7QbDqm+LRrSCYZcPfd7ZGg33o7vwapilQTRGzDpz
OLNCH9MwciVP6aBaVfZCqhFwq48bGxfFSFSwyzfKNIqj1cxXuRhHMFFss/DX26Yd9Ei8NWS8db7+
xZ0btni5bHjE7nt9ApJ2RLBMhQ58lCxcsshg76Q1emHbPuiavL2YvYDUabqf34viwey2A6weXGgA
hOl0LpMXhTMlia6okfKnhe0SU6UIaDHnOdfZSILIR0brAStzZg1/ebfSYlt0IY/HyAhnmWB8aByq
z8xUfRF8PzpIEN0T3Ze3hLiLCK/Df9nsans9uVmQZYF3FjdPkmSnR+u7pOrG2HYd55Tr3q4FSuUu
3KvqhMH3rV4THiWthsnq3LZHAIDFMnNEusrPK1eVCBX58UUMAT7YoctR9XqXE5kysnU7/Kkj4mMK
Xjb75utaZMMz+msWLxK52E7A97WpxnbiKtBBMCFSIW/6NP1X8ISTQuzIhu34nVizoHEDvb4WSmsm
9zFBMaMl7hF0WLB3XVfSY7NMagxQCuddS6OeFta0V7MLYoe+6RkGxRDOTsTKLLeWlVH0SKZeSgTu
aIrOto1bw6DfEkLM429CnqB1OyE0wNwSZO+T+zqV0zhIqP//4jTeS8+ulSxVopueiEEiQJSvW1Hv
b2wkQVj76QITqDKRsOOT/vIcaZ6cFFLtAFsTXiDbh3FdAMpXblRRiTgMivlQrrF52XpyaRlzMTso
GLvQYJ+zeTwK8l9X/tkYHl0dax2R+axbgAeadLA8EIk6IeptkakDP6DBQYb0r1PiXBE1oObimp2J
a439Wl5D12Yp81KrsapWARTKYxo8I/HLBuuSMu07i/cdDygS6nxkv/csZYFGEb34ON0wvymDVdib
NE5q9SezBCVq1YwRjFsHk8e44ikcEzBH1li/+9IpcebSkEq03XxUkCcWfPMEGy0ecW5X4iQq6//X
JLaYF/Bw7z6zUfRMmBn91Sbus90CTxxjkgnrXzL3p3VfH+wMTodnF+v1weSzrqCTE1UJoxHXWus6
e8TWhknHpdRC6VFocXxHDB39F2jKXXwLdUJ93vdklkaQg5O8vPSThHqroQm6GVX7WVY1F/CrUGhU
EUfMOKYHxjASiLQZQxgGXnxKNt1sAUveTkmLa7ZVTDWD+QHtRp4sx9bCkBQpUxGDvCcvYqmde0Pv
vw9jy+I32En8YYGwOhZn822q93xyCSLFzlcfydyZUvcbwvuG/ixSTHlxD8GfyOoobWz0+BqpnsPy
oKceLQfwFGFthJmlbRbKWr7sm4k3j0sytHSTJ4uRn6Q4wOqwewLGd6YfLN+8v21V1BtfhLrYPo9a
/W1bnB98vo00G+60U7DJFX6Ub1VAkzFpJpKgv1+MHl3k49N9FNsO27seLHDbVkB31T2X3A12s+wq
Q/Jwn4JpvIcGVhOmgrjEWLFyN0MhvVtHJxp01Uy9yD+3day1F0SmmJ08xySD3ZromEwjDc6OFCs8
LNqpwNuAihzzBjZNlhqrN+Uo1+he6qtgmU4PWPkB0ylnVYoWHZqMzLKKm9g4iVgC+pWsKxWljk+3
HB3YNI3flgyEBRCki0fLreUsk3uAy3ct8/A7xr+02mFGdRpKjz/m8IFdhQXG2whC5PIbmvOGoP88
32qQzVrp1E3XlVOfs3EaRar511gNkY8doQ5tOBKYWkd2JhdpBaY5pZdfi8XuBVVgusdNZq08bmgx
ePlujv9Q55+bnCYIhgWnkKOZpabzkS/5blpBixtuarkFOCa4TYT5fGl7i+Rsfsdvxfbr1hAlqdK+
5f1uBgLe2v2RjZ21tBr73MK4Sy5w8lZ3YHBGfbAkzlZ9An1xE7n6+3RNASBYi4Vw3kT/OzLcwLUD
SSdWt62A47s3PzL0D7VMVYxbWsaxVRK87L1hVVfRw8nlih+dCevqyQAlvsWRQf2Lns5mTdU2WhyF
vXb4dVzxrXHIFf/veYPlzT4+jdtqmvfpXwPzDuJc/XyTDJgdQIAJ9ZkKft9wpIBhvPhx3gdfQpgz
F9SgOHh5XqILK1oNcEzFnIy1ZQLJtWLrKECewEgrW7pgKcEeanQCQ0MYD9XLMUbKNEtfoZTqgnuq
OApIeaeAH41mGe8ShTBq8d5abCN4Ic0lQPWlb4dUsKXTZRYTzVSHcKtwkBK36Qa4v9/Cyq8IUSQT
SK+J6EPUAE4cUtXZQ3aVkTxJvGxAYRdwJTDuipbDugufiA9cFbxQA4gFTdnEuDeEl5K8OzMsmoJV
R+lNMNWgZwOzBDh9DnxZWYYmfkNxGyltCnyI57rw1SNGdNWg0zjS/sSw0vowI2Vb389HGd5gwtBX
mOsa2OjAvK0RFFLpuD8s41qwa+0iIixQOuigkrNu0f65VlyMC9wMAnnw0bxBvh3PjwwjBvlnMA/f
Gf3AwkKauRkcsIGOr+W6gRaRQcrLguG9/UHF1Yg+L17YWYNmTj0DajrnhISRXoWD6/6fQ5Ykww5k
ZQDBJnRPWPPdLM3Nj0N1SOw7dwqW8ZUdfm3ehpJvZgapSOW9KiD3wF4zWXfMKDhgWsxTTOKV5b9g
8Yytse022cEl1pootfbRmeIRnWvXakzPtltIiXHXEyiEyYAXe3UAGNEbL/Lc57ZfLifOQ14C7bsJ
KnLy3ryuluB5jwGmpBkEnZb8Ey0ER2U8Lrsu1uLk3zkS85yx9/F6PAjb/mzkDcZRbsUhbjsnJ9Dj
MGaIFg/xMj0CPON287hTuHn/yZR/sMXAH0/JiTYUQQlICE4E+RDWsS+rmgbF4N5EKZ6+LmvshQVj
Mgh04aLBl5M12c38siNrFPY4XGfRyKZQKr2Stc3JyIwLGa4M1nL3HGH+trF1UScl0oseFxTrul8t
Pr61zi3jiNFPKDrAXDfpZT+VRaaqYXncCS1Q01drK27gFNf0teZ8GPGQTXUPRXnCt8d+GgL8crKS
908ZBViYpWN9oyxfwtBhFtn452UpyfhtZQycULSE6MQd9ZLcjaYS0Z/dwaToJxm7bXobNE6vwq7g
j7v2qO1F836Y0FaANXskmwC0XVALSN0Tyl0xXdSLbZ07TbAQrSZgt1wrh7jKqwdrrMdOU5Ao38tn
+llRdw6e4qSFmT9DbsHGadnHcZn8CrQkkqTd4epq0OOn+xZ/Qy17WBsmSdWe+GXjY4YVB6WxBDgL
IvpDN5GMyXRW8BkiYbrboJqOkhtghBK02MMv1dlpjIYeuOhvqojiGzxuF5NPs7NL0E2eektN3chT
xjNheGuRhusMmv5m4eLGbbYbyVk+6aueG9x9gEAl/flZbIKfRM84FQ7AQdZu5dQUOxHoBmWLzY0J
UlE6qEnLkwIlJ9skzseRBbpPsOLeuhW1GFuT8rn08S0kMDo+S81XgSK1I9SWTNOKuez98IXq/cKe
gk5nSQXT1hjKxpaBr7keSeBn/SIhmOBp/zGBeyJe/tKL9RAyssQoHIBLYZPUsSmqXdP4J8zHbjv7
twoof46naaDnanH267ukOtlR3h80zWL5Sa9U2hf2O9La+426gxNST2RzcaJcNxXWGJKQndzj7my4
6V3fUuz9syOcCGZmi5rgrfN8g1bZ52AISagKivT78kchN/vjs42p1iv7WX4PX9AsDBXIyDUDD8GK
mxZv6BRxmHPLACswe2PxC/hweIDUyMtO9RKHX5Bd9vyzq8jsvZZ6gEwgUkxbdYdr6kKtw3rP3Q57
LkWPgKcZyb9H0+zoPkuF+k4bAhcnKatpj5EAn+fM6Ld6mioQOxlfbv7yn04haB/00f7hIWyjy5Sw
XCAo1aDiZSPRIpHiKLzZ3bz8cZgzhVmh1yDh3B6JfqQd5jH8yyd9g35NS6oFREObLzR2Eahjpa6b
S4b02NcovSuZrfNGTgsFtNawXryY0IjySl2GTnjkPmzUhyS1sk77+p7j/e4iLH9B9rDrs2CX+n7Q
+q0U/2ZloTQjBWDC73TEIdJQhGEva7AQEIYr4yAAzJcr0LClIR/VXhRDSfRXJ0M9Z0WbaLIxyEsV
zMFgnOpmbY7mY5BPbuu3kM8x4R72k8vhemIoL2Gcu17J5bdGmbJzh4dzHmryZ0xWtm1v+xQ3k21G
O22esSZyB3c5Hh6B1LrL09oWd+ANrKjm941nG1/9ly9ftV/wjB+ckSg3cs9ocwRsw1x4kgtwq70i
87vmJJKD5fxPGB//j4HQYrxvkIeHese9hw66oBKiYI0vt+suqjvshHfjwtULPW3TJ6UvQskwitq6
b9li6ecpfe6LzTsPA+d2GYvLz/P8gIBWYRs9O9S5y1FGSkLoZk0stvY8hvk7B9aaEMazMwaJkgot
049vInOLB/u9BSB1KI+nIp5cQSMiV6opsr2hv70L86rMEM+tbLhKcSgJ23egqHuGQwSVIjGgPeF8
2PH+ox4+qdYsyW8647PrEfGxeaJj0kFH9w6EYJ9zO3PwLU6tK7bbfTDe0ZukwwDunZganSshx8TO
RgfNG/ZCZLWebukcfEkTaRnEIiDmYmxRmdRFIArmrYKv9DWGKh34dcZRYhZrxTk144bMAceAIwk5
W56YY9Wig1o+5Uhk7l0JZNyRJVyw3Z6YBhC7NP3GiyDpnYA3db41YnB/w055y/3l6JmnQm8qAV7Q
hlnNyROngdUTPgocx0VK2+7+SJ2WGHepbbsXCX5mpYB4JzxfHUBwnseIU3ij0vIS52BqX5cdmRL3
isbfJRSoBETlYSnzCIfdLBIhPxENdHzKQ5G7uJuLiQbjLMGM+AjCjviwGMzxR1/lPU9jTX+XKZmx
gN9PY8lGsvCn7e2LhaXxnlH9f1SSjZCISY7qOH+h2VCO33VdAbgpvfcljE3JnvhqsV7xJRyXHWPr
enIgeoX2YGHphwRaP5ARWH89PFP7qUpJdLOytvtcDck5hHnZzomqa119E0sAzTtjBQlnU3B8AOt7
0jByQgpzJIOrdrq1/zFlxvk9makXeJ4ylP+1lu9kZHfATjEFnYaE/o63D92KcY29/rciRNkDnEQh
gdVMfq3KU3RTpb0TVofZa35Dd7x1RD4SXLZSrPvXmS6A3OarhTw0BYUMKxh2Bpgp7R0ZDJs8oLLd
65Yy1DCe+jYAZ5tKU+M5upiu012jvHmCC/5RN5zXE3WJv2l4Pe4FW6CK4MgPwtL5/8+wwLKTGv8C
dwNXQNEzLuNIQM6mYPJowfejpDiQWh5rT9HSA7l4a3v86CN9zTD19GRx9HB/c963qs9bBTtnOJ9Y
f51P6180bvW8qo+n9o71z1fh4irVNoOHK3zRUGL7BAdj5DJ4eTeQ95Uye5gbUxfOaK+R/QXb0stm
v4UIMQqw0C+b2OpiSskWZ6h7/CHcZ3f/nvS7Eat+uBo0jbypzaYtdjxTJ80pVBB8nqy23zELK76/
Lk9oOye2LkU4n4WKYTQCuedtZ4bvabKB8XUyMpms1SY+3MKKNTAvtBxVljndLk063qRPmqHh5Ddz
cfYELjI3/fzBbE2J3m15VwV/j5rsWrG0DvAAsf6Kl0HVdFEWWUp1K7zCzIhjNxGrhRNYkKDNzM7P
eCdoKBgvEOp9Mr2pzHJhp612bhIAmDmhdpNYVkQGhuBsizgMsMuy+bB8kh7MUnB+cx4MYGKPqE2u
Shshu8mP5UmDcVvxv6Q2UJ1IBXL53ZnN4KnOwLu59vuLJg324avMl4K0Ve0F/5VT3AOUNuH9XhmE
+1m+80qXsKe4neHr60YRGYR9h6K0rnShONC9zXhS3eKlEZVzpyw2depgsRtvmRwjKSVuqJYHnwwW
ZDvUkhCcIr+DG1u4dha38EJSFrrTz/4LCpnSQbewMFIO8J+LDaUqPOdefT2t1A7e6SH86d1ASdcM
M3hQqZobMbV+vJ2QpeeN1EkEMM3ELlKbGCIxqOV3skakWmcDjNqWSdnhiPPY6CWvbRYw7EavyDCn
SFFR8qSOwD0IsFfj6whxCMj0zrc2Ydnd5rTsbU/5KZYxyiU7dmz1rQCOrvqghFeYrEBCSZ2Bz+Cj
SpnqW6U3x06pi7z9yJ+aHnysJBXwQByJTAkLJhqUKZ6GyR3WnR7GAxrDsl5gYlhroVn0WIVyne4k
tZktOTViFliy3ZnGlP63HWPH8VoKbzTFqKApFHeYJ9NuTYogiyoVEQ55BhYpr0Q1JF4XhXIyl+US
3/Fo9hhs4lKGzhyMbv3j3ZycXtKA8sFK8zEf57eg5OakJz/G5N4bzDTAvofbDHdOfK/JJUDXIdeC
qBBC/cpiqMYkhVm8/qCgyvaZmESmPLJVGCVDqCQPnzbDnag+/jX1FSSeeKhRWiwwiwYOo4UcChin
rWOuOKFKmnsjqPNm1KntiGJ3N5e6I12hPrGW6Wr7+5zne9yA51O3fh6vPNNZCBNx68yZj+SysGJX
7iBRgdHAT9UyWUolzKn0xYCJdR/dXFdiAHQ+DauSIdDQ6cKBORGrt+jC2Sgav8T8p2rUju0sHImn
G7MqWR6KfljvXLnYAKFmwKxqyq3S1iVGMP7dNRGhl061JMkt1MLB+h0lW1yXoreltl2VKO4e3cbh
/nxJj4y64L7KIabqbjPoDIGt3f/UX+Ts7j0uGIrYd0U29RIZ7JmCVukLhFjRpr92tQcoY+QrfDNu
URc34+tPrhqz0J8YSEHtYKS1D45BpifSG1XZmjH4XhbOqPXkMidAYIhskCqGLAx/nWgdXulYGC1O
QlcWVayi1nXFNJ04q+45aikZ61PcOV+QPYWl3OzwIJ15P2lorNa9w6760mLUJxLDnJbpr2bQ717q
ATFs7XPPruOB1ACsidPvRPkC/7lSgmPfYskf6ZzHhf3NkKysIzsYvzJZP/XqjJ1+bdFW4EPHpQR2
5A7pV15UUqJ2mAryfiX9YeExlS9hO+1Z5wOpMpYqGRoUvZtPp3bNu2k2DyUV6T38UoWwH7iB9c7Z
SBoBcL/XpJAnuRKoJQyPKy0ncXpSzAK+hh6NDZ9D3KrWiJt5eOBkJB4kCeTDwQvlIYF0wl+0phWC
WqcGNloNeQqiWEcRPFQG3J9k4Ryxe6W++mTBhQH2fJnJsroPvtdexbYBsM1/d91vVhS3BNTerb0W
uBIzHcuAtIoetd+rZ3a+MDmWAgSNgYmF9spsi1BRRbqCLfOOkF1pg0+dRVrF5jzkR2TmkivEhuzF
gGJSipfOfOn4U8NfEV3cqQ2qemZdt5IiRUG7aPzA6hpd327i8V/5guOufI1Qw2nki0nkOODl3HQH
HqUtFEX2umsRnoM8w/dn0sK00gEqdZqPiWukrS3aiFHJDdxdvdZxpauZVR23L1TrHOsl+ThWyWxe
8h86MWGci+rg9oiWomSljbPapIsbYfk5hTA3kD56LSM6OBp6FcBC2dinff8ohQl0IMks1gFE0eKF
2sKb0I7biPShTCZNTcS8+gh54FgNP6O8xzcLNw4eNkO4YnA/qfeYuQzAQFWw2x3wOB65jwTpH2sO
A1d4MmaIkHWoZWsr9prEdTRcgoI87lJBEhXtVJNNyMkZq6rExgihTEkjL9FE2+lkheY2WJfE8D+G
lH0+HMYYVOAfYzb6C2HN6dosU1Z51Z9b/qeSbCJJ94GeKQU778RwkjgQnm1+OKNmZ5slnsfovIsy
8cSEh3Gg1fu4KIpVJFIXOn0wSGeprCfLljbEUmX7i2h4QW0vUg/uggGadEy0rN3/HWBZhGo0JelO
2CdqqQhO5l+s9WYyc9d8yVGIZOsBD80WmPs3Hbvqb9pWok3/YKHX5WPrYkdcmCwvjJ9N6RhYUgEp
EiNnzUCPDc5c9Jzjwuj0XAtsEe8j+i/BzNAoENk5Kmd6MgGmzHeS334sHxHYIIKWizgnASiAOk1c
mkXDFDrE5HLjLGtdih4/L0QeKwo38/ZDlomYMqyJiAEw2wKpykKHVxE+A3+1rD9Ev2vUJ/Y7T/Kl
2ZTafALwYsgGWlBFVYmv+U3t//RbdYmIv9Mhvi2tfNnXygv+oqe9COZuywFShqUcN5suPQxYz6nM
E4EnU6frP/r9hRDOIl41RZCQ111+YRxjb8l42ormKciZpA6q+YOStmCQLlFec9hhjAxke8+OpzmN
OXtRAoZHQBvoi0HfhG49alJDihqzW8aBPlBFbFpdjozyxzAagBpiinH/KkAbiT8q0rkPrY6t2F1X
I/oVLeJy1KHji7RxH2lvY7StCjK40eir4HCSaKNpUd4+JKu1/amVFq4VEa/1sLCIZcJ+uKffG+r2
HbH1n3fLJA4/3qK7t+Co+BnEItTzziKg0G7rbDvLPw68lPem/+BorUWUOSv457RpN2OnvznH0rUi
GaTqMtlTeADTsp79WMkYFl27hMQ2TvGlUCUJADmc0oLRS2b90fyCFOkDgEUXxGwWS1j8k1MCqtCy
SuRES6mqICc7y4wVDouaEENwxyr4YH7oJeS0o+QMnbbVBoa19+W6Hc0q4VM1h77UNtsXLtzu9bqH
yKTMt/R5ezbiQGH+5lJxWNMQElPLL87llmm2UG0PYalXsmnqczp1ANKbmaLj9al8W5eMuSH1zbwm
MEv3L6qkNgso63nF3WCDlM1jEP2IGJOaU+aMa1rPC0dGWz4OMg6JvmPJQy/SFwOVhR51lRjgOKge
oLT5RO/FMW4jqP9VCh4pzRJLwUJTPl7OsHQ6w6Vys9gYAHTa3xj7oLLIuhPm57KzhqiHs86+1LGZ
OQR6oGSYO95wloxiUFTEwloGmQNA7iiBslu4/AAD7cvjvKzrh2xqViMtepI1Thmmot6OhjIjX7Ph
5gDZCLZYxUjj7R34pC86bm8V0U51QKlQ19y7W0TzE4G6ZLtNdAs7d/moIuG52ywjz13mfafLg7LC
BuLaW+n1ENIH/8i7aq6Gz8YmptfrHa+2xIBZlcwUHr04P7if5mQ7xV3gzqfzJqAtigsFW57+Y1Mc
SW3Hkkn6jhoSFsuN/bVYLrtKYgWhYRlduIJJ5TQT4ZdMmxrfzaoe2Y84CYZUdwzmAi2DDcOxpxBF
+w8ZMfiQfeY/A1qT3uDD9YZzsKVx9GG/q4Yoa4U3ai951fC87sOqkKAzhdiMnjQfcexh8nbCf41O
XaxWf6vauinfVXRPHzXuSNyHAI69dbCaRtBY4vp+VTczP7ISFuhRQG38+2NI9F3BJ3MafS3Rxh/p
yoPtZlHK0CXWoVkNrCCnNprG7p+ZjrrlJeMHNQlLfUKRCJ/OgRm0BN1JP5xMnxlNxPHNckz76stj
Iw5/W8JhNS21XlPgwyvXBS5WBzl08nF/G0IYYFmTcYUg8zLrerbf67NkNKfaQnI0BLeDAVuPqb5q
Usg+7r+/m8+4jykg9xeCAxJ4n2/vIRfg6i7t1OEdUbWkmOdlPfged6lvRnyOw7XuWT2Dex4FIDpN
GuB5SvJxViGYNOZy1JKmApCddYz8YqhrkNdoj6vvW/hLCFkwdcq2Ch1j96DG2iKfoAJs++3DbfMW
x1jpUiOWFQu6D9CCoP83MBK70/FlEe2oYCkI3nDQEFBYZ8pz5g4bV3QpnE5FBZEp5dC/23uGJC2l
Q93JpZVAazNsePh9+XA5zLQwxp16wXqFqK1ZGAKgSJFda8DAtvATrdxRBQAPGoXcLcr3qQWeIyph
SaOc/NFXlQTbuj4WT5/dEZ0B5nlNdhFbaq1Sm5wX1DxIp2vsdwplHDpilk+XFabO6/OCgxOAa7+q
Kq9erHXf1G+ooO0Sgn0JeYCvmbhcpRRXuyFOAdvw14kRJDUa6MotoxGIENaHTNGAa1GaJ/YIGj89
OqFMX9UUbfRfqkIPQJ09lRKvWlymrSBySFqqbE/T8tWBuy6MQtJ1OooUZe/ScLosXndvYPfwW2Nd
IEfPf5k9N85QkUjZtt3qGVkiwS+pxt6W1c3kIuCLahyr+7I17UNXCKywTk7pYE9qds/u7PLaGece
keE+Pb10V0zUt00MGudgOklcAtHLiQU2U+y3ZR4mCXnZdcPwJ+J4lo0LYvOQCwabOqj9sMMEUUNr
ErdoSGGMKS1wr9cUUpb/ac1Jr+QQnbJBaiaaChfhC+C1tMSi2wl/7tpiAB5HFILeotis+4Unampm
JJrSZMD+sBPNCeadsIH2wcRkqSjQyJ3LV5vxuBs4dsV9cYEb+ZMCE441sz0AdTseg5e1UXdQEizO
GP/h2xhJ84ZZC2eG3HMp9DERmluNilf9WlToJY6I0ZbrEHYDek9ylhFC2Et8YNlzHGTbdE89OkVp
axselTiRxZEAFD3lHaEOCjxQda1kcDi6Y6EzGF8raYpBTTAeGNk13DwmxmFVc03QEw7JCLK3AXy2
OTBmx+gvSBF0/SFRsBOn8E36wvtwAw7RESinQMAtwLIYLsYdZeSzCRY7d2Bm45m17kMTvnYwGDqE
LglWFx7vW/Cp0OMvAdSoY14PBnpfgk+2BZ52T2kl6mP8Rdpuu7iNumwLxyFdJMpgBLJ+6TgOBanm
1KLqOWdV2PEoaWgngtBpX6SlaOjCPNrJ1iUpSDGnSBoILTL5Uua6mxcgQX/dqtxDZJ7kb0Y3Bv31
camlNENoTn89dn3XjPBTF7fdVrkWZRfwPSd+L0JJvyns2AZvXVy/233Ry28T4Kig+5Q0JEkJE5JX
n/gLAwhwJnoZYszmYYTTfjfDHYZeNdyHOBHvegDlHuBHY9+SSk+DgVpHlPHuAYUI0qPqCuAxG5Hc
A1CNwFfS6hFyjFNmwrJglMsX9TE8ib0KhjBFUfNe8f95L7B+o0g6e8fneeYX5YJFoqgY1tClXjOP
L2jYOIuEHLabaHoC+s8bI3FjMC8zJbHZmYkEBv5TTnc6JO6sneld61eqT4U6JRyj2CTG4waYxUFv
AtBHiGHhPDs3CYAcQiA/3n7R591+a7tRcJ3i3GxjDo0z0TUxPiIe/u3vY0Zr4Nik9u05X9B050+4
TG0xFirJGz6URtU3s0cNAqXWYVttxAgSJ97KM0EUpRNDxnMysDh0pKoDgdAJDjFzwPr7AMzCy1wk
cM81+0DX+8xGvQst/JXcH/x8F6DofWq12iwFFGI0DAWmfN+4pOtOHxhYH4j2f9p0ycz7V1AiZcRX
L5VA2n4aB40LSvz5SbLVdaEkOs04sNPf1y/jCNM7y3IFccjCZR2f2bJ/BM+mkM3HwgJ+sx5ODpbI
SeXZPFHl9Tg355QFE6I5tEFHw7blsjm3X6SfvHvjYzxPzrLIRdPidEH0hSY2TYCu4ZWEwHvoG/FU
NTNWBllB/QGU8AHfeoOZ7xLXbNPE6w+4rH4Kxm1thquZ3LtzAwthEQKpkEADSTUnNBY7ocZON1Wd
KKb1bN+nGllF1WHB+Xo1gd4eUg8fN2aihI+xbr1Q2qp7/zmS8Xv0t6NmEQ/vSY9W6PxFJlH7C44q
wZR69iVRqnILqQKqKF1jtMYurOXn7H9odNXMZG1+hWUsG9aMeh+ZQYUFyuGYKoCjL+u0pfs8Zn51
sqvGZSRm/Vmx8gVAAJoVkq7uXX5NJe9mR3sOV6T613ZtLdXvHnkOA7e5r2MD+b0v6gvF/vEMyrbq
izUU0z484i4jGsN1pWksuQBdrmNsINJ8rt5FQCVGaULH4NGr+a1dZjSjgXvNgRV/n08b9OIIz921
zgJPQmnY2RyeDD5Gl4bs2iBzOja6OlVLNRGQejb6mP7BQgbNSj8b4zQxAVsBcwGtUtTuv7gD/EoB
2EwESwuBWzcanxfBu0LqlHsxHWU9kH4KMJKQHbniCaRh6wWNwOv6HgIQhrkHdqHCJN7kUJIMd9eq
YcPD9Z/4IIEqC3tPMEjBZsjmMiEmunfeALGK3QZKX4KtDDv28jNqqUcPmyLLLWvoaBhDQvI70LV3
yLVlP1xMKup7ecGV/VuVLl6kHUNTt21pndBRTm9uc2WBn7Yt4cMUIQcG1aZk2ktfM+tt1hbB66kD
vh2sQt7joIvb3Ux3EBq088/YOJpKHq7YLywLW5ZlTFdpkgPgWPCCcaprqRlb+9YpOXwY6YNOR+XG
aIaJJqMbUSWU69mfn9qxyPPJkaxdtPPGKu/IsRpRQcLiwczeza55CqpD43xP78InyYM4XhLEUfVU
oyGOdg8UQ/dC/2lnG+JOvM9MNOIQ4A8gTSLpasQYeAczzEV0M7djU/+7fUsAcIyw3KPpBDMG5b/E
J558+k4bn/hUwTFTqKaADNBEEXIdd7aoyCCr77RdFfYhjdsIaH+zF4aHnldhCI0SgQ9uGjYf0Hid
72smmF57XVQyhY0o7M4CS0U8z65T2QhE50XGCA+Ud3klkNyNz+CdUz2QfLx7RsPx04Xy26V2WFaj
6rZ9BvxSE4baxqQ3fZcGZp5sKuHr5YFqgeIjR2yV3ZO8QF+8MCODcBVQ4ZitKC0gD4nyc3o7sjIt
NnLUQYcxOvvN1Zf1cZANLnFoJ73fFeX3iqbM5eYD9E9mdnBRXouGuPnX+rhFJOM6KNlHgFUKUNAY
ja5dvHM7iwKVF5sLjJSXWz1b+taYIyxJtd0N1v3LvbyQMglRYbGDOhev2+NdyhXkSC6WOxmO3zTx
5RjqwYx4V4Xsjye609h2GWtpDnqVQl/7eta/r4xV523d4g7VrtXcedQs02/3WTAvT2jvzhQ6s+YJ
CCJ+PsQlQ0SE2Oek0I/fq9Bkwz/xbQUhFwWPos07/1OWZXqJDVLOwrKArIrtQOHgbky3516RHI4y
wUHZkXjnw/pgTT3Lc2Omt+b3sIeTf84T+XnFKifN6DHYES1YY4klj8usSBbD2iMIYnpfumAe9pHZ
Fa1VHuxvaSAV92Igov9AgCDIM8TtScqVcMIpmjE97hmiuiEUlzW3hyhSmzK9r1G7a7nMHXpxVj5I
u0ygS/SzToqL+xJVE2ImQj8KApnDPM+MkoKde9ObZ6miRkn619dzLFl0K66KEeyoTf4l1z74vZ/M
u3ooKqNWx3V3fanuHPcmCfyxrWemZkkIkARZZjlgf5y2pqK62Vk96mA3S57I4XVv1K0vk2X6R6Us
eAEWU3ywUJnKld8nfiLvw7qwmj+HzWH+iAV3s3j2AZSlDqAL2iHkPbP7NGjgdVOvHQs9HN0zq6nM
JP4j51AmMQ2JXfYE4oKAxXYAuuOLDL9viQ7RLkqlGJAPY1Xv7quCN2zFJuJtYJhkfJqrZ3UoiorK
UBXRsXEvR/DWQqJS8GQcrH4XQZFEvcambg0bIDhPpmNm15poJWzvwS7TnqAG0LRhHqHB303B8xK8
47iApYGd0L71vIoNiDFNfdKEDWd6M0ThlFvcJxDWHP6QikLUO85DBTT4O9rU3NShbhuOtMyOK5xH
OcmlsIbMkL1T4kRaMEZ4SpBSnEycFrKQt7KoU/S2n71k2QXX9oF4zRzyQvtpma9jrRth3lnYDSlU
dbFtHor84vaJ2uLPXRo6C98v8KY/FYuKFbolk6P9RqvEUeOiBAii03kCVRwUZ/Frej+tnnU059zJ
vcuH3/inearvsAFtsSBkLymAiMpayq4yOgO/psbC4plkyyAnbuCKVzOQ1kpnzhCvYO4U33exPePe
xkLCuJq4xziCPTg2EJLkxds5sl2zNb/xf1Vfug/hTX3aRBhghe8Z+pERoaHWJ3j6Dtupcj72+DDY
FPegQPQTo3WHiE0Ddk5hrPzfbSCoAiVX1Dw4foS2wveHREcPlPqnfPs42Qq/WFoJ04ZAlA+vSAKQ
35zD9F716KYWw2X5R+R9Y0sP8cHN26F2ESmm3q81wyJuotVwtNSsMtJZ+jOTIMaB6oT9YPvXz0/u
Fq9xoEXqtTO7U9I0bX6r9o9anWWk3zkicXX/4V+QVUQrujsFHqInmT82FE7cyj84Eb0Z2rIYWhoW
I4GqNeKEQyV6f1aNbxCaZcDL0vd4b4qA85ZyPZSSJFjCVD9bLOobk3lL2qcQBZr/xRlx7a6KIbZG
EjD8IQpd8noe4MxnqFZz4lwT7ZizWrjxSrAh5vPPNwHrQ7SHxuVfm4EkIc8t0H3iEQe/usVmbxxv
rcWD1aUzKbroJGsblxxwuub04/IfIKZpM7XYrkxB2SLCx9aknRaTimnEoLXVssJcRqQG2Ce/C/2t
K9LrwQig9xOzmcEWkgNW2tzu6eYCZhoN9hOrDPcgEU30fZzX5euAP5JzTcgi4VoLC1OAdcVee6OG
X5MPO+K/EevxfBjkne95CyMZmY4tXkdMMg9/dbG4IlNiEjp4JNRnQB/VJVEc6xH0t/Zu+IhFDQHn
ZIyE4lFQQGdp+3llsMTCI4TJIn7QXFnwEsLHtNHL7QLGIKFkYFyPZ+cbZJ0kavT+gLX+5MmQbMBF
RXDaS2A5cspGIsUZTGJuq8QhW3bacO0/hU5tRRTB4q5JpQEPHqxVQiA/hlV8H9NuSvsXeelGZ+o3
2pxoJkx/GTIRBSz2hfmAqk4ZY/knvC4DEpK0oI0eg7+w91qG+XkI2YfeD1zUvnDatOhhOBncJypJ
mek2Ko3A3v+KInFiGv6jhhOyX7FKSt6CJejZYIXmNQ8XLPKZ4qU0RBsbQ9JU8ays1Hp94D5T3qxZ
pOveEpelqd5V309VtGyS0GBDhRPDNxREt5t/uXyn1yOFqSpqC4GJSchghQ8TaglkcaO2bJnFvypL
2DTG/UCx5FULmOrJho3Do53YMRlPNV6iGK56SRUYRTxWj9lz18yt/NIB6sm6ZVH7J0W8n8Gnn1NM
yMRQVHRoA/xL6FvXmHxzL4EFBLL2ICOlZVnDknpwsQjr5RQG8L6z+ayQEdhrA+ctXrlK8R6B6Bnz
X6BbxXu5ivRTmPcbOtj+qHvjjGPLhAzRmO0VKERqensLy8YWkLLbnmA06DRnWShbnxbtq3VDJy9Q
yW6HEZ3sLxhaKV9zSERxCUKuKaN0x00yQ8LFYn7NO1QiuYY+k79oyO93TB4vmec8cvivcCtmt922
bLPvTmI88Gth+YIKAzr4gNv//A0DlA7nNakaVzq8Roqr8NvXwBnjMwRdtBQ4Tmgwk8RGMSmkKNpC
oo0QKRrR239STXdTDoOGDE8MN2PTm4nzMKxUEr+xwhxzYfHU2+EZ/m+6cp1HDpOpiomgBqH4/Z5z
KYEeQxmX+ZrnDT45Vw4Z6WHjmm+VODzUJz0Ia8w4TCe6qpVMUEuJeYEeC7TE+zi52uwQncuk5zqK
VdWz4tAeAZRsLFMV/TWdPb6zE68G7PyqF4rMnlxGBBvgk69ZXGvMM4uye16/0nYoebtTyWkyQmBD
/ocEl068VJPUUhopwbxjw88x1WIhvKwIM3UTiN9rsN+iz4nI39cRZJioH7WOiQPRrnlmzhOPOLPf
ohbHo+vUOKjlezfEIUv1l22fApifkrrD1yjLvU4uKGtCkhYabTIGOpSVULIK5a+fnWF7W+V0q4Ys
HsdrQi/UKKR6SlN3myLN83knLpqRtVgDG2SWcZq2LUQGoF6i1HH1B2vJHK/lgj6e323k7hJ16Y5H
y0ztyTKnLfW9bVZ0aY5KQ4rwYUO0k7h/OHRz2jeYbofTmd43VVMZ1vyGpvg7TkGP/574XJkfNbd3
Sty0aAxVlLlZQGORZ3gDqgM0hy1e1X8bWeLWKs+32/jnSK45kKGXyTx3U9cMyLYrO4niXjNfK7OE
l+froLXh82jCsDUcNGCbpatGJtY7UnfzAPVl/EO3LAlcnkOKXLX20L8EXbiWk1tkf4idnm1Ds0cm
qNcW0J5uDGxGm3xZBfSXEG8QhqoWv+joKSsp1N/e3oTcpcLOp2sOVzz56tnQ5Hqnoxj+331iUzi/
gwHuVPMOmDl6qelXpWFtKMX5Kz6kY0A5NTLyIJGBnIqFL19bloy7ViIAPTTHbHVVNawFGiDX+XR9
2VOPjfcmIutVt45n5lc5jzawwKJ9rUF4edNK7/q6VhyNXGeJep0ug6hP7HFNW6Oiy1j8b9AuMbCI
mu8Wn9REzdpma5JM0zZbxEx5WdtnDkjwtOPvpbO7KxccjF3eMXSicZ/R1ZMWIqtNskwMdlZBtBtP
D7gwAi6UT7/e+lpDREgxyUo4MfcsKNjP8l0kOtkqt0aWe61ubdb2gXzI/2p//ElAl2fQDBqvIlYM
HGG5Czcmw1RONkz498UO+AhhJSGkNzwMUGAhilByU5geZ8QdZp1fmaMBK0tjEwU4lQat6BiZZ0y1
/PcScUgHJjSCf+aobEY0HNFrsdN8ahe5mxw2B8XsH5hn8KzVs8Xvwd6cFUpZd0s93qo/08xZ18WT
jmcoSapxgIErmSP2qtXhcV302CBp+mA5gGUIqDEue/8tFpGWj5ibg2PyZLym7L+2y0kvJIJP8m9z
drV6eraPUnA1uqeJSBh98RYScX7PyQSfA0Ruo32RmlExY25MB7TpLNFjJX1Hh2KlHfDEtejVVKtw
1ClvvGzqFYOgtHPFxCVfP7HW22MPq3rdJOez+McOiNLUDWmX79bRjtmOdjf26MBQHU+DqtRwVVvG
1rALoq+eyjUJgGTbLq097df8Gz4JWsNw1fjZS7TWP2WyHbHS0tHFKCM409gRspVCQqfp0BO48kj6
qCDbmpVtC5OVf+M/EudELVvApHEU12PeE1CuTIcbpXiY5Je1pTLoX19/YWmCIgcNxGOpSWK3zJnm
4heLSrm7eE/OM7v1nJcVf6BQ38e5pFV5V1sNM3MorEuwxKvVP/pC+lVs451TMvDvPf1SYxAdQqg1
KRBlMJDJS4J7zu3FpXxjJBXOdJt0VfjIfXNg8JhMZNGCRe1J9hUoyHT6h5Ur433f0/KAuThDfCSL
NG6+gBXRvVWlMUXe0xU0iBXx1V5rEkcu8EtaHRfGwI3jMk73XAb/55mer07j+GkZ/5ctKQfiaRri
EwoHD12Fc0/w9HbT7DVv1P5c7yFg4AINVhMdSoz0qtLzzxxoaxD7YIjqPmX9wBqvo3tgHgZgTkEi
Y61lFCYIogLQ3yVRTpWL/jL2a2dAG4qPIkgztY6AF86oWbXGjVxe7RoSUx5qxB8kF/5ViBypWqfn
H4GGIpVvGCVpYkKdUSKMT5/8Vvea5qJTtKxN3hAPaI5cvOLBL3gTRJt/1KB82oumwgN4frx3ibjF
DNiTlO5UidCCym6Dq8HgbtoSpDgCVQKqkxE1p9k3cijedYA44g1gSgTgtKO4ZzcO+7LY9qvYoQTy
cVzULjO/GmRTueHFTvAd2Ks6d7GfBJVMZCabtlqDRCGk0Nfnrbe3JnmJ6RrEVLXbE2N1fa5Z480P
NTiRWL3d8E24kM7GIP4DbMNgOcZiUGoehjxRf13oWNu1N7x1euaS38x5Hu1WEEbFdhAn+ZReOisX
Tv68HAL1uLagVHbIgJTiKOTxuR/w7rMmQVc/Ji+DHa2L/qwhs1U3ZLOJs5TeQeSCMhDo1X4HVMrs
iGJTrkHhkt+CgX4thUaozYfMR7SbicIp4K6Gwp2Lbc1ZN4WiZ+SRLMyddvNs8aipFS6OE8xbDorP
cZn1DjtHqC0OG1J+T0VAn383cFuYNv1CM0VKcJ/Xhvka58Ki9ajND6q6X5AAsJS+EEE3A4BA9w4b
1KwA28z3iizwSvOhDTR/y4iE3l5eKpqluleb/zLVHE2C/GuPiX9QzQ6+KpIkBxzEd/zTwGFWUIUj
CQny5GmAIEhN7b4IOtDICFHtlsFNdJLa5+EbHEIrklc2ERv/JJhCz+Y/T100OZRtjFKh1U2f2eF7
gwc5p9FXa74QAhtivBWC0+O/9WL5GpWN5SPH7mhg3dGkbllfhL2sVtQLacaNeXNsapkGSNOCiKQB
c7u4TplFUUPim+RFAnQmUnXLE24Mune2EP1jXBklaEIvxbgnR0wQWpTbLYSSGCiZBTt19vJxRoBu
Tip+IHGielUfLZK/YiqJo2pSPT3RExKuEbxeTOFmHhUwZ0HeJgGVH0y+L+YWK9jaaDTNLO7inB55
SnAi0e3YL4q0WTJDvGU4ILaB4RnkqUQsibVYvwGJVuVd1LSIAFD3vc+jkqSNuWY+X+aoWYDpxjfI
z7MNONsgQpqrmEm2O5rpCc1mPPxo1/qqEdDkOL4/4L4TzG1Zw0vPoVhNoQMNv0PCXRyNUMLLIxpG
9jOzfp/14hoIrvzoRt3CPs2C5TR5ymkcZfebVQUnsRNzo5WjgrutLFzIFoxXnNUFWM56fAaI+87G
WQ7ScP8scBK1R63i3V28ElW3TRLaDrSwKWnExRv3bw3ysmoOlnsipBiZRUtzGtSYbZHMMBrIRYwy
9E0/LcVLUfqleNiXDDd9nMxwakze47P0dleVc40vReWIYduYPficUHGX57Sx4l7UFjRSxiorLFkW
IUmOiAg/YAkRz3CexPM7X0GcJiPZ8gdPIkmL4d0XhR7gN2JuHFHMfc2BpVpq9lprE/BUy4eUspuy
jzmaxSJ38aLm8woxvH0GyCdXzBeeKgpYvN1Mzt0OPmqhfYzJYLlnxFXkL7iSUH6m0KQvoDCRsUfu
ARaBcWoGqQ4ykHmwyCSc7qlRL0uytJVQWO8nI0mre4R4cN4sx3tCaC2FWINdOUnzm/Lp8eQfzO1T
PBVnmPVAlcpCSKnJtvktvbgflzgvq3tpRToGMDaWpaqpXAY0RQuBVIxelJOqUyu978/zTRYgbnGr
m+TwX741O5jYPjGMQPeB/cEFi6xDbvLbJYbp6dnrJCWipqfFMZnJWpxUIxPM3URhabCygCtMR/04
qzoWCQ9+MXUAtQ0uoMpZCHicC8cET5ml1/rgdcAFUo8+oOlGtbK1o8WBfvEaGHGWxoEWDU9XCmaT
Ns2YP/bqn12mo7taWeRJFSNq+i++GJC2mcReGfiqSUoRbkaSkHIzReAO8tFWsTYhuUVY15J+nAel
hoUfTBnrHIoREyKlnA61VtkziUSc/73zUnxeuocaqtZCtpuU2vnz5iu4FV9aZuSxDSdiFKqzxeSl
7Y6+auhfI9R/X0nfEZNoe2YLAKS9v2U1Z24n0R4cplLgHm63vsVpBDbDHQsGxs4qXTFaVxFqR+MV
RyUxrews5KJgliejmnTVhd6dM5t+UdLLyq1ThMxYLRh98Akypj7SG9mmFWMZPx2eYS3d8s++Id1k
1i5IXYnDVCLQ9dbSu4GnuUFgFoiqx/YwOv+T5rpWicB+wTcD2AL93vxw2jBvsJOHtVwlLX5s75e7
ciQtnmgPtR88hT1NGh2omUD7OhodzNdKtQI40G8Zf4Sgg8HjyNmMtSpSX4n+mu9tFVSDXmWMmhLQ
/5ZpdH6v3XhZw7WJi9P9c8W75o4DfOuolUqp10W6lj+NmQG8zm3Iz2ahdmoleSV00h1Up5O5Rdib
gGLMperxQGYOER+h0rZ8bxk3u3RMtm6RkyKa3kvmK8rSCB92u0+rVSlhk8sMeYWlx8uZ26eE1b+S
2gD5qlyQWxxeKBNx5gplhl9GdXfwDT3UCx0aMN1FdvDKYVX1YGv827WR34ULoqDzAt0NZWAjuVb6
ObVwGiKoc96v23ki73j/hGQpDpOi3PrROJi+6b8nY41xFH8f9PlOm+DlB7RiuVfWTfJtesp/9pJu
4aTrG5PRHDMHN8cefAFxTVkoy7cuIs/v2PGaCUllFBnWYDNWI9ChOi8ABKLuOLzC3rKMzLTItyUT
X/U25zOdcpEqi222pwBldzQ4jnHg/5qA2Gc4HBorP8Td0F49INHDIir3BA6HD+l+s4ZT7PLtPkFM
jvHfLshEZmv6ylY7fkMKL+/+wqJaPzcvyBjysnZW24kd3TwW0mfbiLFJN231CqDzFap0+xjCt12K
tVldnGXX/MrG/hsv1HV0wQGWQBT2RZSKtrXSllONM0MWweb2BpDUsr0g4JqtizaFc9SzL0EjSy4s
2gdjl4UpydOJ7gMdWBm8ib29V1tBuZQSSmxRlusNk7M7ubSsEY9hQrqWKDScaihmc8PolXL8oWhN
mS9JKwZMQffGNjDwvw6H4AnOAmAnHTvDqTgGum2BSfL7qEVbpafC81wf4fpTelR1VF0EurR8UpmF
Bk9BqRngmckMdeSnYdP0ST9nAutFIvgSMVEKzXXGg3OpjZBNHphkdhgqo2snsl3vwZaUrgDcOLEa
N4p0y82DDDfOHn8i3jjKeFxcH6rrN/odU+L+uPzVD5FifWOXZrVQ4q9PlOu1uymzKFU+gNoDGHkn
rUbQGSGsI11wQlOKeQdoX0Z3F5uMzCJySQcJ9gBFTyKzLG2AARuq4Mr1G+w3syVmOZz5VtflTijK
ONfpO5wEfvfkF7G5+xJn9jCDfT05jCRhTP22IrJi24f+TzQkfdlIbBM86SgDQADuaoch6AJrDCHV
/hpZdNcB5Ezq7CPyATU3EtueqCBCiQLBTGuADzrmOxKkvdyuSiGhGxwBHd6PNZ7wopD76Znh03qR
OEbTutHMSBkdPBta+HNwSg6IQXJH4ao7UMbz8+iShgBlCuRR9gZ0KfMcPOIawCdJh27qYaZR9VOZ
YgkWvr0rmJqS6MzQccYklAlAJmb8dEazCzj2y/duhffeBTmEi8HKr3DmgRw36l7Eh2YCoNMCEDoV
5JlEA3CKOnOit6YTx6lEAh3xQo4LJIykolQfWJhm42XUk7+AdlfX+xmyZ/vlmwLnZ58NI5foNYao
AhEDSOC3f8cScK8AqaIuk78kXThp1TwiYxt074g7D5qocksj0Af4xG8Lg0mrViwKYHIRGZntZXbK
yPeDFBNVCXcbIkJOr9eXLdtT+kYDchJTJNkGAG+6lVjQ1/7PFC9qvMYA60snq8gh4aboA1A8eaVJ
EL6QhNlFtAO/TLvgPBBoyILqQEpY8pxuZkigfE3ev3lpDiZd6U9sd/WYi80e0EvEEnOnCpmPXU8q
EFVGPQoXz7p4aGbeN5xswCfpS9V3JnvahHMyvSEK360pSRCNCfzv/PNak0a1QDRIOnk6rvyuRS6T
FlTHK6uc2x8RgCD19UaEdqj3uUlydKNWelWQngYh9yfub9HYtqkvDcbtRKjVpYKo4XKI9UUvME1R
SstCPNfBWe+LcnEGaqeaZ9KQkSJ0oXUezCC53vzsCaqNRXbtzXdGgoRCVkGnA645rCalZF6canWa
n6ta38yV2lLbXZ1RVQmei18lnPFPi6A/dVxJrTMR7w8mxVePFR+WLzwLuRjzdsfY3Q8RJZnmb4jP
JOG3ydmXE5Zg2UGdEnqWFMfa+gVY0dFpA1D7giJsYJ7hq6gw+4lYj0XKq+s05L7tP6iA3PHv3JVU
jMOQmkgDBiNZ+Bpfh38qeDZ/Jcgcw2M4BIEQoAEseYSKi7SfWnvJUBB7dBFNtnDu+SfejPyTLizt
Fn5q5XhpQZqQsViGYEpbfa53OBJNHljOjK8jDDaFhZgnoRCt2eQmA4x+2Mn8zY8b1wbsV6EQ1feQ
DELGIwZftJW20MtUeB4mUqDD6xEAG0uRWo3HT9knqHRGjvNVLm4yO6G9J0t0FywJPVXQCx5/puMF
ANGJ26wIadr9DQ7OS8fnwD6fTcTdeF0Joh9OZLzUkIkIDqn43NJn2T2Z+hOTdpCA/Hti9jFpWJx6
2XLziPe3jPlae6ObiYJhCNUHyAuRvg16pkCz3+m4+g/BmHVaPMfGVQb8X9XPNjZqMKLpm9h8ffRS
vtmLxFdDgPCEUTqci03EttZ2NwVsxHF48hnTw35HSHT42os5d9qJ2A7f+i//tgNL2mRhXJqOuQ/o
0dOo3jFRv1IOYRc07Qec3adlmM0r3mtFKaeb4vTv7M9RJSo3VafrzHX90OuI3CWXFq/Q4DIZfLoy
OYut6vNp2BJHVm7djKY4oarjylGAF/sKVlXzPBbMJFaB0VCuLWjBv3n2W+0wIUO2xNVscsSvxCtt
kp6ZBHSBAGoBfFmhxeuNpo7LhVXG43o+N/fGADVa51HoA0wp0YWofcKfsd0BN+rH+yq+PmcOL7YV
9PoTuy109kKOVKzMXqfVucekx0W2JQEahL32LnAg7B/KPeZCqjP34mq7Gshq3yEgswSEdCvugwMu
oDIvuSmcbUnqb4pdo985A1yf5pxGJYFMnuTwKCI7FGWjsskf4LDKEWzPA21y0D00Fqt7hLPUEIET
JtJl6Y2I+QceZikdHyX1uJywhr15hWtm+Bp1jScc7TAYHP8MqjSZhEXXaGVx3RvZBZwAVSTYvQ4W
8kNYSZkjg67/KexaEa0va55UMtyBiyVz5v5xGj9tggEhhd0SE8fGrzkqvr/+qPFZAWVAukeHd/HS
TIwwQRU+lg0717rGo/KMOapN2SyZmms1Y+mcKPdOCbu+YLfvqTvwNF3hzrRo3lvN+DCeJF7QvkaF
Ar9I9CQC6lmgt288jAS2f/9iB2J1DlzFSqDWqnRw7KyWZzG4QFf3fmxy9bIJXcXqQ/fMeyBNJMUC
Q0YVdxhN4J7TF/0rdZ5JKo571qhHWwGxYuiSn5a7iPHz0ciSghahUsDX8j2zeOW6fzpm0UV8Idfr
Ar4M5fgEJmofW4WaW4YveDK4k2up4rreOiy4zZnx4WHjqk6+NI2EvJWbFa9tSh1W1PEUjjdb2rfm
mYqUxlVLml7WGwng+oZKhlubHRKrabsKC07tSCzSM24+nO+dbg3DUlTe3IIhsi8JgkdshKJXiJ4N
YVxyKqzYJOa9X4XapNh9/0I16rzfbVsR/fhVyYS1MKk5eW9q7R3QnNGwWXnE9z6ZnT+69hc/4Aau
qoCW32PKKyJ3L9FczgR9steye6JL9F/Qq4Wf9PL9xy5Nmnd9TelSatVpB6J57ynq18nvitLH0PEM
blIYKl6AHWBW04bExRhg4EvMwFASa7JTyU5fxlLVT+EeZtp3rBeWU5e3pOhiJQbox34C6yl/HJi6
Z14/dERXMLqoA4mBM36koFY7CCETdb41gjSjkzpiBkcCAakY5O7q/sz4JH00dOPckxXyZs8jZqaX
m+xe/feYmt+mn/OKjMn8b0FBS4AiTG6PbyilxQGCgBTy979+1wxRSfI5/J/6+vj060gb7HduYQUO
2D+zo/IhGjp8NBwalJ+GHx9Ipk3IOCZuXon8XLXp5F+3m7E+xx8AnpRInYLee4RbTjW3HvgEGAAw
yZ/n9TU6ZEhSSEi3zrWfWAfaPeLiELKEK/r82s3lIfwiR2KH2rindkWp3sT6/hBrpnnamjGUx65w
gF6Qtpiai5UdLI7ZUIXmVF0ECnszKu59yDs5cr2viXVWkkxLAYDlOjUeTwDG8LZ2b8Z49bVFOFM/
fnncE0A6/bfXu0Mcu2U1q/dL1dAG/2QNjiqW78dy0FjzPeS6P6MoLSNLKuGkhsIeB6e9FDqey+iD
p2ixrAzph0/kt/nBZtLjRmmU9sy+Hh2Ge4BgCJnxEK7m2a580qwJAlE8sB0AARXL9kwMGrh5h6LJ
2CLGYp3aXr4fJ7zPWDD8MBYJbIITh6/JnxGiqnQPH8UlUU85ObEF4KetNGleHgGGIgy1ut7Kfuyg
PIKFCaVouEoMi1+Qo+Ei4A2pvghFoq173esFfTcslLa4syK0MKqDTNWtzHwz4etdcHKodn05R8Po
vTHemBHC/wocLb6v0q7Fsvy6qFdL3ulJcAfyY7gbYZUe6OzZsZXD0p+i868+IIZ36y+8SeGHkWK3
RzAB1Sw78tkZgg/Lph0jH3KwELv/l/XPf5wwxPSLLvj/vCfKM+uAPXY6lufduneRLH05Do/KjwFy
OkN9X5O84Zm8EzUS6AlMWWrGS5iVsq4RZEg9JSq1gIzTF5jP2MnnUMLv/kvBlalu9yStiwC/qiII
IYZ6SphFa7fA6D8yRcnt9BCua/YexGwpofyDB/hqlNv+GJc+wt9ByOGr1po790KTQuGfRBNDaBRU
e4YggIr2PHdr3/gyFHTbEtprXZNIbgwGPkEdoUMXgc3ju5ehN8bJSBX8K5xdH5r4BXoxIPnBs7rH
bSw/mACh9hBc/+GIPw0MgNzdwzZbTQS7YJyjBG1kSlT08XBYwI+T18ZerNRSFo8HQCUBBb4Svsrg
T02L/i10lkxUgNP5Jm/CTp4/9JAKmNmNMxUAB8ls2pG5vyL/JrWTy91g0Cw3J+TvJNbPAUYYjMJs
pBet/DVd0cwiQQ4ATK26je9Ywz6R2oajmrzMVT1OroJf6bjlcHgGKmj8/iVYKC2XYaBOcHvJwXOX
ucG7reP1vd1Odh/Qpp0QrM+K/h4fEX+gNTAYDt4c8AYiI9WDMnbD4CkeBNO8eIWrIqoauXvQryYl
iTr3pOu9uEorIQ4UBTGxkhqr4JEoOc2nVItWKI1cD/gE3yFM5GA17g/Y1D0NGXxg2ddxBY6axCcA
t0iBrIMU7NCVaPfKDCHyqsWKkP0IN+rM6c8ePouj2YoXOB41fYOi8ch+ECl9yEznnG7xg+z2ZZaD
d65afZDLzt6XJynGdNOIQdpsSn1AWlJK+x4DkoOIMuFNYx1W6xRQKf80z7zrAV1RomlwGolXjJgS
StGBSs5U+zqZwXAuEO22FETRyz1vozbrsr0RTs0nsIYD2XVPLbValXo3P/mSgqrbXSN51TbPXaZW
GcN6UE3VeGYYDRIP8J27ObBYyXmcQqe7g16vrLOuXNIMNZZE6niNql8SOhhpw2A7lALwKp6qr7nj
fGOjvmSQ2J7syl/mumDx0YC3UsQiQt/bDcaw8MmO5Fxcw5VLP9jK5h27oVS49Lr5T5VOJM8dTWn2
dR0akYexhyWBI7a/rSPig7CaSOh0JU9BhcCn5ZeJXSnMSBBEPHyGvpRI+JIaBY/gWn4uH1GE7xEe
CB2lGp4OYi7Elc0oJN+v8+82H24l0kIwTX4Go6a4hJUqymjjWWuofr/N7O4zOkMTLZOoxo0qERfG
epeo2aCvtBunCrLJVpiuywM6eCc55k46POZx43GIT1XvHbhQMTpypatuzxA2nax3zHB5MlSlVJP3
MHE2w0eWCEZJHg6dgIXFsVjrYRLmf9hRzMIIeP+BUezxAXBxYF/xvTymPeNZTD0PfWD347dfXdJc
60HSBk5xsRIKJCamvpB9DhxmI3oCUpWGSxuCL3pfzNLU70JmmogzsflM5bp8wFY04bJE04DzMKTc
E8lhM/I+hnlezBxGmQ7MBwx+NDf3yDhExjdhT4jIA8Ed4Wv1FZvlOmXzuBbc6S/Dy7NdPhmETt74
Yx2a3D5IVH2G2TWRPnM2ipxQ1UdCwa7pcH/3J6c7m+DM0cE23OFWM9xoHOa2k/0xrh8bt4LeTCVs
Q/I/PeKgWw7tYCAuwqqIAwfJZcSxKGbOtaSqQkfrjves2QzW0oRAI5x/DlqkWdTadwnf3LVA/2n6
0/Tlw5i07SsbPDTfwHRU0e4QdYJ/OKxHLFPIiG3gVpS4E/8KTLSxLmrNLxjz3cWFmSlVAUHlCgf3
YhhBGNk2CVM3RO3vYjbYIrHcpitVBD32/Acb1o6JgjGp8MwpHiWUpWmX1zecBsrL+b7ggPxmKQjc
7/LCA8vK/8lJrrYyXwYDvTL73NQdxr63QxF4iMk6O6pkw3lvW6g/wz6VPxW772f7lBPeIM7nZ4tq
bRQiWZzKTsH2mp/ZTDBD/+dOpoNj47w6fK7ciZ2mB07N5RzpFCdlZiDUt+8GANk/9FFp3WUKsCAI
E+hclO1RL9278+Ja+fccKj40MJfY/iOsbIPlHDjQdqX+7P5KWmDNHxH9c3GSrZsveFOlDOXxjDNz
QsHYAHq8EhjjdM2Jnw10BcK4zBOP82oeNrLFP1GcA1z+g8zhtZyzF9dmSr3cuRf26WyEZ8GCBA0y
OuHnmuDUyNzigyJ+D0SoBiUE0/O4SokbxKG2Ru6NWNDEvA9DXqAvVH7eQv/pVtjSgClWg/wIA2on
WJEWzrhyfRRZHppl+olgqqggFAePhsYhAB/iXqyH+2RtDv/B1ON5qPYRv+ok6HeoUKKSlL/4PdEr
FFrqtvDF2zNIho9K7jSsocbZfG7/Eq2JC3AiK0EOIe2uio9NnE0DR4cTkdlwKVQKQbZNXWhN7sBl
Zsmlt+xVS52nffJjqARmxVNCaztJJRiQ7Ndqd2eNVdnd3AHwZgkASXBNgLJiMuARKgLITRGmc4yD
8TOcMIfvdvuMhFTSQmGEg+NDpOQt3zB4jWdsyQJQ62IX3wdCThtHTb6NJ9fSj2uL69YlUcpRppu2
Htc1Td9IoaMhqRQuq7KtuAVuq78i2Rjnc0o+O1/FC+XzgDbD9KVNIW1149GhZY6YY+4hJWfTCA9L
AhyN7o0P8KQCaw+3njcjeA8nb71YztBq7+Fy83N0dQ8mLXwlKbL9+GP6QQwA5S/mQBj4qszTxPFa
w5h+GBdemY+bLjxprJe76T9IiF9XgyALiosxIxbQfjyyelitocIYYU3ycKh7YZHTfQZcx0UYT9Lz
rRdJGfTxqh0XQjCLTHvq8wY7Ga+bMTMoNuWe45RC0+RT73LoUhkmqAWm0ElaTBfBChhGapOAKt65
xE4vS3VApGO9GPRhwf7V3YldaFL+3hymV7jTyFtvMyU3GUmoO3tKM3ZK7ZsCOWYLzl8D2xAapBlQ
oCU6Y1Q/XXSvDvrJWC24rfh3qJpzTRO91eo4MxUzM9/WXONDn51GpwNDTi1hc6Wx0aaj3O1w1oDR
xuCGBW9BAiiRODjZRCWMApz0YecN7InXt62Xz1eLlK9VKnYdn/rWr1Rgjo1jAxzj5kjgTNLlJJjP
6ro8Kl78e7R4JIJv+IBceR3MgdZejXO2StidvqmXGJWUb2Kod2Jfd8LkLIxWACl+Km8oRfhOggmE
j1P2swDWyKXp1/UClTC6PfHoZPA6dRRnrV+E0GK300NTIx+POegERjejbBtHIw7hQQX5S0YG4hk4
DO7w2Cm/sOfYgYr6wQeJsYb1tXYF+/bF+TohOh7EgaumXmLyw4yhvgbciIRbKejDBbbAKfz2ynIq
eoIfh+3vVYNU8sZkZR8CL3It0qVzEak4A73T60QCCO4OAxZpi+g+eG7s7ahT17NY9CxVXqnA56aG
KBko41ZeihnwOfWYsIDFQC3faURP2AhiUFV0KVXqjHFaI8L558xe3V5yHVibLugactWBxYWNYj+M
aU9s0cTZkWwcgCIUDD35yUWv3mt8E9uZCB/eOIZvqZi5cKjxz545pznZ9dVdxpm/6+5seYl/IYsV
0tOWoaqNXstpUJu+FaBmVhW+RQoi2GWlf/wKTnN+0YKAnNIKuFTKlTKqxLFZd+KNjinzkZMTyK8/
cMBvKToDDyxd7mbLOrDZW6h+B9QY8BN+DgTZkZrBgGBl/JSGcgsNLlkcEZFPmGNgq9LyNTpL3d9+
TJ4ZRDl7gTenAFnYjJmjkoSW5b6z0WcTLTpDwUO18KL3+b6TAO6DNbgGaeS1jOPK4PHMucTEgfIB
pXlFcJGTRJpm4Fiqt9b4lZMUbTFNMK4lVGzaIQ29n3e6eW/vIZdHe9QObyQ5iXddJiQnyQnhKXIf
u9w3yZE6q7XUQ2NYhKYRLdsvIJYcE24KtXsh+7cKerAzNY5BeJifh/w+Hoi5Fu6rmjLnZNKPBKML
2Egmoh5YrSJE/1hxAwjfyjlqFM5H88nYFmIFhen8ZloO58TRseiy7cfwyxcud+TaIWzLBodnf8HH
pYFfRgbcHXVZWqB3SnnIFIN4o2iyOcHkMNo3iEIhZgKfUj5jZgZmNI4UBWOjFtJP+iCfi8kpi8yv
nV3G9lErZjBaZslQ1twou4Y/c8l7lvJOXB6Uvu9gD7+Z/cTrivU83MTPW6O0n6V5oipQBpblMY7V
Jsram8nFVA81uQsq784AA7335QJMZ8Ic/WmpGG0894/o8WcIA+IrvvJNne4eFefxGHzPm0ZTHNtW
EVA5XxRyWx91gABiTYR7MK9Ig/kXK4X9OVwXom6B9ntSqBTkBsB9A2OJMaV0JsVuwZ5tRmVQi+1h
1zGegzCg+gxoaxbQLMHGkRLIJm9ul++REQ8WuDf/W0SghkXi0JmVA2/CYzzWZ6RQLNfb/wOlQ2X5
KCLMZtJMhmmvPrjbg6fOaSR/KZdAgkKMka/ObftbKWFIkdRd+jTvqaGeqajC9u7Hu46jl3LOLXeZ
WnKAW87irNg3fiyJl6d1JQpH58oCChuMjd0gNuLYInBaCy5igM5MKx+AFzItSo04cRyBKlCa2vqp
HbYMuyD0v8xQyfVQScSZRn9VxWA5zrEqKYf3dKndUwTaE0jd807IkeIoAjepGkXYWn8HyHnTtNrg
zEWQl3omTP1j3kUVt2SUH5kt+RzBlFjx0ut7WDVo/Mf6WsFZqSjt8pEt6Ve1q+3GssgJF1iUshE+
I0aIXW4sq7R0byR7TYUrIzoa1bdsPm39OvmGrFsDpV9n19jO+9xOhQWuy/MJBzkOsK/U1Cs7zHT9
mDnLH/6ZnaNlJVnf3u/vA69IJBKjaliz7IHq+7NdKu0JllpWXZigsIrLxzU29mNx6gg3ort6Rvyc
71JJcWfk9O+gYSnD14EXfFEXyWjR7hRFEzaoDC+w81i3TIAQzlF7zTr9gNynyJoauXzPH2Yf7Z3M
sp5tyQRzczYhvKxptY/VbQ1QdNDNtsOFhiL57clmEotAGTGbKuGPGags+kHKykJg+iM53wnmqGT0
EnLE+wXnsBBCI33TVH6vAYL6opqzPT80pP4UQzglSOkRvXCkzHsTI215PubjFi1surt8m7zIMkhs
b0dn3jiwV3ANYdkP944qSw7lQDxho2RVQzyHgL12nONq64Y8P5B0mRLDLx2eZseFychXh+SoGlPq
G+pvMr7jLFgNvTJMko6GSxdbsMr0Of1a4DNlkHoBkwsv3EstrU1W9rc7T3a0BlObtqrpOf3y1dGS
sYqUA+qc8bfljAJHWHRZCBkfIRPf4zSxvoGNWQjYZ2crbAp8wkXuWeSmh5wD485wD33fA+7NRgEn
J7kl5SiiSrnK/tS5BSytnShDH6KAmPzAoSMFAw6u/6JttgopQAZ0AJdduUgke3sk5hM3ncpuE37X
vUwGlSlbhu55D77CDZLnPcepiipZRqohd6C6IUcgTmlme0zrPDp7vkOvavfl7BdY4GRD9NI/USDx
RTBDezJRMY8uDtCabs8LT0jzIX2e00T6Rt+EaL0E3Pic6AI7sAv4VmwRRnC+/yHetdzL9N2bFsEw
dsdIokBavCIvoqm/4LGrbw1g7tsPULqcRT4/fmvynonlBYWvPWYq/Ga6didwOtif6UzHdj6+gL7+
oHu2GI0d0zH2Xy9GIkY1AztE6NJG9kYGO8nF1txXmD0JMqK1h/nXzr6QZk+oM33Iz6H1b8+DAk33
KhuGcWP8HwCmL1jYTylDvclH3NfM7nOaILD1vJ1Lsorx/GPfmwFRORkvwsTXtaHgd59uBJVYrbhg
YR18iebbIHqfSETLP2hZUYT1S6nt4GqkPik+w11/TIq8cLNrEcuzuHUzr5nJpEzVDBftuF7Vgfq+
pVF74LyhmUKIQgKe93L2Un+zk3hDB6LWMQ2nzcuDy3sR1HJoCYYGOh9ZvyXh4/6iWpcU+eWdXqYx
cHvIW7zjYKOgsEus6DVaFZ8MWb2lVUMtgk2YNQOYz1CqrwzCOwWJZ9doccTHnUDG4RrxKTUIgGnE
pjICfwp/kgXu9D1a73dg7DRhNl4PvvgGtg8O9ltLKhs08ZljbyoN27+Piqz6CjFgoBDnWgbYaWkm
9aScfao1gRpks7XEeDJLiuit3KQsfh25r3ljk8hUn5fMrit0obszPimqJFmFNc0om8YPbkCZL9+g
1LLtMrQ4VJmwIAsXe/BNJSH+YzoQp98BlVB6ec4jOOotwOZbMs1inWww0VMiKwUrJTxy1k+ekaLq
CzduvPaIcV+5jKMBBnKKc5Zc8vyP55UPMnTTLRxZ+k1K6jxfpKPQIh+Zkm6e+9tKV/49VAspQGdf
7PfnFdcMIj5TP/fr8OMk1fNmjRUSN1hA7l2vCwN33RhK+K9j5vHWG1bRS6QpcBul5+JWsqcM+8vi
cnX6k5sPzPeF4UbIFf7a9eWu+xMUEZz1Yp+/WLqcic1NpftQ2FvpXruHBJ813wbSXqy2+kBjtUMP
RwSdvXhpBnRKC/jyAQW9m1Bq/NgA/BxB3klx6tE8n21BzDpcIBbdNdr2XKipXEHESOTmwUs1oJQu
WPKxbmzWjE0xTK4XhneHwQ20G0hls/n7+ZP0xWfdgx46sALSbB82v0hiCFKGA0niIscd9xTAFKek
qCMTLJzg/d7tOEO/O8lrMTxeJ0Hs/JC+7uOrevvxm/lL82LfVhmeTVyg0+DfqbFE8d09MV7bznT0
lCG4QtG32/3GGny1MQz3CDxKLNhP/bn5H62iidZB+VR5e4/6n+Tl8skfwGTHUkmeGcaAbCkEfW3F
Dr7mzXFEbaF/qHWNUntz0L96mYa4XRpAGTyG0SRE5CMLVahAl/CwcskJDZ3aFXrtO03et8qHqtPd
+e7umrk6tbs5BAQ7YSa6Z/D1jXbfrvP/czLb+upClqJNjJNbOfevNLhcWiVW91xMggboZEJ/tFWE
sEt7OYHGr2Hs1aPB0V+nZkSV+3fnyyEmvjHMB9segXrzU+uVMf3F9BROh9b7PFbwB5hiyrR9yeMD
kt1hRPPdzvc0WC+wcXraCRsf/eS4fa9PTCkrpa/1kJbL6gb4eoyg2fUWcd22WlqXMxj3U5q5zMaQ
IHyZOf9yo6cHh604zcaGTxYjgVwF9/yqNb9bw51+HApKk4gPqblj/AUHOJiDIZKMFpWnIEIhS9hg
ZyhuYnC3FDCe4cmJWZC5gGc6G29SPgmXcTCvYJlq6vySEMHtPSn623tFLEdQdj0xIKFr0/uH5/JN
LnRR2oFnexT9gHwXMtgHvcdU0Tqn7hIF4MDNmbZbKyxlSXBkzWrrQQexQZpKbqhpqzVTAdSuD4HV
TOySd87cIWvT3RtY4bHCHw20G1R/6xs1bEtwhU9sPxNJJKDmGwIlRV/2RAicZX/3siWhye1FTE2o
u6gu6xRyqnwYf8btzWxsoVFudPJ7CH35pOYBtttdB45mxwKA72jYqkrzjS9MOhcMVTC9qbOfUxV1
uTcrIH1lZGc/gmsWnL04Wpj8bhvZxQEYirnMKRQoagbggvluY0OafUQYNz4ArdbY08xO+zG4HJ/Q
gPjQr1KNlOPzog70vcsxQyis4/1hPUO+SN1sknoYGsG5sE0UR/zK6wLWNisE9eAUMnTbuDHMOEJ0
lPTsY3iUqaHOyEgaLYfSN96gKCT+pfAIUb9jszbe2R+fVTpsFFl+/9sVrRO82xjrbSzGdO6MWJ9p
obPhFrgYW7Q7iXOQQ8trLHqpIWwLmrJLhipjYo7saXmRYgKspUHzyvEim4oZcr86J7MfIcAqyZAi
+v7ncYf/wL39ENQVSLixPJ91EYwe5kFsqxN2ZfarjrPSg5rnFT9otzVtfbLGO+l3YkqtkiVVRkMD
cMWRryMrcN7ZaZQdzcRLAyCZHyqIykNsvsALk/sSiVDkNEcYggAlo5ZIJGHUjSHAMDvds3fq5LS6
g3ZoP9o5m1w+c4z5INQOS5CtaH3Tz8D8lnJsUzItfCbn/hkB3b9ypoVTuSq1TjgwuEoS0rn0Uc1o
gKDryBnbx8qMgF5JRkK18znNh+n5XIpWs/qEiWLUaIuw7UzLxdFB+8p+MYqqTzdamYahjBVa/Sqt
/bfyodJ3qjlRcsAzjm7+awnMXzhcfXS4UnhJTiOIV05m+WnVfSOmjhjvm4ZASNljneqD1xt9M/0U
/EV/EpWqvq2ZdkuQLldFMXC3ptZHfrnhtmrmIwgqgTkkcbpu0xVcsOUr2oh5VTv2Iv7+5qV/gSs1
WMPXLSv+CVToCeucz9VrSKY9lN5rKzaPp2dbvfRoDiOTGzE6mhH5abedPzgvwrQlm9cq8nUV59/Z
hJliIOT8gZoqL73Ermr7kVdpCFG1T2Kl8Sbd8Y/Y3YI7XXpggBXxxMpKUZXeOrJyJSOU/iADDPoY
1mSqaCLW3IgsW9yNtlwLMxQ3WaahHdPqeWz3L74cmooDcMEXNVy5qF7YWgZIP09uy23/UGYv6vvl
gHMdMXYsHg7vQbtw4bupKykzh6bjk2BNkEkWMbcNdRfXwr2feQe1hExrzNQshyl4Vti3++4mSyqn
IVMEan3vkc+DBM2Nu8+xnsYfztlGE8u898JYLlEAdTUbI2vz57jAWaRhrioVCrUfKM9LUl32h08c
HMuwIfBZjp4M/U76RWRWLtXTTBZC6yYR5iXDiHdGJjO5g27qxic9K4zn38xvK0SBSmVxZf6O7QQo
MWz6tw3G1MfwiFxs1jLSVAIrLzBPWJ5LDCiP5Du8T81qk3Zcdt5Oi2OrEJCx4gZulvYrfi9SEZix
sJsKaw0GFysZwDqlm2nMjEMVHWiOH52c76YhFr/B3mue3nq8crTy97/5io+hP3Icspv72Vz0Dqly
pnHbE+kroWD4XIqu0Fy+BeKBXSTAaJNqXI2x+4FafU3BmKtG/Dnhgvni/ZjK7GgQYnCqQkPCVhuj
O6wJrZ8emOE7+t1WKk6D6ZGxyuzjG9X3OW+AlWdr1ub3BqZ4fkC/5/mZEIlZvWNZEt/OKGwo2K8c
raTXFPICrZ9cFY/3uM4m3XFD4+AS5DeRuGwXvWiYXeFNpx+r04QMI/+lsMBaf0mA4Wv9BOxnlnI6
A0x/4bV2u0TAmC+aVoDz1d0q4CZMyolNjN/aHqWWiqVfnMxNORk1FgjQx4tM4XLvoLcv+sQZC6vQ
6eeAVdj5H5b8RA+YQSlXMcL1eym1tnh4qRvKxXuqb2T5bNDM3LRKQ6HLSOvRZANTcUg43TM0TeSP
0WkTZ36tz8Cqi1Oa2tr2nvCREbfR9bRgtbFvH6CK121rEzp3pffd87K7yvL9xMATerDSm0X5nr1r
SOhXaOckQNA75vX0WC9H1r1JF3fhFk5x7bppfiEwuultMuA8R5qmROmiANDBu18gllEOc39TtESX
DrXis6jMWLiAPz6QwAcMYGsJKhuVNSJihWWBk/x7/mis16vjpkPFaXhf5ltEUnYe1kByqoxtb98y
a9kNKbkEumJULZQABbEl1tVOV+Tna5MICMfLGaLflHk2DGgiJrt/cRpEpIVcXKlccr05E9IXDnNZ
2HRTwEmK+W8p2n6tQ5MJ+GbId6YIN289UO7zadeLTak1VFW6NWyaE89QCn0HlH6AlDgqgU72vseC
siaCjc2vHi/I7GQokOkoIzG5G3dPq+Wg5Tq9US6b4tAwJT3xnMgYq87oLidLYiGZq+FL9pf3xqF2
JsnQ+/y7k1ZvFcOAgZ4uBkw4r1oPHJcUiPgIP97cFSmDyUhP2Xyt72wIq0O6gCq3Yd2truhTNsS8
4+jM1wT15MbJ7CnJIkUQWFm2pmlwv7kVClXYjKJxZ6J8a854BTPOeXIKqdIHV/wnoTzbjJKlrmwT
wO+9nqnhFdb069l1muMy4cQXg10waMA3KATvuw6/KCSuqD4hjCgkUHxNGeX0AzznTZxV33K+pINO
t5x5etKCQuf9ej1azsN6ND0dum67++Z0Hd9sHgAKmUOs0/mKxqVARe0zNhBx15ZBTfgkIGWd5owj
Kp9rf7FIPueHF8rLVCpf2IFT4RpXmWDo26EonTU9znMFbM/GD+/cxYL6ZKDQrY+ZmoMF2CCBji+N
H1jAdPCXg5OOobpq6gp+FnbK/rNRKEy3jAM2LBILXih2LdZ6ts+GdlAHJa8UfhBWJ9ufZ294l64p
nP89xsLHegm3YS8VF1mdVENa2MNFo1z4OxJRS+Ug/w2p/q5zNEcGHhWqmOZ4RTOoD12J0bxI1Zbi
5gTSlAoZ5xM4zZYGFfm3v2L8LGplITY7tRpRuq8qoHnGxGHSX9MfKLIfaX9z4f/5LVzENeUGMHvT
jgNzzGeHcyVp1f7Ka3vXTx4h1kvDB8VuhqNY5K7jG6kwbvCfpzfd9ikNPhSoyjysv7wJ/sOs6qJ8
CAroCSUEws5o5+yShlDV7zl6qbgqoWkv4Tk93tuQU/zjGGBcm8EofYGpRBh2cJrxcVh9+cuasyVh
YjLjyaJVzlJpBAHCj2dHuQ3JfWlEDSpogfCfA270A6lvyI8F1pCjY9BICA4eqm9ofbh+IMDtkQlL
LAnbDuAjJ3wjoQAlE98f/yhQAvPI+gXMgaEUm4Vv6FflO5dbmZ4Ais5yKfXzXksN29vYV4AbtKKi
oCPt7kuVqoZmFPobAEZC361syx8E+vIyn4n6jBIRxoac1rU4ahWkD4RtNMXjla4PrZReLd1VDdOG
NqEXB6kGkOe4GiTKoBr5+kxuV67C/CZ25sm4qlY7PXEHXz7Qa1mL33Achdb2nMTfa6mL1f+nGzB4
UWh8nYTj6XAmIhlNXCWuYdgVorXjrj3M1HOiZIOdBNek0cane6elQhkUVMxddBz6/CDYX4a4msia
ixeViNWTWBUfSkNpvznlOyyymJ2i1y44VH89TZ1+lNpVFI0ZfRD8THqtX7xp1DUyQgYeg19hF16+
ana1Qvhmwzovp58vIz7RE9d+/JsMVtSmLuo6QAa45uoPzGLvTqu2FCEl2kbi/eBPSuYA9+fsN+t9
P1veGi+6l2AaNK1xtv8hAL3HzvxcIGZAAGuAyWg8kKHTw1rYQVAgM5Z9WtT6jCBIhw64E5V8T+y3
mIpVNxd7Md1Tr0oiWkdpZqy1c1vGGCebJPz4k6cUKLeV0CWNoXomn9hRooia2BmgmNma5wrUSZtu
A3R/31bmey53PSnzoEFGgKCH5XcShplx9FF4ByY8pDYYgANwjBlA6ym34XFB+pmmEuTvdGdaNBHv
cIxVH27ZkGMte4n6XHUVXAj97YXSFZ7Eb/XfkTyh6gt6f/45Z4xFl0iwSCmhvwk62EKe6/RLjutm
dzrmOxq5NZLcAGkBxp0M7OvPRlFSTcGGrzDNeAtkK7Gz1K1bE1FfPvUch7ofn5Y6AYXJGiXLWxgX
ePc1wBIIhlsDVc4K0n8/TnVaOEia+k7mGaWEbu3lZj0Gkhhhl0aYuoc0lQF2c4J2DFk6zXn/mNGX
cFnYE7aTnOyl3kaiH+otxprl9WkmKwZm7FOdCnmhhAhICpYiGYAuEZoYmqEFemcxVHPdnn6pLn1s
VZSKaV5eOm2wIlfORXnzfXxfIp8AOMHl8EqESWL+u/x/wu3zmA9n8RHv9mL8J22Fm9KOXVmobpI7
gpM5HfM6bysthIQ3rUTlg4mf87C/Pdbfz8sv+Qa+Qkv6wicW34E+08uPyJgG3PN/8z+HkqzRue3m
/A1ShjH2/I2IQ7Hril17lfKK3T5e0TOMbMo9jEMgyAF5gmJocg0t6RoVAhIWXwHL4hw1EwKv+eDG
72AuH77z8pkBOjkz2RQsaIi2yt0xVPXJ0W//8CaSp4Z/5zcxMKhdAVrQua0+VHNnRrR5M9xZnd00
PI4A1F7N0s7IeiMthMSREI3DFlIHfKNEo3PuWzjGy0ZXOdlZodcD3aPpRmac67Rem/Jia87MXJLS
t8w5II+wyhV50d5MCCmLdS3tcJ9KvnavR4KHv1L1gAgiRQQIIlXg/LUB4xK18a4ZCCj3tgOHqjWa
4eqW2WFistEVC0iwZ3TqSIO2JEVuSfMwl8vpH094cNdPoB4rktBGyhYp9MRJxJRGQlcSV/GoXtCN
0i4uytgR/sOAevcRG4R7PPObOT/x22XOvtQq13M2JLz28BsJTEV6ctpeNbx074kLYFICy0TPQwx2
wysFXAaglrXEjZW88XpAhLOm73dkke7rgt0lKzih0Y9CAp9qC76Y+0kct8vUGYivfZG0tW6JnU4a
Iecm8BtGqqyiwPeeRX2xEPQZvm6N+PyufMLycVHP6nb36YgREaA7Rt691I+KO77sF9qf7e88wBws
CwnFP0hHUuUG19CjPvPcC0/Pb+z54nb3zA3w9A3dXSkN3kUwMVyF7xni4HiOcvNKi38WRifUwxDz
IKwu/0fzRV9kzHzHVy4NfWtxPQRnVs/7V/gvUveNOZZMkUWyunakcVB1V6BdlqjxEqPON9z/UXrx
b/KzTBTHo1oDcrDUs5zr7sE5AjbGYtI5lD3ti+QvPIyeHLyTKSg1yiUGJBLsvqGtDGyFZ0SsXbhU
siXClnlEOi8Qr/0i2gmclPPxGNJHzlJhJx/S026Xg9g/RlXhJMxlOjG9b8t1nYw324fR3eZhTpBY
wAuLifnGu4YqnKW1YlRE38DXoUlF/H92XQZ3+xUgWFeVTd68GFkKolb++gN4T5Uz4Z6U5yQmKhZ8
KOz0A3jLfa5iL2twUZhXOnfbp4MduiKiBJguP7SnCBfoPq1QwzLkG5qWjOmyVzNiciBo55wwfVRD
skxy7Ci79dvqyozPoun7dHlTp2zDthFUdK7bVs9idHG5iAJG0icddcvveJuUuA5245w6fHljegmH
UPNBYQISIMu065gVq9Mw9DXiBAA4BFU8CixzlGCinSd2Nzz7G0YXr5X4EVQXa0uptnKwHg0dUBuB
zJUyNr6MmF5fB+UjAb6+FJODCmVpskxBLsW68PMC/phEttKnlxuxxvoP5CYlfvHKOfcUWRHDAcM2
E1dZYYT3lc+JKagr5XimbGMdNyh3WTYcdp0EgiDLmZfpIMzkgEc7ncARXxUm5BU642cL+7NuLHlu
MWzjWISWpLzHd4QfEwKexRIzsee/tQnQZ7sSyzmSillYKPiISuhVUgFZIey/aFZwlNPjvmzDO1QO
czlKYjW1JKtrX/m/ljsoADQQ5Mmw9cIE9v3jGLaWn0j0LJS/F5IwKYJkPj/SFHHH5A1Twan+tNYj
loLdFiNw6DQcLRys8ZfD4nHRvsu+Xo+7NMLnfXCDJXraLl3iHcybxTz1cCLBVzhxemv3wt2FtTnz
8iW5KTZfxY1tO676fMFQekLdc5WCH/ffx3/TrbamLqnYK28J0thJPfWJUjNZ/3Un2/BqMZtODvmv
pvJ6A5JmSDOO0jFxe5jpnOP5yT9fTVg8UCj1E+O5exDyhyzdy9AnNqNPhEKHKlBBDaEdMit5PXa3
jvwPyTq/rCp1K9aFF3f2965AF16MVgOAEZK18BTLVJfNIWBhPsYBfTUG3ZGnLCaywbZvlSjXOBnc
l1gwTZat1g6noiUmfbuEFPtszpYXWnj7lSc5I7Y0u0S4cwZKX9OEHiArrd/lUYd2+HAH9ngcuy1v
PfqrLCwst1litRPtupARNPxr6r74GMG3JlAvUjIcm0ZpitfpPvME8v0wfrqf7kM2wkAw6ZuGPEw4
Z1gZGkuNGC23BDVovwmL2yH8FJ+4TWSxPqzQHtQBxBDlJOlXb1n9sT7Aw8nosDsMRw7Z0Bgwu2bA
Ik75Rv24NCREim49X9ZDkQ0x+g/lXzSi2d49n88RFUjFnJDiFDC4rbKVbcZXo88aZQeWe5AJZmNG
EkiOPqldualusET+e+qemdllUzPxgZ7fi/FLK3Yg9yX7rKIQrWKIA0Iw5lcWxqLW0Zdr3EaWAOSj
9V6zc8HBvSQBSOu68/98XPGZfTxXa4Jute8dGv3hOC46mXc9xWh+pHXz6ba6EWxGq6FHDv1trpMn
BoEImuw53AlJNkBxdzaF1wc7lGR1TzXMmX7Y6mwcix+qTqHTeRG+FO7ISpghs2XcMshyPhjLaWhC
Va2ZuWnA0KtS3kNmkWmC750GcxtfjgRo1LotXar81Dxs7m825w80RD11U51QONTElhSbHNIliKay
L4S3R0xWKaxvqNxzUVTLuNoMs9xZDQWl6fvvwMP5GossP91Bvye6ag0Pqgyio6UgzJ52NSveT1Sm
ZkIXEMch6etirXQ4+w/AvM1SekC+ozJ1Rh41m6zmrflSlJXZ0mIBg9n6SrKVNZWu1KK/kJ4H/A2G
LITqDn6UxPaAqBMqialtsXayPBtXNJ538aaPWs9TO80kIRkxBLwC/zTuzrYF8lujtRaQk3OgfXDn
DhJ5V+xkAdtyd3jhP8YIun1cOuOwD2psSJaiIxa+EcSMNmidv8mRMV4yW+GL3kmqMnxx1mh0K3Rw
aCyYgjAdq/x+10M2qHmvxpQd7c6ef169LeygcjRwZmeYvr4Tv6yX7DPN/jfVMkY45CmHv89ft2K4
mLtvS6mypCgZupkdhBSytegxvRxmw9ENGlnmKQpDTx3pUpQ3UHrzP9W6vd7qDJO0Zy6yL9/hXc42
9YLbNdAqRO1u5qwVyHFCkyAodWJndZoNrgdtlD4tfCvJHUJF1uF/pDJxQoTNa5OQsw3YjWQz9B+9
Y4w7/ui6ySyJv31jPEYH6JHbsoElRDNWDMjytF3XaZ9wdY6APsBAHPWF3JkfrP2DaNiYuaWzMClx
SUxv194CCFHwlZYxuvX3jYCfM9lkWjeIUj4BYqf0l6e6f3EgvCtCKgBXzaRiKfQ9nghmR4tzFSps
/hgXZD7n2yh6pJb1kGGVnJX0GzVbAklKQBW+F03KzHCNmZPf5PUq7Iq0Dn8pYBSXBtrCLdxJfpXG
gucVId9eCHkqeWQbCyMhLu6STZqnHsb5080g/h3O6vrsblcF7xt5jOIEqal3bJAwmchYlX8wWxTp
eZzapPRAuU74bi0f6VPiiFufjWkIeu9winzCDj7lV5dIhYG00torv0EBMgsGB4a2pAtxrflihdzQ
ipL8CtIwNdR2cxA1HZu1z4mG4C1RwRWXy7v/O5ipc5LkYb+WUD3ugXoWI70M3R99U09F8+/zfnA3
2SyqiXSCxP1X/HTGjMFimGhH7ZMlaSUx69n6c7dkaquhvBZ1FlNvt1sf7aGbSVV4os/KV0sRVv9F
MKK8k+PDqCTjV8STfxJMO4A6D4J71eFle+s/G93id5Yr+wqUNGjk2uwuU+dygpQIsHEDklRPyvE5
1OsmNI6BqBYjFYOe4USNgsrxGLuy6zhd04ZjJMU1imupIts6N3OH+o5p3Jr3A2Y8m/7/JBB0QRpG
MCTXWtGkl2ajr21DTwejfiF0rUPCUe5TqGIte2lQVSFYLIBDBu4JjS/8ZyujpsaXG/zTVXVy9aaP
CQ+k7treLqGKvA7NLLyUAj6SP3W9/e8nFOSzllfUYPI9MhtvH6gM+k50df5lrOn6lGsY/3lJ6MNY
BnpURPTord5/9UGekBFP5/vg7Xf+MAn8Q7ietJ5VyuA1HTcpSnAAU6JSK4edKzGciXgsKixRyrLa
Kyc+85t4jjp2774X85Z2CMZw7VyCAQzSp2/uXugIFpfcVGAFhTKab9zwAcktoZ3hzDH91fIdaHc2
ssakCc5DMtmZQrvrbQW6NKrYpMC6l6LPxaWWN+RKO1TK4FB8xCqj81XerOm/w/+lw2tFhtJOEDKa
RQspEMyCFNAntTVgXSsiRFN7BzNM9dQnloaEzjKvM6ocwZyy4e67107St/K/7Sabr8QVAgqt4SEV
KtyajreK4jm2vLlV/97m9eBKJEwUoDslcQ9wLISHsRolNutuQARmhoL82KKpALPij2B/gLvv6vU8
AnwBB+7CFbefO3jMAFvfOvPNPyVO12xlsQb2k1q1IbfmFt8wmajstxVivakz72La1h1WswUoPiiH
Tkj28Jm7H2uL/StmvDfXDuqXW69n1LZr1lFeXTRk4t0KMdKTyEY5QROO3UY5Zxx9Z/aNDepFIBI3
TW+fzZBOl9L/L7eIOMKL9ruaGTe1HvD2MpsU6L8mSof+kz5z/ExZ1lGf7+6LTOV1h2LoIZPTJDqf
aLRea5aOUdnPeJdOdyr/N/Gtewqhp/dDXINdkpK+P/jvyPiKeL6UbcmoeuIFpt2TKWGEXCfOURl7
E+6slrF9n1yRkVt8EwKeN1VGSEuZnLE9BSDjsN0QGVPuft9k/dNW4Oh83YzaKko3v3fTUVeN6ubx
mNDcQPrULDZ0JkDTHoaQGQS7HqQAwbO+KYUBtnoFiKrAaws1A3yq12cAVegbXcW5FT0PSFgCXxKQ
X0kYpYSgLeBQ067632oNxCY80orsc1lKkOTN8gkBuCg/bqZGafVIEh6/sPgMRF9nA1gykUVgP5PI
sVjpmz916C0CbgNYBehVxUEkC4/qIxTIvIoG2tv1sCLbSMRXW2+Y4w6eHRk/7jbpcBa6KSSIdOnM
cAnxn6Kx6FzwzR480/XmM355MahuxIpwK0O5E55Tw+CGBy3nTAGJREOCrxlLDuCKyv8FOXomuEZz
BS9iIwAReqCu8wEnqZIDmvDphVwC6VuDIjqb68ab5snEGw8kAgjLda3vJoPmZ9yYIXoHL6khCehl
Bgbwq11QhHY+RpIMH/Hj7MzyooYhh3Q3fX67RwdlaqAIt8eqX602d85wi77wwctwMrpJ/70gSvXE
7or63vlAkEecQVZ8frCeMYaq7pTDMV+Cle/pN94FFQ/kelcoYoAfpHKr771vsk7TplEepMRsNULT
2VIA6jvbBRr9jN7FpHfmu3Fo1w2nkNra2qBiUk2QrfUtkEhUJAs7uOQJspS4WAssOIbYh+VkUH6g
EKwQZ7NSMa/04yf4DY6nu2GrimmMd9BUYkYFwkj6K80RQnjvKETNqpj6VeeSLh9/SjIxwGp/GefY
SfeyXNsq10OqO3WbD49dSi8YOK0TbDgGiND6zNMxDeYIFokaKnmMTAecR0gKVtRPJ7z/Q4Vq7VVv
99AkEPKiJv1Wcpwgp0SGnKwiVebA3WYvoEWogP6ZMVNzqZe6eGm1CWbgmtFj1u1Y2SAH9nk34ofA
Ve/r3lfjl8+Ys15bqxWaHglrinTzlaJuzaaESSP2UCUqZyWa5wMXN0ZNue0YuQ6OJzwptMu4obVe
QuRFngd1hHn5gbxbDY6ZioG+ANctl9jnwKxjDRr2vrFEAblXJCnrqrUe2D4FN4mezayincgJbcGl
a73vxRaDPJvw+jPrE4dpPlDCInC8iYfx2ZphxmucwG8Bg6r5uL5i2JaBUmuu0rVoegHBJ8Lyw4sr
jAzr1ZSiz5MAArRtI6IpR9a9G9C+uv98lJydNvtkfrLGeywYOUeHQNuM3m5kr2fEcUoRJnB8NdYL
sasFg7ZRC77yelO/mS/BMvna6kpbOIb24ANh/1jH1xvXFQUmfI7zaGdGJ2gfvdza/gyoDUEbqM8N
basn4ZBr0bQdUXS5MAz5Yz1F54+jV4GFGIAdAnL68V8UHzTIQ69TLlgni7lgEvRx0P2aB9yd+wAS
zwCfIkZP/KgJIBnUc/HGsO4FQ9rN7sUdSnKqY9567ClOoqwdJb4mx7vGKs61jMhDQNWCOoYDAndn
5x6k7CMb/sYm7QqpHLpXYnvMG1bhWY3yw4YM4i2ez62efIygbhHxmDd3uBb2vPEqkIbkz0/8NSoM
bF5rcDQdvqtCLnWVFbUp757LCRnj452ei/peFmgntTxgh7ZshbukTrE4GLBHyyG93/AhaCU7+Cmy
YYDyPmKSIEpWYB3Fa3BXmM05xPCxBxtxoqJAqqaQytMQP/W02A5A/3nItTFeKSyGUraEZNn6fNfJ
8NiDOzxjjGSrvxd1HWCNCPFRODtqcU+D1qKT1UG1pVioxzlMKKzv8joDKhK/oCy0IwCqtNG7VaIi
Rnxk3gFJDsfcOMnyyof4SqTREsfjvG0/UE+3v5BOOuSKLBYtd6TmzyTGthRYOzIFEP37KparkAT1
i5R+gUOR7O2cozsrYu6giVMn6wdrqhKIrCuD3M7xBzaQa1JxJaYR8Wmn2xK+SMf8ud5waJilSI4Z
OCKGsYvLlPpye5eQk8y9Km2tki54pkZ/wWRHMT7fKD5Fs8h7WDSkuEhNqcBWQNmw+Q6ywc/pOJau
7KIbN7NIwecQRyPQ75eYQq+QnpO8WSgrn/3rOkP8Lj2zFVluvk9YnzWMey7uKVoUOqUrFNUdn0Tz
dVPJLe4kT1V2wI12x8zXM3q6pCIEaEUnCwEe0GI+8cOAeErjD96ljySxXG12MVgJNIur1J7I29LB
WhFjQVJ9slGXPqKVii3xaTV4xQWGLzXBYcEmBdI+V/DDE0wOOoDx1UlGqwgLcFLyYwlL/DmJ+Dnm
G0kv0Bz/wF2StBYEiYwe0b/qjG55rOOnaTkhTv+Y5EHaVB4pV89ECRgIYdKaELsHd18ByScmn6fX
fdUM/WgYXSzKe0WAxDiydDM8iPwOGHyIWoGUaB7B7hoNq+nPSZwticRV58QTMupDN2kdps7svdDI
iBEEfVa6NhE9r1TEfAZ7Mcx4X5K6TR4SGG83Yv5not1xV9x2z6Dt4UrPq++oz2iikzdbRDgufxUj
h2gLcJopQvKIqXMDxio2cCE6oK4ADbowQR49LLx9pGo2x+IfuhjY9eTX40WkoJP1dm+5lP0V8Elp
Can6fbR1IS/Ye6n9UrSOE6YFVGkAZVABiuTabS0XzkDTn7dElh2sj5VPAA4MlYiziwWZ7dP9bKrl
HeD4XOVe7z6ejEglvs8kod4ICVrG/bf7bTCosjDj/C1vByBtGj0Ustx/Viz9oHUFDp9hUccrB+59
GOgEGWYn+aUXcR5Rqkq4nvANoy6f9wVea7dApaZCLzsbtmqgV0RA5/nVywYdA4ce0LNYcVs6tet2
CpF/ck5XER3l8/uVxyHMwxq2q3jTZD56FvtuwlRsE+/KBY1gBHSpOImJDKxp46veI8ITrMuDqVGb
Ci/cPMF+D52F9Ph+C3nOlSGe2NhTkd3TYmaUQK19HDYEd43XVMPa3Lkmq67LV5rq8JzJTeYYkx78
VgX8fpR6P/Fqce7B1Mpr4USZB5sV+fLQkSb/PNX5Lxkj7CB4iDJisDYHpoiU3+LbyAmhhs0pRhB7
/RwFqGVf8gHPvM5bppr20LtNOdthTr5AVVWA2RWqX8e7RlykCTVXQDmQ1iGuqwiyggJlV5huVtNO
Bq7TxrwzOTqqcRVmOt5HJw79Rl0aREsAtafhcCF+FCkzE0UB9R97Hw4YxnY6rw6gDAiISfeaKnc/
YwroXN98gZSxxDzXBsQsEX4Ih5gdGOAjn5EOvn7JkLii/MHQ5pdzSrLKlQA4ROnGnBldNwdmhta+
jyVaAWcfCVcTPMj+ugr3RHhAltAFqlxIUSFVQbujpI2FjfmpY2TvtIwcioO2C1L1wuxUoBc2WlnG
N6T2fv4EfqUEgNbg6d0bN/Oi8e92hwKhtFG7Fdglf56QhAMRyDjp1B/EAf78goHf0jxbN76vIPOX
ckycxPdyju4xJ7aucyQPt+xz2uef/oJup7RsbXCfz/uWMaOX8qWbDcMoW6OcygwvgdKbXQF94Gpg
BiHcI0PMLzmz9oyk2weE2GXDqW5E+cU57iszB6dpZ5MIO1vKy36HcAsCRWWuTmenpipyM4e9cXI1
kaw9Vsw8PugDwQs0go9YjlNWAcjln9jnInkeK0BRYi9ZEP/S0Wks7C9LYsD0WBNvsof0xweHal/p
PoQRh8zhiSRXxu0kC4NOESbJFq1xzdqujBGxBsSt5B86u69V1iSYm1b3HBg9rc4Pc8TiYhGQiVyH
orkCZa8m4+MADYZAmY0+kyqpW/dfKB/T1DUkt0Io8kPaMAqF5IG1QKztpyhgpwKqvpl21OzJAscq
AOzS2YcoyLsvQCDq2aCNHmjlCRX6Rq5627hi6f9Xaf40vV1bi91+JIBfWIbRiqilD/iQRHyprc0o
v3uJEffr/5IInWEDdn8t9F5suDvf4mVrINDrvQevqdyVF80IZn5BAEj0BtJ2g9dThsIIWB23z/vC
oY5TTdvIEZ1QgwjReWmOWJcDAj81Nq2niFc58FQ92qHQxiZoQZGMl90FxmO9gSunOThyOJ3jznlU
awHR4OUknKcHYoMubL3Xu7Q1y3Agmcl9lFoQgMtqt7Fy8lYNS3yEtqRVvAPHHyQlFAuPDMTC10ON
UTyRURUR8HPDcb0enkL0IwaISfTmy5FlbYWsfsOvw2mr4LWVfVoyrZXgU6EDmYlgLfdgJy5cGc52
EeIxnYU1/V+OHQOZDgPSt9n2xBNtS4MCQpD3UEEEFh8xdfPZTDRGwZRQ0wsuXYsafS6dRGyz0Knh
fVSR+7loBSfoRyX+mfdt4gy3+Fej8ZqR5kQX55hT/4k1S1cRSfVqRwcHJXSle7R81GRv0TnWxBSG
WDT6aVR7WY8as9yWn520HIun1SyM5XE4uow9/3Pdkz/OSRAdwaa5uB4FKJjM0jg9aIjncvtPDzON
Ik340TundBKWcRgB9VoyfyccjC7smQg79YFtj5dhS20WV5wFkOqIaKOkERkmtX5FqCk+fykrP7I9
lDAjkc9gQAJgUKGX1r4/77ME/hTKhRJ34MAQFsy4tRH1JBFiQ07ZjdRKshLl5g+II94lRWJJIZX6
PTN22eLQzFWtNxc/hhVftGFlebfAw7y6c6NLLZtbxbcgaZ6ntAnWpbhlKk8mpHNUlVg2vxSdAGfm
E5V6UbzQeDs8vUkSNZCaou9qfY+ZjmnOWMehJSeZQLzkUlOVjMOHkD5SZ6oSiN9Uwh2Gd3pdNIXm
s8gMu7ekYO85adjD0JKOhVkVoyXrWEJtZnvCn+lTJauEXToEU3dKZ+tXo8a3Gi7k6b0ug3CMwVdT
Mhj/DV4GrHoP52Qk8YVjTGfNcTd8fCGN3kg3XYCXMCUMcfi40k18avp2Dh+vTnL4EESRGietJ2eU
7Clts9aop4ymyBzE3w7DahN4QDqlWEmvHt8gP2tf78jtM5m78/tzgKYI0h77erA4Nyq01fIKnncd
f4PNBN3R4Tj26dlYFUwIoqSM4WcATHxOyX1fiNEt4zscI4ZP9OTScRkKy8yqrNrqDunpRAPOiA6A
9QIUEcKU2ITX9yVyqlqTo+yeQCnWzHKJgTNCl4o6EviNSkxranxuOpj3K3S1vxx/h1PtWkfHmI8A
PB+gpf7vDT87EvP8DPeXignv+RZYdBob1H/sbNNLr1EL/4lAC1RsB66Zv+KKEjOXWwiNYNn9WF87
Mq2CCOxRZBervztZBzkQASIPWhvYGnC6W1/C1wiL8TJvIO3JTr2b78OZcSAEx/oPXKmRDaSu9zne
t0MZYCQAfJOpKoBhLbVl97XH2Dkd0+vEvV5cKzl9UTYoAOzSSrr821N5YEazd/V8VjIqxpOoDhNv
LyDxud+pq9XcM+CjdoIp+8pgHkXa0BDni1Qo+Hbfsa1hyrrFI9cI7lohaS6/kEJCEnXxVSDTmwvK
cer1nYvSFnfPsBlKKSZm5PBym8STY6RO3rVVI8Zgw69II8bfxjo3eePf+hxMdKDusEKQ4xxa2uJZ
MlYVCrlBCVxcg2BFVzCX6RlDA0VW7KbGKdlTLWkUlwpskN9K1Qmzbqf8LztlTubKl8t75DdZ3eRc
W79/VmNSAvNuRfaxdkRdWMrcKuPeETkAA/9+dkxW8/peUZAtxF7m/kd7xrmd/Swx+6jGvI9NVbaU
HpR2UQ7iStH6gaGPNsGEJdk9Gertf5/q+adaq29BOO2i7KJqBSXYJmruvs/7RwQQWsRbiM4GtbfT
AmgHCZ3SeVF8xMCPjxfKraAyLtCGp8H5BGzpfp8slnphsUv4nqSSCggUxeIJwD0QA6yYD/Ddu3jP
psUA9DWGRWCUPuukS3XW98PErHnJOuu7oTinFWzm7xXxpDhtKVZHD4CCszplDsvqUFyfxUOYY0+9
f5L6kWeKQ/u+rkSfSIFOwahIcEkHy/Vwo4M5fpkntCZ+COvc0GwM4jXga8bGTfLlxl70yDKPNDUm
6zhAlV0j9S6FpKh6N5N4WLmGwXKQEyz72VmyTZ30gj/Jj0WIMmsmiYD/wWHuLcLMkKoZjZ8oRXy6
uKsWdk8Rv7UbZ5OXWOE7LPiq34vGDEE3SMSDIsnRwYtLs+KceWGvG+qjf4+vBjRIhBwbIfbsKg1b
7Vpw/pb9bg22k4R1Genxh6EpjRx8nBW3sJvCW0q9UZpZPBESwQmU04PDOsXGM/GedDChtEdi8LNz
AWFEZely1hj39DCGx9TWGa+lyzS+ah/PcSueyjkMupD34I6nAPGXIgOJfRnw/G2T13u7dQBDZw9g
GtGNN/kzHYRHb/xeMZFw/rFDDR4XoU3ebayjIO3dBm2JofJOwp92AjLlzPTljRURz/5pneELDvrX
z2dAXJaB49wZaldQd7DhNGFy1ooFcKRaeCryJ6Wn/uJwNwy6GJCFSE/2IkQhsPxfyUV+0Ji+DOor
I1c8JCeZbvCNR8DJz15PfZ2hTZdayDis6YaZWwOo0QxffpKFXyvzukXBcJJ09/0kpmea+YyZcZ7k
0MNxl7idwRCrn5X9/Vq/ZXUUB3WBLNLgPw4KQXQKnwfFxaZgsZb6pyGlOOyHU29WYbIJ2TMJoToU
FrKBolaHtGpf+3B4/hmCvI/BMRiLMSn9jXdbONl0quaMN7zetRwJHbw6NSg4KOEN8PFvrvgXiviY
/+/93tDIPnh0LVR8vO7y6GHNj4H6Xmq30sOHbXX6V/Z+IicBGsj1eCz2o+LEMeNkFqopieXonGCM
FIwL7dHDbEYU3dNwFMlbHrzuQ3vzrxCVaz8UNmklOQkBHC6nfafU7D4dOJj3bGt5Jg/peEsLzEkW
WNkhvoZAjCTAyWfZIUW1oP1ZnHlAB4je+TksvjzIG1heqCV3RKvAQOiY/Pu0ce0q926uFEFdFL5c
1Z47XFvFAKIRkN9BOzgywdSlJAOfoynUInB4TszZw+OMXWYzZ5MfEjVxNaIajaAvl77GyiRUMb7D
ku2aRnVEalG7btcN0+fn41iu7KjHx5NPjNJVVsRcqHKS4Hf1QSBwJo2PlxwvBYqaBioP4SBTC9WB
KPpVOEMURfbI7U2s6Nl10MW3omygk/nWtL8eYzJUr6GzA/lQVvEgj9mqmmRccLHJm1k/d0TCQXLI
pcPhNBRjWVQGHe85OTY4ZL1Liy1/wWQYoyUyrD74mw1zY5eJkMQLoFajDqBgNzOgCnHyEQRnkSD0
/JlN1hxvA3IjO9hYvcxqmeqVrk3qXXpnBAxm+LMCqhqgNPozfyf9X7SgiNjF12fL8Hp5dy7vH0nN
qbd7bjw4h2XvdaiQeN4gIlj8UoQJKsiKp+/EsoNblT2KI4zDGzdPcoh4NViOVnpMWTibvvNBOZpK
wKOSBj10TCF9Cuauc4n3IaPNpFI0AittndPRNM7iD8hsXWCmpbybvYh2PlzxnYlno80bJXKHfdgd
DkWn+BVqJa/3I9yYE4UginUght/XfgMuesXqQLC1WVEgZ7bhi4BKRlvcTBxOxU57aAZgjeOrllPQ
cfyuZtHVOjm9K3K9eKtQgGO8u7KGFIQJYqMUIVfy2cIUjkcH7S+cDUTUcb80N/Em3N5pMZgAvJ2T
kcCRZGTyE/rxsIdahD7bUnw1mq3zBC6f+70nH8fUsXSsdBxQQ6I9pca7Q4juT90vVZCewaMLRy3u
lVcdfnC4wAdNpAWOSIq1yms1X3LcHCgSqQT00Sg0ZULtvt/EobSiqZRPXAfJp1ND0nSFXwfnAdfX
bKVV3qIXwHBCvSeoTBoW2XmjrUhmbatHu0czhAj4IuwL/3SYAn2jQalDgtj0EWDbJwVhXHHuk3q6
yzLenriQ/vAzvnwLuGBo9bGZ6aPqA7xb0u8FXxbAdDqMbrtox6d4AMwnVwjyJpIaqImfkia80Nrt
ne31PMcI/89a4Uw303m92OkQxGO4mTq+wZnUeTaFZLcbyWTOT8mp6upRlCmrILqNDoigtsF9inFF
DBOC2OxmzM5RXkWQuLgzrwD4ko6IKOkoRBkRaTbCYCrr6h4kovPPygJSPjJNbw3I4iwWgRRikJRa
WesGJdwzVok+z6eD7R3y9p5oB97oTrCIITBtW41W8hCA9GjyMWEV98Mg1O8WQIq1cgFCSiHWmEjV
XFMh1CcVymUmWtNV7/D+QmK2h6cHdun4pIOWIC5qbje1nziPJ19owHmjRCwcp4GXd+euGQ08a9PN
b7W6UT+uYDupt1Lc4uw9J/o0QowDVAygdn2BzQZ5GjAXW7QVPPq6cA2yFGcrU+Gh2dr9wfwsM0iH
UrUUA71hhHcKf8hsBySPjrg6o+wbYb2pthM6pN62+7JFHoEe/iROegzjGFa9RhlfRF9RbEgusw8e
RlSzTWUuHNI3ukIRVoMpukAGDq19R+z5Ni+QAxvc4In+2W4EkF9WnSxAuzh/aO5EQ3SE2NUq0XId
NwfJPh2YLCJFD1rCrQQb/ye9g/GZnPH4R5pw+8APBoJdMjo9WzlSrPqqOQJPGaleR8GfjyZWbML3
HIlZ4jlaLwhu944wQ8t0tjK+SigduvYSf3UnzozAxlQOxGk34OZfSub9RjqWkV90SInzfJ9gXdHv
00n9zj6VIAYtE4ykynp0e+/ugPQIbKfcXPBn9SRBEJmkcUHUyaHeav/fRsIjdXq4Ek7G3GRdUXUa
ksGP1KRrIqPc6AK1dhywZVCamzNY1ipcBJLE866wOIpKz7aCbWLIXf7ZHbc1tbA+OyxvYM4a0Gaz
R40Un4JzjHaF30aXZG7LITqUhMSYGnY1N77pjKlHWkaGiPfK9Y3bjmmNdFGBBhQm7A1rbdRJD9nR
PQz9/LgNxhBPAB7Vqvm4EX53ahz6/D3mL2kGdK6/iPxLnVuiX5H/3uWebHu2jmU+TEaJJUsoBpzC
nv1rHZL9FWSP2QSsbNkBV+4gkjkTBpVCn90svdl1TPNe6HsWTAx8HzyDgsULwZqzEYt4wjcwcam7
4Qb8g0iyo628PqXj2oJXLPTGy75fJNpgkyzpD3w3xoXa4NYpniGf0jza5LekoZJMgB/FigbCthKd
EORAoG7uGDher1MScjn+4GcjptRJxR1xvInuaL2a5WNb8/7FtRMVBdxY0btwD65QK7WNa9BkBkT3
0r/ffsVV49D7wB8p9yq+KYb0UFsmJEOUjGHBEucgP9XX8gEYy4bKgqpvy7NLMTteCKWdjHxjakQ9
VjSgM/Yv+9klF3XD6Cb3bVboWda7ZYwSH9279pOkHh0h7TEmxtwS8tzORnkPQA4hhyyD/maFyg+K
43F3KRGB5Iiec+X1g18mqF84+l8J2iHXdgL9uphE2IFu3Tbo1BSdDsMTJyNghL+5u8extqlNJ7So
gko6hboCX8A4FUBJ2wNVEt+yW0qU8QWCOP/xnBW4heeK2MxKyZoF7ofHyB/eLmJv2jLyibfvQAFj
lPLkF6ECpT1uLjf7WbmJX5Puiv2xYMZ6IHLQzf35gKSGxjCofwz0xIsB497mGtrjA+XglE7o68+v
lf4YI+5yHJQrKgzBVM7SH06zIj6AFodOsXGJxbGTk4OIrTP2ZJUl8BwfXMqys0E9m5Tnpeykx/wy
zQdqFyjDt1zYXXZjyNKEUT+jD+XG51a1/DhDDm9lC3ofc9rxmrIrPxlclLDhiKmLFD0Xgo6svMxN
hxgUTNB+DssgTkmF739bi6DcfYAZy/tdp5RvJIQiQNE2YU5Frsmp0jtYsR2+/21Ar6BEbUm9J3q7
KyeK/rhSothz8oikSnNs6iXZSJj97RBmHqBxT5nCEpFt4YrpeXrlambUh6atkG2gwsIf26e5Zy44
MbGIvb0rGJnihvHFCuleAgtO005Rc/dVGhUmRtbgKk2MKTQlvf/Ad3eGyYwdI+N9pUeG23v08oWs
ZVfZ86qpTi4iCdjcMuhubBFzbgOQ5Y501sGxwgj/KXsmD6B/cVqQO6u7DlcqZDQu9n0IRu5P1IsC
tIwzaXuI5KEtVtvWbnUUPsfBVXqfrVHRatoLKCwqnuhOviUbb9aWSXthvDvUXHqlwc166BHMIKQ4
XHS3taX4rdHfmc1X9uOu/uirtVw/JvLOeMjFIefPJQBZK7+ARDHZbPtgpUfq+gdxgM7EjcjBK88f
uCFmH3d/ZtO33CV5+6RvjKL3xqfMKI2cNfJc49wCwSYbWBRvz/m5OrKq0ERnt7vUu9YalD4moEP3
noyya220ckyS93KA3ry5O4TkBYpg0xbJ6iJwkkgVfUXijxnGp+ntrEuQGixDZVT38ksZWFY08DeW
XR5i3ncTVDZ346ov/PXgtsut+RnfXk1CMSgdSjK9GQAMh1036mjSPhLdSJF7JoxEAeWqBgIL+am1
I5cLY0pnc5pnJEWPaOtQqoxNEveehD9Y8OFY9Qi++lfvJqS5z3vu2zcvjPSOW0pND2EiE7QUz8/b
Jnq9sqxDUJdQdb0VXrLIt6SyOatrKMC6juI9t8kyiqzhKGflj9c2sdSst/DXZtxVqFN7NIGlpRAN
ypwXIxPJfL8wgX5RcoCMMv111beHD1Gt7KT4/hYfzuM3W/nIvcZuTZ+JtVf0DTRs/irP0Ean1jyg
Rd+um0XCTLO7B8T4XkET/EewDTEwUgkeyK1B3rdW8HgRvFqFc1bwwpAcu8YPJrXa6IxNoD3JWhHP
A1k0fB0G19+SNH+OF77XJ9lV5Lp29HQ4gZy/IJTm69vl7ZC1jMYLT+z7P1J53baxM86NwWwGPWTm
8MbxGVtvaj2cXlRkirChDrRj59CaK7zD0YlJhaC1CSs1o37SXKeWQ/jaWB+XnxY/FJ57Q5bq8lxK
m/Geq78iFYkAqz/agTO2KBjFuoLa3wLOyELugo91Ed7iNcyxEAbmqRc6UQ5D5LlW7ewO92r52m5H
JwOitjvYdbRYvx98RtZQ7ZeW1hgMlOJvJ5kY/OR6IqRFrToPJqME45dlgA5XOo392QW9cmgtfQ8+
MFvNg7K8+r3EBDK6Kva0ESd9AiHey2TLs9BAkF8JYs02ejWYxsySuUAM9VjGF9GUrEDe1y9rTw0l
Ogs5YPjRz0N7UZnxcPhsOvK21aKxNS8H4IyAY+y/R4qiURUeDlV1m85H/zI2zajV1AfuZquqF2vp
iU0XbtohzQHY8/0pqEA7S2wO95jmd228PcE8cJzWLXbpMH+T5g7vLDgKrp5cB1+l9vn9qsBXOYld
pK6kuAORSsKMwsO0jWFE4yzMb9uG08mZSIMPv0YZJMGXEUuh5PRhmp6slnzR1XSDaglAPhWSvCBe
sVHE31ULwFVPgbGBl3PLSt67gaWyG+MQoRszPl5Gr3zSYi3Tc5mlPelYPlcTj/HNRu7cp+VoSqZR
SAibLsGt/5NQci6sggEQOVkQ646mIRsuNZ3pR5i8oOIeKUTbCK9NVUSm7XpVc/f3iVZOyZd4RP+b
qOFBPLo2qzhuNOTB1nbq+N5bl+K6QaIAUypUySr8SLgbRXh93GFPKkxft7xGXmC66/Yozd/7kKbn
YBRQ09j05iZrm1se1jM6jrLnZHxPnBTysiqF4yagCADOqxA508vbSt2FXIA1Uuce/mu8iy3JV5ci
1tm03y3+Ee91qlwtwTT8h98lyV1jsfa+M7aJFtMb05mIP1b0cpKmRJvvtbSb3yWGspB2hyQLFuNc
SB2eJmDimhbdiy5F4LkmO+ywaT6mBdsP09d/6tO6quU4AD4JfZx4e1iDX+Ih6LJh6LUMrgHQBLyu
sG8BK/aa6+SsjOh/VBAvLoR00z5mCW/rmSrBwN1W3ggD9tHvzmBkM/tbdZ3LUXzmY6pxAerhdzxE
9mWZdCSTla4mm5pho6xV0JGtMgS/XwgcEmm+9k/xmWcmzzhFi6spCGAFxQB2wL/XMgAXpDSOvP/n
Vn3ix8ex/Jc7HMur4Nr/xRxf53LpoGpTZz5rC4IJUVALidZ5x6TEKFgYWdoD06hWa8UsoM6UWgNH
DoAH4H+DWOLb9jrMT0yNyEBKrM8FLwBpQV3X7bkbxOQMUddc+ssUwW4shul3gp+dz/dTnmjqZO60
oWhH7xkJEBF+nLwCSS2sbFWvEh6u+czTuc9c8H0gKsRQwCE4WySIW9q6S3/x5V7JJ03Wds3Vs6nV
wE+bD0tOanuVaXRyPr28NUEdJl8+ElhunhaDYWcy0QaQArb0fKqgZbcBbOzDJJY3xmddn1Dumg0A
95FGSH+iAchkqnuWpYAUu4hz1sK8rHAlEDIJsuN7bydsnddM/uMxqMgxnaclnQ5eR+iNj3z+zhqU
+7PYRgl7DO44JPQrjp2de55hwKhMve6spnClukg4nIm40V8XhRw8RBCSPPf6Zba+Prq3PIFHiJz5
PUnTRNiGXyV1R1vAbJ3FQEUm5MDFE84cTNaUBAgruEuqLuciT5xRYJWn+ughYC/Pd7lbiCyBmlqw
Gpjxw6hsWjgQiFCHe4FHI04JOplMiQvJ5yaVAlIY+QGsY5TBiksd3jopNV2DGCP3kKqWk82MYt25
woyUxRFRU/8xj8jH2PsRY2bOvOMQNrZlLOR9vMbfUec6HFLBq4GnbEkpx9+g6RNBu3Cq4M1z4tbf
zAN9D6kv/CV6KkNfOHXgujeB3/E2yYwwikczPGXf3yLFFD6rG6gZx8VLpwSXbaMkiXo1YEc4n4q1
8sjwXN8Y0f1+atl9B0pK+PgvEk2OqGON3q3hvOLVn02IDttvR8+JKeDv8FQvBwWgKc2GbKYtbciO
5tO7sOcGLFFcf4OdxrLbw2Z5d3QBBVJA/VP6ba866ILRBqCb3xhw2d6I/KUxbR2lan0Zp29CwLeC
Y1a6X0Qemk6X4Rlg82qVQ8478qnxzUXC9ozqAgNIS8STF8dbAeruluE8I0W7WTCjv4zxgI0kqnBl
Dw/q7GwmRrfVH+kLNUUF5WQcdpdV9FDDzWDi7i6ggJ8ukPFLEmR4kZYmYkLV84eJlBDCf8yQmqKK
TZtzXh7HrEvtMSdqUblGOk1CU0YREsvhJvUUrEsyEV8eAjf0oJ5zCwtNypRiJmO4Hb09XDAiTjOZ
W5BsjpBd4tHUfYJiELFAvG4gpq5EZ4gRAsZlSON+nc9qICptFWXRrwgpPfZRnmBfn0Etdo4X0geC
IOvyaScCXrjqq72vDd0ZqYVEaS2C47anoxPrPZ8k/0OsemK3DPrV2Br94ytzscHIRIS1X1yaiMfM
ZmKbHhGyeLLfEioWJlaXs6XoYY0tVEG22flM3HEmeJ3O4nWpXoBTaFh31X9Zw+ZCOSvZlaq4Alx6
5LcIXKTy2RgJdWWQiInZ14jiFGRtaX6UL5Z/pmAKveIOKP0sNFBNiSMPo5B4WtmoZr6bn+Ab5iB2
e8RqIXisu40cYKEmStIHc2YgJmNKeHnQ7ACyfVcJ4ZKPmZIvJ/mPEWI3sTdhBl+5b0pdtqy+/gPf
4gz16V7mkGMlx6vBkX00vNAcVbTM7fTaEPl8or8D7qo+lEJGUJHD4yfkwSi1/3SsykU3u0G75Qrt
Y8VYuy+lsWB04Ip1s0vr9FXLlNOi/O67Utwq6D7Nih7xwmXEFo1neS0kIkb6+ZApqhYxVD/vv9GM
JRQ2Dw3HfEF0231pkbNmF1HEMZlJLXMkzSEy80bCzfQEcSaZfbf0Cc0kB7UhMsHPcVg/NZAsLc5p
Cj6XBwDiKwsCLkynbawKycy8IUnq1Fy6/uPLuNOKzVysc17SMU3sEqLqyhMQTyse8Gb+LT+UOnrZ
THGko6uZXAyWzZLu5dEkTNODGVsqlyJEMYuMyeOW/7NV1KSDqp3MIX6wiHyhchOP0QgGStMUaRyH
izQhUDkVK87TqcelPiNylTyUfWMsV9T73AriCpcKJo+c6cJZ7/YKB/ZtFubDjSFib3uimzsJ5nf8
1BNUY+pif9umNg1Y1Bddjid0zYrIQHwAqHONzYrGOYy6Cu4UsqhJfCl3r5N6wQ2zm5fLkVtpcmui
3RsxCPrSonRl2iHNzqLy1onvoljZmvFWtHhM/eeEBHMTq1854GSvmn1Hc6Hwn77FQDA0GR8kAsWY
wzIDdwfxDAtkISXGy61zZjlO7NEEKPhSIRUdqSyuSZG+Cr/5lZ/DZOTjSFusaC6/BJZfF4R/ZeMl
F1c8IYOzPooJKKzQNycUp581h5CsAdv7I0qxzvgHgSwExoHrhZjMIZbNgQsSnW1kZdY4VitLB/7X
AEfd2Vcvw1StwEKFFnAKjvafpXbIxxkAnzLsQWMmfxOzkywaI2YJl47sCQ9EH9wXnBon5FoGSbie
BsflhXFDd3JOFsDCN5O6Bda3Xdeq7CBJHe1kobz2jViyUDCPNfk42dO04gdCznNBIYPOlJd9KVZp
L68Ca/di6MGO64fSURVd1GnUcmI84EApG/wKo7wgGfdLbrJb36uKmzSAU9TalzwVgCkerWoDPj4U
kRmDYY5uyY2Y2evgolqMmAQwo/I5xYwVkYaE1CHySD+a/kp67kebJRBz33zA46rA36BZD2lFBNcG
89ZSOTagyKM/Lsd/x1ovmGJ8KO3TlSjBt/u2DGHaR3A3g8dukZzincPopDrZVwVl8Qs6y4FfxTQ1
2nj21Y5FiyAaSUpi4eMsKN4Oe0DMrIDJ3kFtK0HaS6uNpm3z6+OdGaFqAKQzG0HEQTXBW4+OfLGh
ZrXk3ovIUH3KkvPu7RE8d0XF4F/LDOSEZ6bSgGjiPQ0HZKdNBfvsw2BblkwgTq8wzxZFhAAFBWXh
Czu95w1HHVUJ46fd9t4AAKJgFCEzv+7y/rhJKxWd2xcq0iODkwW8sb3hhf1Izaapv1sALNcbtyzN
S5M1idNVYfqVXdtnPzuZHomGstKAAmOcQZimCTYm+J7X9rcVnq9+ge1q7rapD11A3W28qVZebXaK
tcgZsOeapAZZyG/WR10zzgVW3i/X09QbYbDMSAv2O53uForPa4rwcmANjUrTOuuX089xdFjC5vPz
RFXD1MCjy2OBOZL6vreWUuZ39QdqLwlmzzh0SB8lvk8ZOp0a1S1ejNKa+88qHp49rm29pZ4WAiXK
YqxWg3JZzkt2xiyx+GrjRRm3xNBXJEDFUu4zfESbOZzWJwkCdU/Niey3/VMb+6QGCiR6ksoGTfuu
dA349hDQy0VCmaYbVUZQHFvjhf4gLp/0WEiuVmqCRkmO3/pXIHblzv5hEdE0tS6xWNYCWOmF4TQQ
fpdZviaRg+aYeMjfdlLIxgYyhpqYUIyzN9ejyqyPyVgLb9whbhw08ORID4JXp7WLDR5kZtfIYdo9
a9cXzn8zMNe7jjSl3Em61IJgClfZDqqYuv9i3at8T1viuuRhaac46rc4Xa7yEjvHaI3UdzQURZFD
zF0CdThtF66jfrotfS3mDGHkzKwo9wY2vqq7ygOddf+QKrSZ7kyvGWza1+3bJ1L1C/nEChvCtqFs
ROKOszQaxRNrQFTLzDZiIsJuCkTuY8vSwMMyX9O1SeTdGqIsBi1Zta44TEVojdgrsnzrA3Sif6og
apfZswoUR44k8WlVYXjG8PzCS00Y3DR2sHtEUaVrLnHzphXo3+eZZRsc4SzdHxbyNox+5K8fNec0
gk9nvAOC4bNHMV0kBFRDImvdFomw6JGGZTRkJfExXmcZ57jB8GhTpvN/X8qsnEnhls2yEk0SxcE4
Q2r4sPGbPLcqN3j6aKM9z/+9t2nhxH0LxFKeAWL2Z/iMVcEHPrNNhSnUe9w7Kk7RvzUzcf0T4YaB
9YmpHdwSTEsbheOsfC20OAIyufgifi3rWJ0a4rfcYYs5VSiSK7IhHDIUxzRzeBPCy/kOAdX87Iq3
yYQI8amwla50rOFbtE7zibcHkiYprSg1qrd5Ub9+ck0Sfh+BCFmYVMJ6iqferVFmDObwGG7sUdKu
dJBZFUNkkc4AaXx5aNofrM4jo3pigife6T1E65aNCVFI+5kzO+MDaMmOXI7ndwpamWQ/Rf4zOiQk
kaKwkZsXfOHm94MzDLpZ9t3WXYEGiLDpIKpIwTfA2omtY4L/PWfMzP9VYUdZC6bGLqGXVy3uTr/M
kwnr5diyvDzI5b26tj0gdJR9f8FkA5uF/FMwoNBf8pXPEhpJFwRJbYSDLuzfOZAgp6n9sd8hIKXS
ggJHzqCJI8gVtjWpXJS2u8KVUJpWhPpn51KlRafA68cxSlPHMbp/sn7l0FidEIEoMM2Lz6h1tmky
rgWHl0BRLtNcrVXaKm+ehGCDrY/A1Ootu1tovzmBqI1SM9+1nYFi4iowQSepc3rPGy4FIub6fe+E
WWHwLUmCw+N3YJFHjDrC4EljGa6w918zQWSlduUAHF1cgQMns9l0G3oKASB6pMoEk4Q7cBpDZH3s
aKU2ICMnjErRRCGOhN3r00ct/Q50Lmdssdc1tV+vOmGNQOU2Lo7wCwcoaR57kJBjPgDdAh4VKkK+
G7KGIt0S61ZpEma4emyhfx+3l1qMzN6gu7zvF2weOznnN8U0tO3fHRtCZfr8gpukUAGyfKT0xoex
Mb14F0tCa51+CUxvYnKchwa8uvw5ifXEUU+cpYkbe+8syMkmIoFM84VTALnCHIR2yeguxHqbl4Fi
Jsu5JaMRv87uqHi/UXfEp/+SH6KTgmxNxCT6xHvJx+7U8TyiYq7Gp56QVU4lJE1WzTsBhzF8EQx6
6UaPCU422TLsFdpWUNbjNrQCDydBHif/eF8nM01AEaLgjuYXRgBXIdZLoyKg/gUx4EKP3iXQlo37
51s0hlhUgEU/oF3mYLWV4GEDWJ7+bNo4MgDF4MSWBWUIqAkupxtD/Y3r5mkTpPM3dosLSCKB+TTm
Pam7/MlbhU2cIQ0p0leZQsw2/3/nDLCwCzzlRFKQZKaRrSWEtcjUa7FFrvJeeT0TmQahVVrDT6GC
17ig/joRHybatB2dw7RsOhiia/KrW5DS+d+AuR7NQUxuRqSnKU9x3W177nJednSfvlifcDaCe0Ti
RqRQGpC1XFpB1Bb3vw4lYQLZQki9fA197DgQ5SXGkb0HptKFLUa2WXI1h+kHTdgYJ93WZ9w8sVir
5LrEAbnLgNKcfxrujI+xoSo3Q4NOpDpLyMVIiZF7JnO+PWuS0mPrLxZmdmiUCm3b8mkEi+6IhQvd
xbtGLCunDBkprYQizVkAbv29IU7ZeeF0dcN0Ef6124UACntuRN5iKwvMIGZJFGxNRQUNeMEFHciF
QNNCFK/ntermzRqSATuVCMeOcfhrkGzQTkSSOKvvY1XGE1K1cDiqEpLqsDG3JI30nr9xaP5/6iSC
9k2bJwm6VN2oH4f1gy9BRVFM5o1XHFqS6Jxczr0PcMQX77OXSdcSMNT8xBNem1lsyhYx8RoEtJ67
F5IKRYUr5H+S7s16q5zABvhYHXSxR8ND7YAFV7S6CfCBC8gJXDLs0oLKbh5/EF6nrj4d1J6D2Qip
asCpm8/08d2JgxP1rtBxwunujtsB7jTUVWXOga1mIbq7pcIluK+YnkeOvLPfgCLBODQfTf509y+q
Mz7IHTL5GxmlLz58C4oTUEaOzgfJ0dNwiB3BVsQkchBqtyLjXtpY0MDqI2GqvtOcfBPrD3YnHTWv
eJMt5gWK4VzXxoCKwPfM9gk7SWpw1LMsyHTwc+lg1sz01AIYjgqAMaFS2UZnY9Snnc2xeNxKII4Q
/Nbj4ndWN6rWbuG4WbRTUMp6M+Q1z3bWDiLpp/OcKmIgZOIkfH3ytZozUYXjnUsjxoGUs2sNUW0z
JCX72jQwbjgjzqxTa7XN9T7s1n5+fOfqk7VqiMqkvQriVgj5uep3SBiBerY6Bxj3wug4k6ynjyPF
cuzs8D/vdjui9OcTqkWLkuhQEzQpssWgrVih/gmae9k4DrYV5AT7A2VbkJpNi8rFrgM3aH0DwL53
yHxGxBzNJz+eOV9mkqfmz/1fO+mqLC9Rhi6kHp5s4bvE6zg+smLlVtJxBfPqbZklXwvbfHYqPkx+
C+++HwJNSCItlpPDK7IyzJdr+6JHFI2TjOzZPf8DccRQ+U1cdftTcDfjwV+hl6Gg/rEldhb+8FN6
ZViIi49T7OO7xpxquFCYb6LUakAMzDmozKi+u8H7qjIJeKW5Efgx4rOfucekyVmN68ViKB2hAULW
8Nx1GKL/WDfVQJgYHhj4IhK3SiaWMDV54eBd4o8UR0HtppvGPbNovbK/Lec2tkjjM5CpeWU42BfA
YP4JcZW4Pjm7diJr77VunamYcz//8mLFP7fH/22rEhqPrwZwu/4CsFJvaqF9t94sIoihVSQSZpE+
Vo31C552VGQu0l0ErWmUejlRJS/mRQAug2AUSTOZMzx+LmlPOv07mHBLB2MNLiR1YnfwFtXHt5ZM
IuqFEHn4Pz8u3sALiTyvf+T7QcqCA5Q3reMoF2y0V8ESZvtPbLGfyMRjAWO4Kb/ManxeHxw8sPIA
vUfNUTP0PAgIZAhQpM7OuxLVrytRZJchD//+EUDxEch8cSjjD3hA4AuX8X3MUOaARiBuzooduawB
r4M8Hv83zU1aQ9MaYGTWl5g5rBlA0xahaVOsAFW9ZI6T/OGqRIokEc8ammLhPSoDJeiAyes6RtqY
wxzzdU/VWCXmBgYpi1jJNpMzTHM6TaRtXFN5eR9tu6erSlPA9ooHbH4CCiYm8cBZF9nNnre6SmC5
OLkiBjuP0YsapM+9XKl2LL5yWiMGBaMGNNdMtPoKPcGxq+t5C4/FX64ima0MbQE/9MMbdLKlVjMK
ua3/XbZXEA2N4641d1g4CAjJ1y1kFlkk87emZcT34mbyeXiRWrZzyAOvgfbJW6n01T9DXF3iulFM
u83uAzwKQ89AnXTz2Mq7KIKpQqrbUHbNGHaGoUQdTbi9OmBCOfWyi595pLuAb4f1tDTJv9rwQFxS
Wb5xFa5KQbkmnEYMV3HfZEWrLNB9vKyaZYLodQer+JbxS7icIUQ8EsHUk7XYPs+QEsrafBCx0uzO
geIlDrGxrAusABCHxmkK+TY9LoyiJzgr6pKh4R8lHNSU8nFlpGxeeJzgNcuu4TwI4pSg7JehxgYJ
QftADw3Dm8Ff3lasb2dfFKBzpHVck74uGgO6nNU349PUxTdwG+3StNjG4uTgzTSjnPciBTB0r7n0
AokqVBhwyWGAwIO+7QlQRUAiC01w1nqRJ2Qoo38+wf9use9ItCp2AKQPsF3ZH4Rdtte+oC6QhIB5
lBI2JOBRWIj9fwvvTp/bnUcgQmEBqBFyPx8SQP/LoyAFfpENgfdgk1KVNvcb/xV/cH39USWOkWY2
J3WNllZIMhTTJFs6P2aSqo05mWbAVHlEm2sQbozcabN0Le/gY/QNQkBRmDzWdAg1K4h9WVjnSN/e
GEst5PLB7/0wUUm8tQIMz6pAvFHf5XS/UasGNCYY8N4IoBG9fa2LOs4c0F2Bt+z+3brpBMuLhFfi
rpZwWvTaCCA9dsTywVxKPkALay/W1i4vX8hmjHnw4QtTkxpyo473cidYEGL8hCsgBM4NPLfoLuQR
5HNvhrdTnh18H3TWpFnMXPmkl4bnrVN4L8o+49p8VRxTw1fOTOlUy2+ohDDqnTCFeL5RQ4OKkH8I
uqeNGXwpi5ffQ/bqYNNCs6dxpP0qy5XdCFLLdfQah7Etw34CI8m3Xb6dcEHTouUkINzLc88I2XVV
wNeiksFs5ayZrKjvYcfFJaFp+KWSE7Yack4OQVwCWk8DeatfdCjKlnwy/1CfKiQw4smNV3DS73VT
u9W+KDko7fpUZUvQsgGmql5sNgFQsUjzUb0dhkW45WiR8PWfuhHj9V/LV71cH2a7kwZFh68BwQYc
RyUu8mevE7RWslCbB4DBq3z6eR3jXB29Ng+aKgoCqaEu/L5hD2PoKFwWGN73O6TmyGfyFacMcsXA
VQPkqLYGgLbI/po1rYN3YVMgwc8mFUjpghniOh3Yaf9fyv19zvm6y09/9vp/gPhhzDR1lhyaX+W6
05iqFrjLncwuRF2G0RQEQ4O8zw879OVpDq9xfk8rq2EPQxebDXN+KNkjMT8rv8Gk00JR73emzBaZ
2Z3KhmAWlTbm1bp185eBCdXBCDQ7b6aIVvWLHvxFvQfEc27cWa0WofQs7t5Bd7gdA1B0KSz1JF/U
J1aksdf/cUZr99tujAu0QR3zDgZYOR8tKEBd5j5T8XtxKelMsXo2u7VKXryR00hsi9p+RavKeqSu
WjYggev+5d+N+pmXjicxGuuaSXumIdEOL/IWWZ43aK4c4uB1iTsLHm8d+CbgJUT1Ii66UIRF7vdu
pfh5z9fG+PWP/vkHpbfpkCqLKUZkPiW3sKiM5jIqEjtnPdSjF9qtNmyGO2HP1h+BKUhIVnHOAxhV
REYdEeWjYMsPYOZ4IgGvC9AGdA76XTomvN6z8QT3w5wL5djBh4nWCF63RAEt3MX5OuJNp4WbKNKO
ARISpxsc6X8sMqbgiSIphUPKRvK8hz31uhtfPy35uOO7GKT8CEnEJuv+n8dY0+R5/ARcFPc48KPU
qxwAIQvEGhtb6gfDwQxt431etgfptN/2GBX+4s/IxsW0zxwDvsqTWQ5zlAtgo9NG1zr2TkQTsJzv
L6Z7DRMLtu6atzr6L/yvMY4nNp1cSm2RLv9i1pKLJV1dbxO52pMXK6sXEMjhWv1GgPUy5vr/dKv1
o3M/CVFn7sXOUtkfeyvpuGm6E7l7GM0lw2kQA2jrMqkzNbGfxoV4Mipgv187ahskhp1EQbnXJpsf
IC4imncT2URNpWFgbzlasHiXS2FgSaSNAolfcyBMmQ7Dcw+96Z14cqLJmIthvOgBLqRq2g0Bqlco
dh8EbvLYeWhxu9KUPJy1FvMbGnPY95rPKT5XqW4K8dBaD5vGjSBTxBjbdj+0mgwLab0BhJckh1c9
RCpdpILkNPNHXflq9N6xN88O5+aDEW7FDTbkB2SB6HzjzwgKZQgNHoVI6J6Yph268v5jqA+8NW9T
IkAtt5k5jdErsKJvvj2fVrAwmwjFg7/UFaLZbmqJ7E54WIco2CP7oY8qNJyAWAY3UkHolUJMGcdu
Wo8j4XTx3A/1qh7hKk1NzeRBvJUP5zZHFrBKu7QAaRmeH4HsFGI2ppkOT9zUQ6HylYaMoYCvfINZ
F+EYfeinHfFH58f9qc4OTb6qK5FDdyTKOJtiK9QnR8sic9D8CGCiA22BjHBcnEr2yLKEcjxFeC3l
zxAfPWnzlHXZGXN+Z/8QSmZUVpqppEtuAXf0Ec5Hb6ulw5lI2cnEGU/A5FvikE5q1t709geX/Pbi
uJ20zsQLNTmKABe+bHeTOgyKV5zFi9XEjkVhl/ifZ1+2Ao/BJAbj2puRPmV5ze6SzjDHzbG339gp
dQLrnYgdRXn2eM4ejySfqSHFVovzz6acRXEbOfD9jR2uN4jApHumgFdxOSRDc97tmfK+Bif9v93o
bDGHCC5Krbbh0N49/hpJP8cLYzskz5bm+BML7IAHNTRJne6cE0YmDLZyoYHi3RPy/9irQJ66CyBo
NvqZdLDKSXCJ4VOmpyWsxdkAg+2OZemWeK5dwi61TD5zHG0E6OgZiP3hf5ZRvGMbES+lYEzIdKt1
1cnn2uFz5PuAUPv/kvNwgNGsN/Yz5fsu3/NsCpXgg2Z2FHFyojkUXAc17ziOU8rFPv+RuBBCg7aN
ozK5r223/sz/ebnudw0jSiS7g6ObKZMt6EMsEcOqTrmBRg4IGc5OKiufHwZqwqAvwiRvje1mu01M
oUqV6G7YIM2klnVX5CjXz8f+zXBJpclVkklRRGK0fXMHLE4ZrGho9nyB/yEEr4cIvMv8Rct3GUDY
Aal9XwO965sH4XweraocPHMHlgG00JCUOTpgThR/iSODrOGoWhX0jycFF86HQ8+YjUDNc/Cm2cKE
1rcYDmMC6yzqxf3Vp7fQ6J4HU6FyRG9eRwrnFQGZaSB9Htn4ZZ6t11p/5FoidBh54wV9Ega0d6dO
Ss1L8XDUy5bNiF8ltMAkDgg71k9wuN8Bl9qm3MYvqiemKzlxxx81LoPegFj/5zViNQtiKLMlzzkq
KOjub7fpLdS+peeQw41Kb8XEbgCffocZQ3V1wQ876YrqvsArmbbQUf6ncLRkRVzc3l3E0tu1D8fG
+pzVLFHgGvTlHbHCjc4cnCFyYJSwzKApMKTNJHgbK/HKq4ydpkKOViNt0raVfj1BrdKr4Q0+4pmQ
p9BapYpunUF3W3Url60xqwx/H2VMcwi13e1YS+EfK+9d8aSBgZUphWbK1BWY7TNQFA48Q8oN2L+U
NUAK2RP+ExIWNK/UUiund4P+mUS6+7FOiXBWI6RgjUbTho4KwT3w06B9cIHku227Zo+FDoD9rY0S
E4xqdgrKfafgnytrMPEJFTEaIzoHGpgD1jeryTajC5bAFebM5NRcxL5QYVDeQzfEsxGSzNSS0HY0
K3TX6FYu0LsMB9VOIOkl2bgnutZ49TnCTDPcCa2j6E3H9e80nA35dIZ/bUlmkf0EeTgenxWws4PN
mU8aH68p6lYrj4anR8kUCaJuRfm7uZY13Sydm9tB8jVQv80B27f0Q/z8Iufl6T3B0kHmps+dxZBX
rk/W8/pBwaCUtfq4Dy2MdE7lvhQ0v43fqm6ItL5JQTvvi6sQypjjIYaDQ4HWM/gKGhzQKoiP2w9t
xMmHBm9l07PA8Bw9Dj07BmfhLUbcNLDFZ7hwpLdIiCMm39FDRiawH5kqFdspI0UrxXB7E2AGhLtO
RJ7qfLZ2eohQMAz5UHpiwJ8fFtQrBmk+96SpwSMJQBjHpSJKuwTduhe1gPFkQhPrEMW3bzyq8mDe
FID7gXw1YDQexVoRP8FHMuacFd4VhtGZSW1ZMCJiQMy/OCNvo9PUUc9titjjGjWuiQ3ksg62ThaJ
kBjaLblox6QScgk5P29+NLqtmnZKDqjcHs41v1QdQuDf1D5t3aWCZzQ0YuEyLdQ/sEfD7klEYnz6
AOFX7/lZ+mz4G8Xf7XLrbMZvERhb7PkPTYjJPMXLy/KSdvF82cupw4tEilhGU6BIXPZfjPA6/KWA
hIEz7pvXnqrbgDWiGKMN8ez7LEb+Jxi/z84eq8cICEPpl0OOsKai3ID8LFsrnC7+ieTVCo4ggoYf
qAHGVATcAKv8kLPpnwGWrYYZCyRMojqNJB9kJIF++kLEZzsATMFGzUF0xQRz7MTwuYp/cV8NdSc3
UQWuLxToGKRBZzwclhtqgON1S48gjKj/+tjYUnn27gA9AULaKEETi53028ekqY4zCOQmKERPXCdN
WP+6B1lJsaVc3DsRHZeEYEKRPKF1TWTRno9uv4ZC7yGmHVmwwBZQMPMzrCY/NSG7QkiWkqlE/qU6
fKFTDRPNddO8tDWXRwL437Se8t+PcY5hpN+JcVtbNmWr+EwWzf7Gid2tknKi7VdpCm6O6bcaHso2
HCPfqQPSjQxl54EsclKUg+Y4ZL6Cil+InnRpJnw8CPdxt25W0qmRJqvM8B2irgT45KrFTilszdF3
ih45cA6hMh+CTM+44jP9KDi2nQ0AivvYUTl9sUj7KF+sSGx4TWNJroq+j7aTZ0iDiSVBaNJJNF5X
feOa+2/WU1FuykfwKY5VT0PE+vXbqINabuMRpbuIZ9Si3J1tdEV1jOAfXjZGTcnYRPeYOVlyidbp
ANwmQn7QClPGBLnqIs/hC07GoCQH4poaXtloN5FFjFxF39nFwMnyiXpXFFUdbPypMvZYbnE0JYnm
rxlHPozOTnEm8juSqIwrC02+4p3CX2fWDOIFFnIBt+FfBj438YZlSG6+hdRGD6IsZun1v8bXlL4l
9C7wVylgsmq+rq6WvrCr5gZMoNJRcaDChQnnFvSmZAkE+p11lA+gyqhrHMRy66hLPzP1XICrdybG
KPlOA9CYWmR198UPpb/zzUbD0Fr3cigRqonaZbcWb0BJppuxx91tijXFUSlnGXy8y/qNPjF9+TvL
rXo8+H3t3spDHxpSetyjKkBSbmkmkwsfCRNIqcg2lizB/wDQK3VPM4pQPjb6SRQAIQCd46/k2JaP
9Guii8YgVk+kvj2n820b/7BDcC2LnZkcD1VtLFgrTMZb8P5wdfJeUKj8qdXmgnlA4Gu3b8rFNzDg
dQIS4IA8na8ps7JrMqPLOoxzvl45zPFMS+BqFmIyCErlDpU4jOZ/UvAwb+rq5yZcimGGdN+2guhR
tJQQrT8rbNHNGBsLnvt6/EElhFQH1IscgNNt8cXQD1uTsE2+0S3wsIdkIeAmv+T91o0Ww6NJXD1a
FlL3M8uyl4RSjtNcmNiwmgHZfhv+ad7WWLxhWMrpNkBbRtPsnMZJuliaNdFO0PbL7OZDk7soZLoR
DbnyLchwABOqtafBqGJbTfZvjlx6qFn6Rq1zq9nNRetzSCou82WXIJm/T8AEpeCykU6F31GR+njm
UXRtbh1nE5zzyGgCm5pdU3GVdq16ykYB5zimMRkSVxYWsPCEvIUSFDnim8F86ZiwiuU1RPZT2sQu
pT7NjF9unWRC3fJPfO5bfKCDnGCG1DmoRWxHi9P7tqSNkHxrOhAYL48jEJGxHQxiRkqTrlJz9qgK
4lyKahggDf+BWdLgjb1RccrFLv6zi2PbyJo4zFNoY+SmVv9Mzq2/iN4CGyPfmIVCsQKiPfQ6m2k6
xElQvVh/z6WIg5kXLF+dkrlS8We2SNcYAuf3xUQcWZ/TWfASLWCvZZGdgZ+soCsUSo2J34A+/QNm
eLpFW8BwVk88mSamf1QqIVm4L7esbNxcVjSt6b8W01Lz7yXuyc7CVf5mZAn4S1nn7ZNZB/XQQDrx
xHC6s9KHAWXb1nPYvRaNk8mOh6/E+uL+TYp830IVqoflphiwL6ZJ0FNb4LdLFQa2XWEIBYbRJLF1
zWvrWWMW2ZMp+tQ5dnY0ygZNIlEGfIBjgsPP0QPIidhOb3Mfeh3PovAW/Ati/+eg82FG6A8KgdTl
mZz7AKu1Tcwjht1l2KhVoxlra8eIHvzMPL97Jipu32CPibqjjeP9qOePjAGhKuxytctMt3XgXJuR
AuT0g3L/Q1P2s7XOJW8qye/OMChVwqQXEjSbfsTxSr8vUfbAEgnOMMYk6VVaIUGGSAp03FX9cmVD
NhEJlhPujRfY2L03rYgUApyAwArDjqLO3pvtYgulBNIvUSA1WNTpmhVckQkgWoBRzW9NppVb/Xax
OVvtCe1tJFqnsoeAU+UtqIb3uxetPKv4d1RBRc7+kWX3Oxjf8QNYdbftOtZ6krDGT7wD5OCiZKbd
/o8vUr/k+q3c02JgaLj3E1k6ExQlS62ItbER2DbhH1VE93yq7SN7NyN8E9EwPc1Cq3ti5FCkjNEf
jmtZpS787/SFpkCjvgrUv7LK67tcVT1Aiti8Vxkt5u/1K2iZdbRQHaDjDmBzL6ufrNVsVw+aKR0s
WyLCClS0Fx9odpojN6l3HCrns5kT8MbXfYt/+z5ogz9UvheSV2HgRaajdoCrUqcJrcPHyQfJTSbZ
rB6Galg9hKrCFmlwtvO24miCKiObrps/ovUBE+sui+Exv7rIZAoO7qjFfO9GkNUz5eMjPlp9kNpI
3VhHtJnY2u/P5p1CS8ywQdqqOX42vNIkSxFcrqxCW8IDAVAHW94gOYKQEyolnk6r/8CuOb1QuzeU
i6MvkaJBJcxNe4VHmDo+XUYXEaI2k4Pxn3LRi8E3Frfd+XawIbRjJCftLtunkZ0GofcgdyftSLq9
TFw1brluMRefe+WWnz7YzGgh6k0pohN8bVxYgIY31gDayGLQXjPDjYZX61Pwje/cnj6mPv4ZRiNg
mp5vgYw+BunojKDDC1OacLKvhrwBdMhL/PxNXhENdUt8QmoEKBm665gK2NmW8VsQUaPnOOG/IT6R
aWu8LywcyMzvEMKPEbSpf9xu8loryBqFWtWekp2Nqnrlp/Ffxsk0r69yaSl3/nZHP6SceGeKWfrK
7Afl0/330YLBA6v5Vb5+PMHZt/rtwjzY/ZocJL5RdakEsaq1PlXeKHDOEFok6eZqCSffxMJSc233
CDYvVnrtZkPoS2WGPT9d5icD4i/nuU0piJXeyGNMdps//5GfmLyJmv6Oz92e9LBrSBM3uMq42ElE
MHcXokgJUbK/3nAmd0+RJ+PPga16AxYnFqkem1UMy9KIDaUCCOrvRsklLt/29TJHRcWSv8c+HqFZ
HLUm/ugmw24pOxTMpqeJ099zVzj34NGyTdX/O07tdqFPWdFXSpwRRG4Gy+gKuOzkD6SYh1+HuyKB
U/CnBt7YjWZExvbxbyrszr/fYZj195y7jHgz5C2HKULQdSpdAa2G+WZHhOD3dUN3A4GfckXx297y
sYUNUGGSV8jRUeSUyJt4av7G/IzoHFpHx0ZPBhzklqih6yi5w6dWZ4F4D8mmakLMnUOk9YxOkAgu
fzyaFH8csV38N+IC9Bn8b9fL2zS5AQcQWpLOk5VbPY9ZgVGn9vAPBiR4oROZvHKf4YaECjPOCRIi
c2R6QjCJDbBb5S512x9SPO9Qx1PpLF2Kvf2uy7bVgEq7bWsdz/FX5wvm5YHSlqOWxg1R0BTBmz4S
p7+CTVXQ/9UoSCK1J352H2ZjBaCk+Ki7gEMoD7h+G2lNUY+WFdVHGmVhUIdee2SckxVO1jf23bjy
K69yQrRnQt3DR/pff9P0ppwPv0MVZSnKSTTYJskq1x8+B0hQ9aqPqdD6YKcLu2t3X6pdW2uz4UcL
CYsLjcoCQrijXCCC2pT51NK/hM+Vszz4FIGueQU7o2kRTane/ru+CM+nJ//X7q773Msjjaq/JQOA
NrYGKXs7+CiKdR2Kxc/M2iOhN9MvwitebyoYwI6+c2AxaDlM/HWjTd173k6d5H+BCz79aCJqfyHI
egARvIvmAoR+vkpAY0nCCBNj5KnY79Fos00Q/aqiK86UF4qGbVEtzFcDmJ5I1a3ogUneO2gJp+1+
870fN62KQMGg/65wQu5tcASSJzCkC2A/8bIf+cFDAKBcmB0gFqC4d9K6PsTdH8NB8I6u9VnWYEnv
t/lRIyW3NqK9RGiiXojLTkEq9Ggq0QS7O95vuaoKQDCflFGY+21QT17YwUNdtbCjaOYO/73kzBez
16XKT01TDB69o10vaEsvlXxBccUlckA7CWcKPgnk0tX7kANiUvpT41vHESAOc2R5sAxlOYV5ZPmK
VFUVbvGs4BrLwfcAeDpzckk5vyyhhghcVoHAEjZlxvKf29ozp9gTJ1SgjfN+0nONwUxSJ2Iot/dZ
RQy8GwpL+2edkW+KWtpECuDSNGEn9e4o3ALAFFxJmGPukfrAnRTilLZv0GjlkOzxi97OuisUNglJ
e41B8WZSgLSXe3PWkl0FGSUWxeVgmhsMPvE9tZOE/9xFrQmA2r5TRvfv3n1G/qZ2nblnWvYWD0qN
CtuHv3sCFuKPERhKvEPbLnzZZ9IIt5Z2ypniSktgMSrZdB0/vQ8FrXYDIPF3Pn7vz2+2d2pCRCWQ
cWQDwjhd2pBTSmK9EoUBkrgl1JiVEf0G9hMXnSOF06Aoo2CZWo7Cn+cRQLEPDsizyxgf/BESewJG
o89ecG3pSOfTBlj2I6q1p6TH6t94ccuAbewckYvbYuer3LHgtXdG26tUzF5FpVcJs7VFRkYycvrn
KuPKcfBd9xToCciG9S3+haOyKAtiD8DQVGNtToyuTFNrwcZdPjZNI79/w16EKqupJr66DomIkG7P
aY5lIgEneE5SmRT/KsUY9muNMDrZUZHHvDkkVZWUScNUGvLpb3wOfITeW6AEkOo7/Ds4Ka3uhLQY
PJID9iB60Ws+b17mnwj3X02ivSacku1FKtFzP8x2fGoupqLT95bOLIEyE3MN6G2SKRZ/7jZb/f1A
O3Z3U/F+++RCPQZfCdVYnsWuxavGM7TT5XrGCRON9fcwIwIDKkC2DO2r1/Vj9iCzvnVgtCBVvHS1
WyE549XV0XC38MOG0USriyRUco7L2mxB9QdQA0R+TkcwqnY9vI91ETaWSrFfHHuuO5BIBgOsk05C
RW2+BsxH1uQaDAqNRdX24tRHuql74KzzyomtYLFrtjZNaQpLhs7wSem7M+7aiyZFH+lbUMahVYGu
nSxb3fNOAV+CROmZpesmE1leZAWcfp9NJZUHLez6GNNSPMobXekprhns3z4iGbG3vvhyxHJVxXiJ
ebsFj+Cr/UFde3iaphhXlXyDRP7aImBCwSUbYvRJfzPqEQazGJqWSBMfSG00cwhaHO4mJCIMlpCV
2q+4nvJ2wa+zFwhhjKanQK+SmNlFxXdoAd7hMXNGArn4JJk/YMC/XPog6jaxLVN2XnPl7qzAIDzz
jwqCnyxXBGWkZZObW6kPGur31Pa8Zce3hBjbVUP2RiSfuJrIZjJouYL1TSGbK0kZcE3f1LEGgET1
4FaeNQAQ8EYe+8LKqei87Q5eLydPsfbx6SsEjqeRWEDkE2Z0g/Vqw/B1CA4FxkmiDJQbLqiHA0jz
gzdHX63gS4Aow6KgNkQxY8uH6KU250Js1urqoKZ70g8atrl/KZkHNCiAzwznIRIubD3CRv/1fZsg
KtveioK5R7AHhe0qWZBO1e34+aCLUf1lB1jfsO6k561POgR3EE0b1b0l+zJU+WfYweGD43cFT/1p
sjE7hyWMqneKWLMZvDI+4JU2ip1USfCxDcs9ucel0WOkbgHyk6ESUMWoOMATO7Mlegx+APkyExcB
bVrE1191VOn7i1dthiPegoqEhg4wOiBw2UOkGmiKC9iA4wAw3ekQ2DuuLhWVIVu7oDZTfaFqEtDi
F1NSApRxGq6d8u06S0rFwsPteZYJfKGfyQBeT4zooH3HoyHgkywE7nKU42gkLVtaDpyNTUZwr9UL
XGV7Jsrp9xXtGdbhcQRv1lH1py119IYEA6+ivJhEPeKdVVLZGW4ebhop0fNIM7R7qGvxJ/3WGV4F
SQQ2kX9sybwUTrt+2lVfTQSBwb6crYpuKatfV2cwK9y8MQ2VvavYweEhIxpeAqz/jyW12KVEwDB4
4lIXpzmMNFM+YKgpCtGANHw6hZl+FYaCPP2O2xFzmVf1EcOBYg2ISNf2a9mC1BpCcj+eaUQdAeJZ
c/aWN9noJsD8SXmreUM0zgKp1UsJC7N4fb3W/cD3OJMVwKeSLoEhbZwWPDFzb8op3b01fXS65+VY
P878Gm88ynA+S3LLqXf+xDc/XGpZdzlL/a107xROts5jiD7KtylzfuPBTffR0dRog7x86PnA2JaM
Ppgl9UwChy5ANLjf4eoRvqCUop0zrLxoblLJloOdkvxd1yKkipwtj4dVB7JreHMiP3Mb8WJoAX71
+tqf4RPkI2GCmGFm0DmMQfylTKyMdSATR3aclqQHZHZ0jtGY4+FmLUMQWcNq/B0R3igPK31ZAOND
Wq6nEYHcvVHaS1vLmCAV1a+HooJmiRkGmmzgy8Us3i1tocUEWNmEKHd2ATG7aHwOpvdP1gETrXxE
4Yz/GAEAPyuwrTaTN6F5BfZqvWp5V4uL7sX1x80VM9wZiRQVGSaytoit0c3j43yX0VhxMGKCzV6Z
Cw3GGOy8glrMLE7YscxpKRT3UMrh+CXd0BSnHUqWymaf/zi2w/zaCCgosQw7k7KhubSIMfdKb+eL
8y6eN1XUHdEBhJLGsCUNOeCn9V/JBtGzpJLihlfDCcz4i7lp6w6E5rldy3xNBPXyHUj1swVIt1LN
ov2yqEyEAha2+y1/9/HIocCW+z05hCNxeNqWyBMWYLL0Jxm7Lm5vfNco1rBc1+x9ZWtJcW3VEHaR
GU6XFq3panSbdM2CAw6B9lzxsUUUYMfJKpcfpA6ZQC5RvdkMoYffQNs8cO2lwc6BwdOnRTT3+gW8
KA56j8zxa0sxNLWieKJPhuGCArCM1w1/qFmeiCPzK03EtgZle35tyL4ojmVjoatbd0Lu8hUl1aA7
agPET0T0tRGtYpXXJ4fw2uHIg/C0Ly4eEaFaR4Zru56g3MioUXyIfd9HPuHnBlR+apIhwjZcIWaK
5V4gMLSLE311XFTavR/Wl4NeN23lIeAlTMo0gbtTUs5AIhc0SXXMaQEqCV8JTOdKfs0EYhnSSzch
3Cy++Etmw2FQtnN6nAqyYeksII9EkRGZBwXOZ8+KwMHXe8md5ZH8Wad0OuSZBTB2E3mhFZOqAiGo
WMrj8eRDnXk95uyMlVHzj9ScF7Tv/3k9/S/X4RIKW4kObjgwDekBqwebLi04Od8hDsIGqNr71PXD
vl+x6hGfBv6omL4HywBcycM6bkSpx4jD5G3uj1t9LUnQk2kHeBZLCE3cJt8myAjYyFLz3z8ML2XB
IrQdxDu5RnZfmmF/0Gw1v9IxG+HeQ/Nw0jeceQzyfDZzlarNeaSda1mMjYULhE3dk5nYPHqdzIrL
1rk/nKiajeZGa+fK8KZ9RI2yiMVPOISs6dF42n8Ma+sFxX7DUDccX8Y4VmemAO9z+4n4OF9Jkz2d
dpazVw8WNmW0kwWwUKMqWDNZ8geoq1xxRMrlkFOXP02S9CCv63lJBIiy7OBWo0GMk+qiGwduGH7c
vDhJr42qcEbOYr+gp2ZxrcPujouga5Z9cO0bTytmrOqm6F99NHRmYY3Om5K1zzrdjeb/vcLXfMhe
cPOvg+6QMVR49Ez39HE3iTjGP2F6V+gjyBH5k6wYCoX/D4uqRUi8iXvXMk1jHjTpecLyWP0V/1Am
Ay430jufh7pWdK1zPqvtA6KkUFNuwjQvkBoHEjTZr1ITtneK4hi1W1YKUiiIHbTrx4rMeiqXqw9K
KeqYPVUg2QfDOGIjUUB0FNX11eYWXBB8cxLATTz8fLXwlNQLNvgmwQGidQmJSmg8i8Ds+ABYIZkK
TXjmydjVjxdQf8+C5W6bKS7CueJuGiaYGib02qY2cZuJtItO3m6VbqTOTnWZSW8M7Adl+HeCo3uH
jYEVdysI6IS+xhiFY7yFxOlaiH7fIbdtCFnSOE1u85dQvYnZnL9+q7i4EGcwss8U4865yFHR2nzK
/gwkHONlcknNV0Gx3Lut6+tINoOJjC8I0DXkGtDoI+YMnQeRvR6I0dx3xVjSxUYk+D7TQ8TVNL9y
xqTigtBG+kMHzYMoiqnlNi9hjdCr5D4I9yHpeAEV8yY0Z0cWop9mp0uGMLEtDks6toMWj1Ps0ODY
/oM6vqapfuCL3VKlTKw+m7vmDngPtR6kVDgIeP3IL8H66cI2mKBBdsihG3/ZZf4zdYNH9TXYA43e
9JbaArCUDOqQd4qkFyopEpbzj9dektAFHD3INU2Zkk5C0CficLKzZuAd1/PLzcFr9oE1M884f4iy
4pnG33IsDjZJYyX6mZLJu/Ww0e2Fm4jCm+zLzkQ2B2wgLu5GJEGiHTGK0HD8FeFskCf9xo/mSbnA
GqLzHoF+3PfvnFBkM1RFOGKbnobi+jBv+3Sl6rqXpmOw6WJbP+MkvdOThWnbBXAiFeUhefb5MJ0D
pfdRgo/0hoprdSnzoFFedvA3pZlegXLLNSsKp2R2VkRDJ6Vy8CU3pBA9gXFAmV5M+ETW3GjsN3UV
ZARA5f8THZVg5BWSLcnjYccCPlY7/rAcQlmtoYmUCcvxpxJXVno5AtCFO4xiFiNY+r7sOPTAOD6C
9EWvSketqliD2+UPDpUxsS1ThrVVC3S1tqYTTQNIbsOxMGVJP1Rm2hRxOBMJfuoSIhDCgk3138T2
1SldZwaroXomNYScUeYyAdgbdLg1QEQUPGlwtaaaRtS3vHXwO6tDJxzPvSP7MJzhjT65gCl3EwRn
HykfAZRNQRb8iPgaxBxe+LqZyk15hHdGG+9QItnMvW4u+ZxKfKKsgxING8CMn3vu7/71BAm5zy0l
X+vUpzkH6mBmfkMs2gwmBa3XJC5J7NRv2cFdGEQGkUOJ6blS+k9thSDcDbZv76gBSmYUEh+NqgMu
X/laRkyCUEj7SbCKBaH4uq5UwBb75T0WxT2/DfCj59h6xFniUMgHOAjts0rpnZZLTCygLhsDuugE
bURm9wQBVTz9V9KPYBeqMjiX3qsXJc3kjkuZQVzrwkJtUU806cnetZfA54FlbDg910y6EUlmhXCv
/mDk1X9YFQ6DmP7wyxRfvMT/0boko/l3jbQv7HicE1HMhhZIv8xD9VsyqE9kVvVkxf5UKgMxH8eI
35n8W0+loOyKP9hoBagp1RiBuop5Zvqzr1sfr7TT2GK/AozpBVf6CMUoPY+cTGKwddus+GnKzJSa
+3ij7mjL8WUU6ROADmRMP/ho3Le41kiOVv42aG4Kbv21A1PfCh8cV0mhUgu54TkZ/zDw6v9JPI9+
TNIvuWn+kme54ei6YvhmrC532FkcGLSr+GO/3GS88XO44hwfKo4YWbknpbun9DE/Q+Kz5C93jF+K
wBDaTxq+P+jwBMnjPHVTWjMriLq3yNPcUW55NOMoAJqt1kRAo4T7ELya8GbKP5yT1ILDrf6I2Uaf
gHPfG+xtT/kknnnQsHEbS/dJjFAGnyR+Bx79iFvclIYqWwrqGlji2AR014DyIoPN0m85LNktborT
dpz7V9rCHBWP2h0xo0f0rn3za8Oor3GWIFq0r5Yj6QNzT6bH3Q5CFc5Da0AZ3z43d1V3YzjFK8wz
GHdB6/B6RcTWSXh53wzkJpGZOQUsg7eYYhX0NHZhw5JB1bFnyLjeuSxka9wPQSKD+HXd2KJ/eoP1
PeD7Na+r1kaK9+yL1yjv41VfL+1h5UBHzsvbZfsCQ7S5Y36D7MC1IR7Q3E71s9KP2hhpM6kUMSSu
Zf1aQsgbzOMBBg0tRG8F0FmZY4OmqyRv1zcnwklniNRfHyL21qA6+YQSr0Z0xmuhjZlUiv1j3nik
c1pP1scPz5kIH46jjqGXD2xCMxTDbNNG9S/QMyKu/J+UTbqd8Mp5qF7LbGw/w6IUy/l95wHUgNjq
ytpgM9hyQZei9D+jcK2fEmHP00QN18jZwy2MqWXrRVHzmwX9FxYIMuMBAp0w/q03+6hU9ycBl9l2
uZ4rBsDmalkxtY7Op9UX/W7lwssofhGHtZpkCkbivNGJgY7ZDKfD1HDJedEXrO6yafJxCiFQyu7q
xKmGbsUMMUFJOA7jlk/v3VUci05dawlnBcPvdBMM1vjFuwU/CTDjaKDeqmpR1OoVpFlwSOJX82Ea
t+FRoiNkP1sr4xrnhw01VBQ4CZxcY1HGbPnbIZWY0LfCzRvlCx+JlOYvySuVotkwA5zhbmblCHJb
teB6A6pIAlOvuEl4CsJHvA/cNW3KOpbHcGfxH4UbJ8lZ/IX8t8bLwH8d71KuXi0yYktcEF+uGUbX
dIoxqRFRsHTNUkFwWrY1YGqnIUW+OiZ95U43tBd5hSJK7k90yI4cDP1G93Nerz+5Jn6wYqCzHEf1
z3fFWwgEDJdRvGbNhxIVfso+U2j0oajiF+/mqLqJ8SjSQW6naSN7ffCsI7HYHp+fMnKEJMJ8Pk5q
cbBKQ9u14smUmOX8nL8b9+pQCNM12Dra2eQHKDJXX3yQKlOdDs4o1BjIzn0AIcsT8lpMcE4PdKXV
odlcJOReWCoMkxvgA/CYQhUWhfg1qFwEhneqkavwOnleY7s5GS279WrBMDpP+K1QD9GAuR8htHe3
Gq6dUKRh7FjuhUWPc/F+5YoWZw62SlU/39GY3Q2iudxabkFh/KHeqlAwUkXNVrc6NWLpNnxPMafP
2xOUe8NlfRbt88P5xihdzHjDjobhfcdZds1tn7vTEMVHwTR8oOPCvQISmnOP+88nxP/nLRimMzDk
XLU5sGeqLdtyhlgKLu/RK5ZsCrfsaokgh3v8o0tCAMczHZb9ykwNGQt9cHQH6Q2SNi88gohGHbco
btwmjaJwmEjQTowPvFft6h/hpRC4B30bkPLcjYon58QzkmxCUVgWbpG5Y9KnPQmYS2zosQdzi4eg
GLj/IzQVp0YXcyBWVOhuGQDdD46BlkixRkbLw5rXsXsuyvfE3lQIeBIP7pB5i0B/kX+4xI1bGDdA
yC/ulFWxmAKg9RzedOXBKHw4gCx52NkyRmqdxUCOAkxFhL6s6S6Pb0iLZ+Y+gR4OJvfBXC4l5y0U
9kJnjSmNFLjW6Dp9q/Eh1NZi9pA16cLTo+0YRp/A3VSBiiJVEAjYwKC4FAMKsbzDInVojuPCSC95
qrPCNjgUMBriNEnTF4k0faA7vrebIjDnoqJ3nNHhjAN+mNRIo7G8FRzSGbooOrW87ijmVvcA+Cix
EbR9vkr/9foE7NLo9dpdMcVQW3TWY9oFCjGnYe30qJ4lRgBCVQTnKPwmYAh4mCR13BASxlAL6UKZ
2C6b41uG9se3sSnUwb6FC7JAEwgzczgxLXUjfhJnYEG9vbCF64aJ8IxlCcbKeyhnsev3uyx6TMmv
Oes5rzOnEhKYBBEnxmg+JTgOUvxT//FH/r1bOwBlRMrdK3BUkORduuyVrNdW+iL2178wowUs+PZ5
fCWVHJbH0V/JSHXTsi26oou99UWWiY6E3TDUhhhEm7wuXv4RxH1DOqNHVjRJb5j2OyZ5tA2LvNq4
JCuW4bFI9M/vuzjAVQs/m7XDGf/B95TP0UpxhRhexBYz2hrV8/7H4P6iJ7sGXltRr3iCr+hVpbGF
c/esNKi/jzo6zouW7niZ+2Lwj4sorHb6Qnl4SCIGwSdRHlPDg35oqEjespWHTWh1HsylqaqbLhjy
s3Q1TKPQT65quiGvD6HUh905//YuBguvEjWlu3OOEyOHvfCeN7+1SVsuSxHdyJRWvqkUT3DyumwE
ShuXW7HcDWQ85hPR2qDnY4M2Odb1+zznuJBKDAhXhN7Dc4SDbUWS5ml9LTpHvSeNZoueTEwM0kIO
pO8jTSlX4U4tDIhsM5qRv7X7+rCrjudMb8WfSBFz4Rd5AweICeC8SLENjbtQMhREym5zJrxlRMI8
RxfvsydgcdhFUzqB0C8gtZyKWhZjMy2ci2FlltW9aGHAWDHF3pnWOyz7vvXPHLYoxa8+hbmsRyOh
kOG/IRDy8LtoOoQwd5Yym1xfw2kgXlnnkxuHgsl80SkyZCqhS1LQkbFtSQPK5+Mgg5VERc+DNBPi
/ReqxLebfLCIRdP06TTc4ufW8t8G9qG8kaujetKi9gYMhcHi/fHQd/iPzOQn6XkG31c4Q6ynOdCD
2w3bT8mk8Z5VWqDAcUSWOzSCa8o4GwZTKR508NntF+99JRtfhTkIWXfszNfdX+fGGg76Ir+ZTCTg
Odcd5QhMfUpUzZwp+2t1pukABdE7VDHtYHttYINUk8W/3xVt4yaTFjjD4kyM4U34QB6NxIjWoudk
f0VIo3tW/78EjvMaFS/d9LbMMFBjWhPFTcIFHc9Ac7eNUhbXFMleTUdK/T7SgEuS7PJHEum+h5la
bXc8kY7Q54f9gXHja3sJ5oP/IvlLGMhp1woRPCXyZfdMZXWbjH4p3qebIHKK055nQEbnXbJ0s9UZ
iRjCvw4PjEAXTGQjM//HToxrec3etxv+n0VBG1RPR+yYj9BhP71ggMNa+th9X+YQO5+vlk/YNycH
k2+yPPymE0ySQ1S2BplsZyYO6NdP14r6VQybsHl5HUOlrIj+ThEXLIeHUNn1Kg/HTstFy/1fKFWI
5PT+1JHAxA21IuT9427LdH2m98VMqBv+TuzXIkYuV07WZ/RPFee8RjUXDvAE4t03Tb7NpM9LE7ox
c4OXj2zyHb76dGToRN5OVhc418XvdiXPOrjlzF7lZPbB5H61hQKx1/0th9YdVpqpLI8JMeztJ39T
p7EJMYqre9SVKeKg7N3aZuEkOtK+BfK+rU+cJmM4O/KXtIE+HQ0ybjZueaFzHHWDpSmyNVCnHE6O
F42579aeX3WfwmRTnqHDnkkJPtsAWiXXNkbWDTbFEOd7nQwiRuigVvoVq8kjQsaHXbaTuMJ1gK2h
GG6EnzJFFHuqNWra5BTtXQPlTqG6sPOCHFKJVxUE+GzpcLLf/XeGJZdDY1oXd036tV+DgCT0AbfR
LQPAj3Afg3MXIFYM25mDCBdWJfbZySlztghAymIjoaoU26HWKD/ebUQS+KjZdJaPWBDay+gHRpTy
q2M/dbnM6/PtfZr6RgPWIUQbcx3DmxT93qT0OHN7KaPhETR09O0+xs4bMI3NZIPwU4XJILRhuc8k
ZQRsJmBIVoVFlpaRfbYmPOczUcokC2mcRuCThM/hcbZ4Q6JCFqzPPkbnzvFdLftYjdP4Fkk5FSVW
jOcF/ZfU2zijsEfhjVfpivJyFQUQG3kl/ptRhY+Ib+I4K2ZSDy8ynPuu/M3787lwy6cxFJx8Spn6
att20jpj9yxXOujAQrJABpFy3Fcj/WUTYZE1NfCa1tALvEam374ulQjQ/2MB88m9HZsOS0x69cTb
ISRJslzUZu2LlvJJ5VN8F24GKauksXOJvFSl1zGE71QPXzWw9jdnW6hw43N1+QYxl50mCyXziSi+
arGclgw/V25qRzEx/B0YKGr6XZhuLvvCUJld47Ra2dhHIuN4j++u49VzhrZEjXpLplwh80EIUNMX
LmXs391U5290Ga9LSXnLFxyD8cC5tIHRF7BZMRocmpgCoQfV62xqQCNtZnLS3JJiT8VZfT5HbnjC
jgv0Y963sNIIpjyXTsUTbFU/JQLmhw2BptX3loWt3k6OIMm3d+PRmE+dpFDHOwZTFWKMpZeYx76u
Lm0R+CNEXzpvpMGqqTJovxp0Ts+Ej5PtA+Dnd7jPPQ7YLcb7Zooykwl2baHeUGJFYM482nC9C9YO
fiRtS2cJTCa90CrHyGLsQvcudAtpeo87jH2rMC1b+zed0YsqmREJJfq304htM9/YlkFfOGCAaRDh
NMFurX3Paf1CNjPfw9caOSIaV/jJYr0/tL0J/zzg4jgaMLX2s28OgZSuPYfAqhSg/NZRY1DgW01A
Nt9hu4/Jup9N2cCFMqzq8y4gT8iE1hKam0XQ8sjz6b+MjLRBKvbGHke8l7IjcHtjzxMogeERcYUt
x/VpcVw4cVeqwFSe5e2muxn7te2rjs5mB2eN+ig9P/b2XcUqw6docrRuEqpawbwA9Awlx/TiNjYY
ITXXSECMyKnoGFVCzlmOLEPQetxdNKwk03TKDzW0s2UrfGt6/wWjqXZcwaupArbFr3hk6Kh/loaQ
g8J1G4s8RM5WWJBSq470pEz+gjFKr3i4oxvcJBcxsIYAnmVV5O4Lr0/AS3rMF0ofAh+4D2hyQNly
ybp2HSPCOcxu9VpNvNApF3/dQdI3eCt9oxbkr3vieUXWf6z5UW4OnKZ0bQYZAA6uID1Ikf6afk+0
0PsTd51wl9T18RvwGivO6v+nG+CbRTytZsulHyOPuZhj9dtjdQMPD5+06kH2qNEH1AWXpirLJn9q
KBeq73qxduDOTCH9ePIkiBGiivVsryi/Ra+uDVG8U7wghXdtVyu/SwWhuVjaJWDripSBGsHB/3kf
VMBE8K1GWHtH0CUMH3tQU953kRZe4Z386KnU+U7iPBuMkvTtX0TcClismOXgAEyliGFfywnBzo7X
Bj27vg8CGNeB6xuzEzrcey+QbBSYhKvOiWRuqf+dv/i1n07TRcynzZe8TOwteglN3mDzgj6Zb/wv
i5US4gJBKxuEi1lUz834BHkA3G59NHSS62+f43CXkyJVxS+sJS1g5IuT4tX0WpS39aLfpOmdOqvI
jCfuYlOPpBxjt+jQObUPVMasFq/hZ9EOMZUNgn0eoUSiJMoahnInLtyMR52vM1YxmY33B3OyRn/z
HEcfQGt+g1mOBnADm2DzyWwVU15QWz4Dh6vyR6c3LR8OkdS2JcNtl4Bgg2AEJW2SUtlrqBzfgSUc
cbdFC2HdDPGuwoZDfbAIvutmqpUqDFoTSAjm+uJ6b/ALyU2fVAqB2oP8UkY6BC5kIvaVPCbuzY+p
IyeBb66a72oEPXiHbxuPVVDvbrAiTC5/zwNO/BXd1dUoDsLEOEsvw4y9tkSscTHsRg7DksOKrqc7
ZOLCL0Gf+AVMg1kXx2/YtMo+EskFjA4UdZwdyBJMvifRRHvos0HNDbIc6bbEonp0mqUULkJLxp/x
xzyBjRVSvN56s/E1URMeXfXJcjOKeMiq/Pa4xzMW5gQAnYpZNSBik650kOOaY874FH/iNr8rgbAe
2wG59zGBZtQT1Z7HJWpQsy2Y0xFUAmsvINRU3RNO/L8s8ZPIiroX54dTuZ2ZAo+gIOB0vi1yjxmN
Q0UmM2on00miUZA5iqSPXllY63nzFlI2jBjvp5C+fApN4eBCt2fNyPCGpF3uAF1Fd5Yqlxi0AgpO
DCBKr3PSD9TY0/AyX7bkPFWLUy3zFMy3VGFRm0t2MHpOz8tnxJc0K2+qMSRbh6xDwXWFCAQPSyM2
mkOufL3spuoLk8VMwmwDunKmnSfaMxRWsz484G+N93qiluyJ7tRbXAXKkGQHoiDIlSFxkxvqjgcG
cjqMSbgp05Q8AETUmG3Tx1jShLcNOGF3l3bW7SsRu1TCStuXO8aFmwL+nSVL7mWWoMfUQAggd05C
CEV5UmfXkIiX4xTheQe36DsPAVxUoFxtrJ8xx0wJm4My7iOBAyPdbljGvWX+gBIQGbY5s8RzuYmR
7aRfzRIAFsxxZhDT/SofNYonVSf/9FnlgnGZPAFchf/SGumThbxrqX/44fJf1lh4FJNLAuoqxRmv
CTC8IqA8u1dvOCRWhDAb/WZCd54/huD6+2xL1PBH1IPK98hrEzq6NAfA/uEJtya3gLWDnhmiybfh
Qrt+cR9LRbsmWQjzTOEaXhxf3r0TIkRITE6y7f2IsQyaDCcxgnbx3bXS/MnKROVPMqGYN5H6ut2o
wQRI/YzQXRx8mmvvpgJUfN890qO0tD6OFDRHbL0Vo1Hi2p57Vrbj7iKZvLwf8mPuIRlVh4rAFGlV
7GzFmy5gnl7TXI2fZ0aie7XvpVRO8LpoXK9+nYMfgF7oOEfZ500HifNNDpuWl2HdMYRk4sRtqKwr
NxlHEwS+T4I7QOzr4++emE3Nx24ed+xsZ9I3LVj59jKWR0gjiCAu2z0shD35bJeN4FXRPlFlDOLo
oMYu6O4b3qTbhx1yTXR710bIcwx5Gc/QKGprI7I+woE+iEJtHT452SZgpmrkbQ+M/MS5JdC4AZVG
f4krXPJYVh+0BOyx5BsIwiX1NDowrQ1FM+e93OEQ0RnYXILbxfj31RBgY4xdoOB0FlHDSUGPKmfk
9UOqnZ+xeaMbRpLdKFMm1L5cbV3Riq9fPmvzoU7PfvCC5u3fpLew2SY9Gc7i9Zg6usox8aeOwAAy
NcF6lJu3keO8im4q/eRP/FMySHjX0YPVDkaJRuEGuiD5kr8zj+tHBlKJkYZYLMcJW5VnpbaRl6aE
mzEVZM2BlJbuiMOxx+qBDIIwWTuPkLB14bN1o6No2cDiJllnhjS9YfprmRcBLaYnIHTjaDxQL3Y+
xrUcwWgCk4R9hbCedwLpOhPGtGfGQWQKC6d2Tfm/lLB3JMewEg4lm7J+cF1i0PHsvTODguTvwnOU
ydsd8oes+PwT8SMDfFub23gYRccJ0Qwef4rgZp/ZzU2mNXoKFheSe0ROLjbVRecQIcowYz00KWu6
ncMWOOIxVKKr4mmRhMxnc5U0i0YsAbaEt8TzEu68/xY13n1BTp3eaEnGG7m0ClksQEMhc3B92aMW
ujfDkc805vu/cW6uqBd4zMY+dzWGC/nYEXHZzfObHTMC1h5YdKUKYXoGREKUnk9HP4Gssh/hNeyJ
KGrTTlC/uKobyROJWqHjiShzDtSboDXo/EUXCFBYHc98rAtXckEeHoM6ctz/+/JPT7oUo695dXq9
az4a+O9nfN5p6m4uTm3BZdx4SOeaam0PPLSybkyOMpE9GWteASaBmkzdchk1fVoiZj+/b8ZsODem
oQxZz+i2gN6uHx22bOAXrV56wnz8oRESQAHWf3/uX5UeXvlb1pQ/SiPHtz1SoRuTvUdOXG2QpFmD
sPqBiy9nWkM5wAPkRcPfp2yzZspKPrtd82fZG7gKsBwje30X1rJmvUYyZ6rtiKsNc7lfbBsYZ8u0
F4UALz2q9tnvZ5e0uahf/7WGAnxdQUSBs39giEOr+ljDfuf5Xcy9OhlckxhECASHNDSoCFNuGw6b
HN4/XSf7iuZRld4IqF2T8xo2/XPx7QRBxJ7QIUD0ekgj6YbJswBsFzVoPExaWfWjBoI4QyipvVo/
9owj+1Kino5Z7Vxqecap2L/9z09VxOlxNzGEJGFJhPBx8/qd0jm0iP56MkO9qm89RP2BjwfnPWp3
esqv0DyNiMfNZVBYJImgX+U0QR9CmhUJTsj5XSZY6FyOFWq6LS3D4jW6vgfwhEnKwg98iGRTKtJx
I2SCHTXNj8TStYV4lE8Yso4dvMXMl7qi+C4rC3d9f+DodXbnEPywvyQE2jovEuOQ+2+3c6jRNojl
47q6eFgM1cdwfzOFeufkRTCHVZ1xGL3UZ3+UR6sTdS+8tmDIMz5G7T3McWiH+MnEYgthmZ5pDe0p
nxYbL35my+n0nt3UzkT4BWibYMn+rOjn1v/8GyJAaffGMqXJL/k7B3eynRpQIb8y5CpSOM8ckX27
FZSAJBPmr3Wnv2IBnfozTeSiwmOR5VaxxK3CSDN3+TR7Qr8BuefowscROiz7sfcOPxxqdaGBaXLa
bu+gjVyUAVmcJqJsNt8DqdfUH4ik0YfVfZ00TNmkMuIbAMOJAULFfWtGDsJbot3a9V3xVhgcNoRR
qHt1YAZb88VD0vH8PDph0R9kF/6YCDM3vE8e/2CJeM9AmgBmecU++QsUKHZvJuQlv0UHQFln4L/f
0pPD4X6jWnd9BRet/rj9KFyN0F4JwB2Ksl7nJ5oLnxnfRrK/wJczedkF9AnRrMY6KQ14GZ38VMmH
GKDlxzwQDVCSe5j7og7eB0TIzhf7v98nYr9CpidccdmKXMNufMawLbaVHzS1agyUiyOulGE6rAoh
znwDgkx54sfXGeV5lyWiyljOhU6sUZ0p6barGAv1qpPpvTRqcdcainTFAAlaG9rRTP4fb2KHWScP
NAJ9q4F/WCWj6bPv71C+GmCmJt9ZmENsfgnZaLmBcgPVwK1p/7yPJUf8Iq2V5OT4+PmhfgsH8X6f
eTRFhGFGBN27me5jedYR7W1+6gqmeRhTm+x8aQpwdHfIDIW/+rLMeCjycOxrKnkNFy6X9d5dpJaD
yZJ3f2vrrkUpyDpU9W89e1LVwwyAIrY2T79kmLlq8khfbO2KN5U8IMXFEhknZ3SMMNXjgXFL/tLC
qAU5b/4gIamQcDuyzDqks0iZGL4iNJzgLJ4RVfa5YScLtT7S/8qwjbZGHVXAp9tFhwYGeIxxY+UN
xvWOlM+TKcIG2HiTBoM7LMUsW1XkuFS5cRs7wIRn2LxYFzKDjzURPOsf7a/k3YnvlKWutum83LNa
pIL3K8Haw496dry5IS3ESA6jAemjRwJIusrnl/PlLbZtILbl/X/XeLH4CcMAXyxneb6hzR0wx+BX
tGzWp6kgA37YJkGUf6Te56AFbALdAVJXevoRUWxo9nAg9QjFelEcJs0Nsrf70TnLujmsdxmbC2M+
899QhUcbPTUhwa0C4GkahVGBolhkkOFVwJ8Jm7UgIlzJSsCORNIdAVjWOEzun+p2W4O69BNGj61c
s62zwSlQPdhszPqz1HjrJORUHZifTHLqKeo1GSpFIxrV5lhZwDm1pZsno2y0yfdiB+OTCn2Z1P+m
yDaN2mrP5w4HmrdawBjnT2nfYCdWp/lutJ6fVbYq6oHeMBGI2d1qzYtK1MZsGG2btOEMmd5w1i9o
1wK3ec2ZZl2LodNygpx23MjyvI7MhTW7wiLTNtNG/kAHtG7cYwiArOsVpjRx1POmYCVG7CMBAWBS
BniVQZgim3IogzI4pfMSMZu+oEcbA8nSV1HFMhYOUP7bSO40bap/lN3tovuwbGHSVUKbNXE7zxha
BZT4JNagpfUPxseyjnw7cForYDjSjxiDY1UG64UzwEPNE0s3fUfUVzW5pKvRw/SlMDr+p0C5+Qbj
Q9D+OCr/Ctda77YxS59E9t5du8VNYeVLMkkkUtIwDzynRkyb1ucSXYHEer3naCQwuXK9+mTPtQYS
YX6kxXrDLRs1Nfe6bcNq/MMKc0agDwBsX0cj8mmGL2fpE4dgg1nX9B1czUShvB9yS2exaxjjctQ/
X2ASu32a7zudz//zV80QRLMJAL/QDZBC534zDfXiUrjm7wFrYsmaCmZDEUvGgfcHvRAQerbSlbPK
TyHT3PCu+8rYUH4cNZi/mzhNsWiFPZ2er60838EnzhTHsdEewkkbvmI1hA3GwuFV/OJPHa+Ye7b0
LSl6+WAwA5rp1+sl+/UGI16wS1YaZ2jP0ua5PkbTXDU5T6HkVjEg9cyG2qrIEtBLhCcbSqbGiBn2
0xXo4Ha8vLM/vGnIPvErIwCNmnpPZJgwHCHDi5mYauZmdIViYjV//AEEj/AUMDxgd2P4ewvkQOZd
3pd0y2A5IHWeuY6Go/Yu9zE34jaC9rB0XF0khVDPLWJ8o0Ku9pghvIeHNTCgk9q9Q4wwsM3+0Who
T49akT7CWfb0crFTkOHedLuMcBTrafLg+Yoo/mNqNuvuXrKGt+zJiY14PfAkuHw9aimlECzpHmUN
3Mm3rsckahNwvPFFsyabmRDgdgS9kkynCYx/SIXjAxfDflJIA2GkPc9gWwivYfM6aEXvXCY3z0Ko
l3p34C4sm2BeH2qlOAN2yA90VIkL90nYEsz0Ko6FFVYs0j1GqKWeZjDOdH4E5oBd3EN/NrBf6XcV
ttRteJHzwrVIgo1k5FLFBptQC7c2KZJucHL3hoaoZEseLvibd+My0YSBgyKgbSx6wRcJzYPcnM2R
TbJB1e8403DJnACoTHi7Wc8GSWB5J55hqKixkpy6srqHFmcPh4X8iHy6CVNDh/EmfAer76hCQ9PO
G7JSntU/Dqpu+zBsy8BaJEUL0bKwTmkE8cCpp26gJzzaO4adC3PQ5AYp1U+MvOoafEEOvFro2i/s
YVBKV4MKmVKsPeMEuiGMuRVKRqykRYvTXwzsNCy/1PxcWpblffz63HoZBMCR3zBhH1ZSpbepwg1S
l/skDeKLQVq5wuB+SlZ997rMnkm3ELeeXZ/4Ncw7vZ4TInXRNcFrq3qWAvMlGfaPRHq5gz4Y1g3O
fVQfKLJLCmxq/DEQGIMKwEVyr5ad1eGy26WcSJXmGL/vlS6kf+4aEL+1fK+fIY4GMQtgkqQV1vHp
hgmlDvzqkB2NZaU8DS/bOAwurSBdYL7M4A4/cWtjc90fdP5nwzw8+cE20oTce7EkYz0vWz4k9Njx
+pWdgZ/UcovMBcxnGKFEb5IJpe50djDeHjvdCuni2vnLegn5NQdlrGDAAXOM7Ny9qbXeYze7iUc3
voa1uBVXlVcZMr3SEv5CiA1+TIkiEGCR9595Sorf8n1JuXjItdq3ZITlJDnfmlh+ze8XuwDHzvvN
a7GQELlck6NAl7psvaWSbaVcmN9gyU0uFHyt9R84S1R+CtqUBxbQdqvd+T94WMj87bXdQ5LNgbjg
fF73yR9DECF3X+u1FX2DP0VsVq3x3ou/QyEaAcijntB2D4wLsLBRkY1EohAjQOTRhBM5Wbhy+fL0
OvMVZhIQBDcMTDcQgsOiv7p82uoUMFNlj0aerW/ll/yrchHAvCDTQQsuzWKAS+aTAvtI05smeccN
+LJ9hN6ZbazaWPaR57AlTEiGBfKTPSa7kDQRwXrpRd1O7nkZkT+9oRw5CzofIglyATBDILD5QQ5k
TrjEBM1qxlxiEArODOX9xhmAOguAYT11xx/zTHpwnzNJjDmKTrXiNIkKVxZKIzdhsl7GWgCn6ZW1
XQPeGZW5b/6stzIzUz8GuauxJpoQfa+2sc8mGe1SfPkn35Prwt/+uGm738NFzkrkJhNwMCXRAYKq
z/0UOGZiytNStdDgc25FIWKbgTeub88eHlSzhIYmnuwfP8VNjSZsmYe2h3wcWQYq1NHkj9wsFAZr
0wiDtGvc4hf/fliP9rx/iH5WN7QvHSiC+V9MqXl7AQlar8ZK9DlND8raTl4wABHOSSauwMudy9bG
+ptXCl7OGCNpkV65tjq+3SmCc270QF5LtRdc4w9od+cHwNYXHBxxkW8OQkR4KmT0E1ExoewvSLcZ
35zO6dwa3DCtF5bIG8os4O2vwcdI3M3WnZV4Ai1pF4DY5AwoNMQA2xSFjnh76ki7tCdrg02XElep
4v4NUe/HDDC+dRSGZPZlpfnWI1nggEtTHgfrZM+N0BX5wFt10aDi64cFDA6w0rqxG0aKF+L+qqRL
3D1GNzKaVblefQ2GRbOUMt2GLHsyZCdkwokbJOaSUlRbOx7+EWOANTlW1XuKpg1YGHjc72djB4i7
jX+QYtXwBQObaCj65VqlYcT6I1zuHew181iLYcRZkR4Topw+GAR6e7Yaa3xrE50l7CbnwO6mPA81
4wuDWPxW7S/LQ1KNBDqeSmjbpBERw4L5hVc93K5vtsglW07gcaha26+Km9/HaPvvr/xGAA6n5mpZ
0ZDBjFWhDBLXxD1olf/vPGwbGp0lZjFBSwyvLUHtgNcolwXHG2QAJeWv85KX5fxWWvp3INrkokSO
qWpzkKOApmb7hsgZz719QJrw0fJU9r2ooPA9WF2IXjjQqXpI0fV7iGm0yyR7kw8PPYRFzj21gS5r
0F7ZocccD5KgpXVJwpDXDP0bQPpLculnZ3LYcL+bprn5Qg2oL2SY8jwCX/PDx93cg9zeXQAOFiAu
Nc1I2V1r6Ih07pKkr0SLhh604YcuVKrkBBJi9y2UVHLUeGcmi+zFpEMyeZv96/T6do78nA0CIlhL
4fOHp7u1DcPhZkMbVWyFNxe8k4BjYCCe5jgocgF7G5VyvyGSRJbrt2ucqCvrihbzferTwvLIBA5k
VruCEazrBF3dhoE723j2/3KMWwZ+UM173lIKlbYgg7Moc5jx9UBvPE4ZjctaNUL5WMwZ6vU61+6u
t4zX5DhJNbSMUYhQ/dWPC9rQa/FUnoqoVXoVvEBeL6IqKOe4EmHuyfHkBJP76FPq/EOE5cbEoOMi
FmphN9a+DP84IswStGGUsdD5GN3iCtX8sWh/c5sea1J78ZnwoD8gUWQX906NvkQA1adzKPagGxj0
Oplc5gPsq4AYeEOByweBtxNnRIKeFVE2tJ63u5Si7ARrebiJV2Vg7UjWEJINpZ58KDW4YZ+8I1Ag
0nFFj142wVuB7ifVR/eyFjOju1QhxSlW4u+DPcHAVXwCkNFJGIR8hL2aErCyUxUJmuHRD1jURWMn
T8CDbhrzgZX6RzSlpOf0iZHfwWjXrUFdFElbYv//GFu3WWOpqRZNTCiazJFhnbPoxsZKm5zgIDHu
xEjnDlIuOtiS6taHlz87V9+EWP6EcP3E8uoqaqw9KCqFzEU+0tqSlGyCN7hTXofD22704UAbQG9D
+RkrqrIE1GcbowsGD3MQADuAhwgjZH7hWeZYkVCuNxbNem9RKrx4pPNgHpp0g/WM4tkE+pHLsysN
dyjA8U1VmRLQuo4/5bZ93E7xkZnbXtFTaImcGV7y5VtkIqbxij01qip3IoqDjK5GkNI80MfbEhk/
o21uzUas4DGBAb94EtqKl+Hlkul87Wdn/ulDcrz2rqt6vfc3drqONzeFO5piKHK2l4796sqz00Qk
GLcphMTi5WaQ+jSZ7y6D2gBWPzih0TJ1ehDUIvcJQQpjJ+oZ/gd0XnRc6BUW+cmt0uXeC948HNBh
ZuT1eQQra132LmAAQIIplo8iZxRiSBkc1ZZ1fptPCdahlms5+Z0Nq/igj3d9OtswP1kcluLfDvOd
JhLvQEk0Eby1xtLRNVM161OwqmkYoXsuWEuNpDh7RRnFpTUqSnpLRG8eb65NxfPKsrgrnKCAMij+
jOPNkCLiFPtwrYDHiaXVKlb1dG2PvPzEO/b1jb5aty3Asj6mZtQV2CHjhf7IA8paU8LPNM9xQ5aJ
eJM/DKU2+4GVyoQtLH7MyTFW5gtz8/HKG375WXGc47WkaVqfi6TWci7fn/3IAuN/SZkNcGoTZ9iZ
PcmEsb4dzZ/5srWllD5QYPTKJOfm0kNcKW+ZTrDBrgU5bI5F+ObvrRihf+u9emtj9qEdDAVlzKC5
dJ5ZU2RDpsw9dc2iXKA1QwGcvZOa/oHHgUX3+GuNtFaZ13MUgl/UleK5xLMHWT8wiy+lQtK9AZxY
JpT7bf7kHdXQ7KjWTS9czVTUd4UoptDxvTsD+IioDQEci0UpnijAzkiwIdWD4cPJTOl+B6WqOP3W
kbnRLAwJjzcuzWiP/WiMKqskt/Gq0uognF33HOSkfdJT+hXklzXyDInFp6m7kVW77wrW/MDbX5vW
nx0ZbXsIMx5u09p2pf8FxXcsww+K+CMpDg70CwpAozfBCuSC6E2xcvTW8RktN/UiXkRFaKTAycFA
pZY3QqKEt1P7nSKyh2zku1E6QAyVfStjoBRaYVnroD44WLb7V2kZyp64MHnk81feB7vxTUslOZ1c
Tp0k3VZNChNJg7/VvAyu8nFjpucf+PLtR5JXdqYbB7bBu76yC1p9yo3hUYg0wKsEjnJs5NGr5AnH
JWkzh79LAYiClVFJNgT/msVsfQ0fUehh6cE57MLaZZu9Bo5HIJb94vmnF3hwcUIwsRkswoHfCDqI
w2pFVlvSk//do1dp3MDBRDdyt5L3Kh5E9r5W3FaJlliFrE4UP1FaaaOl4gboJ+7d+mqGxqSkRU5C
p93Bvq2F/tWJf2SH/1+VG7YaPJztdJZUYOcuyChZqwA5qizjhnatKYP0w08eD4XnA3utQ125XZKQ
gfZwzeDCQg+h7fmw6F2IqUJwlsblhlOqhTgBXEvMAlpEe7HI8YAsbxzD5GSbpLBqP+dvxgDzod5X
x8vDkzi2b+/LjRhzmPXryrcymtXnfNzUXN9zwTFXjDhopV/OZ3aKwW1OYDXvC0sNcRVlLVSIo1F1
/dO8zvuvP38Vz0f6JU0gRGfVK3ip9yzDmXkzUFh5vPYimPKEPJ/ilcEoJUJctTZSgOyCqjKlc8ih
pY8CfGunmLnwhsHOLalrgJZJeZHixHMLqvw7UY6ZpHgn+qnPv7OxnJiIlFXOg9aDCodoVLSJEazW
yr53VuI+uRT8YbAAOHnVMuLDinq5FJY+PgYw7g+hRx2LPXmSFDdXsaMGqfntq/eZwEejg7EQbrJl
KIEQSdeLiLdB6NiAwFijZdoXlWPyf1pvHjywgv79LEkwkiuzhwaqNZavdeqXN1IBVJ8YlAAiNVdo
b1TtMSPp45tFtN4aZ8tFwpge338saDgycgGRMg85MDlqsfvCR5hrX0NQAQ4x7FzCuLyQyx8LdgSz
3yM8eCLQVFEmgQjzVet8UZF/f5v/T14F1QXcszKhJGXLSUnt9yBjOVmYe5E7SPJne9IGIFnzjQKl
LJVCQUB/2MGydPcRQw28U9TUjphG4sy6nNwBR9sADD1ErJIb02Jj/FVbCJ68skYIMX1+JNyLZVf/
eizOHZ6ioR61Q9He1Gi5RjqvefccHdQEFQ+2GzZaWgFbyOlrjHhg5vcX1baBCOP4BJv7BfZWNbAL
am3NDBJnpPCISGux2gUaIyF5VXr8Jel7s+Sd73n154WJ4CRUWRZvrgCTHsVlf/IjUBhDMuRzUkDn
037u9Itr/3E2sAndN3fVjKDIZsUccod6V7dmdYCSQUdUNL/Ms7YuQZRcrT4nNL19pkj+/o4MLhIF
aKubsPUJHElLl4R0hItwn+Pf0/08IFumgPFyBF0idMhFqMStRTA/XH5LR49SZUEYpH/m5ri9iAUL
Z0Z/W5Xbmezp3ebRT4EnS8E9eHHsX5+k8Ub1XDxYfftPdZQeYLNE6Scbk515qY7CJIbLjATo/nT3
HtjW8dlMgiuIbNQneUj3Wq3Zhpjuj/Hsykapig+la5yC5kvnGQy4CFYm+oxJPRlBT/DKyAseLJbQ
CZRVI4fSWqpmpfd/+KblcZBr48Mkr9V2CgNmY+Qa7cO2ilv1XznIMra5xWZhzEnuYgZBVkFDZjJO
FqapzZQfx5aiEkU808pEu9LCqG8nI767GE4xDrMxJWN0W3VoizAVBMZSiRfltFtMRVD60pntCeEu
+zISOfMzJwRkodB7b6/cu/rCP75IJtWjJ+DTU/lHoVPd6MDxFtLVHgwdmLKsn5vtF+T0RXO71ez0
8BYgo9nI3wD9YD298C8t8jXwol/RLUpyStuILWfzwaaiZNACp0jCcIcXGohuBa60qGvpbMv3+9iP
qquQUlX62FVvDPYTS4SR7gelogdJVG2esJPevmzRMFZ29Ooi8md1SGw48u41aMf+vu0f1bhH4mwb
FukSSE2ZcXPJ7mGK9C6U5FVkJ3I9n4Bs9lYdtFRbt3BPjEb2vIDImnXXYYk4FhJb1fW8b4lro2Tg
NCYkWKCmqLwcCE3hN7Fojzib7wKM8W9iHA7GuRJZYRTshhg42C+kjpjAETuYjZDJkHh1mER8PUBQ
OQvxhGaJwn7GWLPlCdDx8JeEPNFzfjc1BTbqUz40w8taS2YqJWm7cUPt1uYInlKY25ViQTnlMhOT
1F8p2/PZD4A/PFdNTPAiFSHiyMttW/IUtsGDIgYO7462XwyArTaWJ+0Z0qQKHmgGNuen9vZvLykU
Y40kw1mFKu3gp1RjIeG2ot3ewMyJNls9OqAvMa/UpEEFwqXNa1/YlV+VPuVtbaoK+iWFqfd+lhG/
VOnW3hFzk6Aals9BLU7OdwcMO/KP+N86s+yfYDRwB3teH02ZmaD64qB/lkqEt/7hSqk/Ff9P52fl
STx1rwpfr7MjsJumJOWmmliYSNtGkSb7tEomy3zLAYtE8Zch5mYrM53IClwZf8HNND1rnS12i7rK
1zNaKAgElYwdIttmy0PMsFGJiX4JMo+YZlFQETtQG9d1GmdsIR5WdXkhGzvBmwYObqwxJ4SQLVce
v08XN55kUu5A4APWDV/UVNcrQj99pHw5f5647q1wsoZYpaYe9NziEc2s4vaWffh1bGNUKNLdYshY
gEPnJKGRbeftpRW08IWwuvGTnWBEV1jfN1MtbKmToqPwy6opLq9AyLtzIhU/jlM8JEcNB7Pz4eBc
J/9aFDJ+U4mIVDIP+XpGo/LvMenPZ8tLCE4pSAOHviwNTxjcWzyAF4hBWzLzRGvLdMvvNv1v5fXX
S1CRCFID1GF1ExkPn34S5qXH0i+eJudtjl7mqaZkDk7x9zqea/GSC3m/Jmsh1ARCpxBlY3Tg+g5U
CtmDiN/eltUcTNFSlFZNTfr1R0OLC8sh56HuJS7isRArPr7ujDGIkeED1lXlobOLzF8kh9y3wUC2
SRj0QoZsL5qDwqKxd8HYsxPxzmeJgvUulSenXazgNnfx0GJiW07BAUaT+7j2pykuoc5jkAQtpSOF
ZAkm6jhHBMBJgQtcxgP5Pv36NYW5ENcP+DA8CUm5EWcN/2gLXcrWMdENQGOyh04znlNqwc0V5iMN
ju4+V6nep2r6zAQdsDfPMmrwli8307GrLrdVLOPgLRSZzVu3Lr2ZJr/Hjk5S+pCganM8mnI6H5cP
4PbwOrNicwbjMpvnivKLOIbyIDoY2QYf82XY5GBuS9Fqhzop1unajlGiTJNJYiWGb2s6ksupjUA2
JOWGTHQEbUza8E+qdBHQozzRmYDbHGg8QAr8AsQcp/ILASWis1iAOWpxDPhCEdqougZOMi4oBcGv
c+mnZ+vaCPRakgWOHC+1Iw2BBFhx2KeUhxcRSxkMtUlIsUWdh9+SeJ8lDD4YhDWYN7EGSP7p14tk
yl48YeXvkU+n+J3BZX9zrimXMeKesQyFyABikPKDutZFZ/9XVapYskr3BG36CWpB1CT88pCOPD3y
M6atPCRQTKDUYZyg6nJd/Yl8GjFQVzEymILciSUq2rbmYDXQwzxZzOmAwLp80belE3HqL8SQVO8t
thsVsekBjuZ1l2Sa+3Nwh14mcjOKrhUY90ZSgLPxUf7GTbER6nOcKebXN8yPGxwK6BCvLAp23gLV
LJnzI7WlGKHVgwN0TS4m4bNCHxz/ZkQy9rXqJ27FH8UzRkHxTeQivC2+QI0QXDoyOtEzeNlUHOk2
xzSku4BgUrOA8+HGBgm3DRxNjJTKep6Cpp/h6vcsDGeoLyR14Rv3WkNjdaLZfVCAxfquKR4XYOpS
yDdWFXW+xSEAKHibc4PoKc521W6ZOukEcHqVp6owZ4pDL7KT94HJU9TIDjqpB8sFGAq8gYDCZ4mS
7ya6rT5bpHik34XW816yk8aeTAONNmpvzVDZUo3Lr6NrAgvC0iUtzNPv8j8Tjx99FfcWy4u9i1s1
qggGJPhhV4HAOdOEmhbGkcoF7FOahGYaDRdA92Q37MZiBAWll+uiekCQ4IkouCIk73VXd/hFzn24
Gk1/mpzOcwgm3KYvqxzoTYX97msWAWeC0V8N9UBI9PfX4ccD84h6GlQsuAwfHk16HgBySQpMsagq
hSIzZ9jdiLvoCU/ekX3G27bWsiCzV94HCxiSo/pBqpSVMRqsR1dCxkdMJ6mZTf+j5KvZ6agI8JUV
Jh7HUiYvJgKBacXkEHyiFI/EAXiHSrXIhEasGAMKmY1zeeDku0FT7sOqEkLjw5p3/OScv0Ig3du7
EFZlQ7AKO8fMBEfjITzBOeCA4jrTyWD4k0UdhsKyEPRlWr3LYe6izxavQKZPEk50I6TYh5DOMw+Z
hDnWbpcmtKdozISi5LnLiA2cD1PnmRKAzrxf8soDYVakMcI1/g8YthF6CbBMef+TD1DUMeB7XK6O
B8K/YJNTv6GSJk9ULJxWQka4xJCV4bYrSLl2SJpGRI2+Vj976QmwKZ//gotOorbIHSnSsjAd+AZV
Tsw8oupYIKb6tJKBHPX1+SrZhyXU4LdBEftL/U/cOP4UUBJtp5OKfEj9iEKy/0Hc1RHmTHXfmYK8
qh1jN+i3XSMEJ+keXKfJdcmRfMWC04BGM8zSro3u5EicyUdqbJVJfg28pppdQFGbS8F54MyR2cYQ
MHmWd4V+sjbS1JSu21XdunhFUda7+C5AQ3OJpIIcQenrJgEo4YN0slgUaSVbCbLEwFqhtquPdXuJ
Dl0om6JaneVotPJEb5t6OZmgo4kvlK/d7509oQPPMbxDL87tHd0fTOEm0iEang8BrAheKPsgjGFt
qCOmiAJrLjV/KaduinGbjOIUY2YqcltuufyfoGTHvaCyG1zhKiHreuXuP3t2mQh1tnog0CYZoK+1
FcYgu1VzWpyjOUUJFg5bG9Som7a05wXG+BggyBex3sBFVpOZB/epfTVCbe6ZrWZ9Wl64wddfxNcO
loSZRpa4snZSy4Fp44OWe+U20smwvc0iFbTQSXCf4NWg+hTGoxGFm3xlvY3XsJyeLkhTgbXTtpVG
kzktt93QyVsKcWfUKCUh1mkdfrjizFJB8/EMt7xnHkOMJv3PT/lnYkKI1ic4EXPKmEHT2fPRar6V
vtj9ZQOJMmrgdurZPanJ/kApNNTaa3Oy0BQBimWn9y6t5UAgcW0D/IKNrr0kQYe209DQAdScNqIF
W/4WFg+42t0rewoewYGreRAYdpmZS5dcMdrdJkEtWQ7KFA0xkiMiI/Arovcg01t8xJbjRHLQyTbB
pEIcPQLddQBQe4Ryfsx7Je1wWwoaGz9vjY0uKF6Cx5g0Q6dgWMx6QMQoe4lLeLOH1VOTGCf0+z8e
P8/rq9tvmtrgbPznto6MxYIBfA91o3QLM+1Hh4KlA0+HON5lNkRsrFu0LA9I6q31RKKLnhgWod92
jQaaVkgnWaukisAbz1HBI767Lj7pK09Jf4KDE032s+c2nn9IKoQmwQHp3xIIiDPSWJFipWymySAC
zQG7u3mMxxEPWJVkBXJw1+h5tu9FOPsGjzX93+NqudGBNqHSAT3XlU1UdjM6XsuJ7OVrwClIn8VV
aMeCmqOupQTmly4gE7pNfsCdW/1RU7NY2WkTMWqF81kAAZVXYgkpb/kzRBgSanCHhqfHQV0wBR3y
1pkJJ9obsBlgDokTyXNa9Pu3m9D7AhxKnQRy3Zn89mppaJa/XV/MN0oqxJ97rpzfCx/E2eXfiUhG
Aig3B+QL3SwKkZXtRRzUJKJabIocrgyH4YnJp9MekKS52mVWFkWcOvOd0MVwbT0o95+CrGerxwOJ
VsgzGek0jfqDo+gqa5AAUL3Yxn/nMBleEEFojqLXzySJ79DCG8sFOx7HYaKVcYGU1yMawHOzUqZH
WiL9K/0/K33jslsDdkPVrtp56Jtwhsrr4Cl/0JVZd/o/Sb8AYuzrNgRuJeAjo+ThoBJk5ydMlKn5
flyaojJPGdo+iadYJ8584al6b6eSwIJiZmmPPRkyJ2Ducx8gsZGshBcoKYP+org9AtlKSd3QReu9
i2gEy3Zktui86ohd2geboYQvbYVQ/DszjmysUYhPGicDZst/RKNaSeeApY1OVMl23NneGttqaTGx
K8vJ5+Me6Z1p3gTmYUxXNk61qp7QQZoKjsDI7hYiV8296sDX7AW3tdzJcmG+hbGEBq8Tt0OF2Y9k
nSJYefJRzzXELDPv71ZLosVlHdOWpt1QNLODw/tzxMDJc0weQHpGRmMEIvsOX2PYFN6BdMkwkY1j
/wVEpuPl94v/GXLThvmsEFx6wA4J9k71Ox3cfhWOcH++iDlXOU2SdMoYjfHVNW7Iuy8ZbhCpuR1x
CE1og8rh/fyAsGtrwHDunOGBd6gi+a41yIvvpAcjX2TSRnuQACI1rJ/2Whl2MBTO3QgAHEJWAQ1b
pHDPM4v5QgeX7xH4eVwkZPWwYCt6GPGtzlLavnsi4GTpELK+GapsZdSWvx8KF0qdlR5lhVJsgvYN
HN7gNY/mzcfc5J3iMyxdnggIg/gtly37Tp8WuVzJ7cP3QRWDdq2/Ilfa7mlruRd4YRMz1EdzyCxy
egiyqpPQUjTT0NwKRufINHT5Z4Ipa7nY3Gj05MJgyxafq/zUtsQDP2+phtL89s9ltXXyAccmKyFo
O+w94Hq1K8et+XOUAUXxV6d9bEVfqNu9ZVixN36YPtXs6mF43J3HAa4a6iIr3DpOUDZmktHK1rjV
uvMhej5fdD2HuzZ/ljHt07TaOM5EJ6AVmF8brjwod+A5pCHb7s30FxBlLxacX6mwUMwDbUgcDm+9
/xM/9BOtM2zysT1UDD5jsH7KV/TuTfF/7J/qS51pRezE4baEJn06c8bWrZRcsEr1Q3JyMC6kvMq4
2c2CrMfK20Tf+VDExROXIfX0EpnMwO9/IqCoe6amOrkBvH+N8fpc8E6Z5HLMghNMOBwnV40eLYN2
K2+TrpEg36ZOGlIex4khKQQStG87SmuUDGvl/9dttoJ5+dkRYX/Q/8VGWWRUlLe+4Nx5ghUEBVu+
GGnOxMZWURhy3lrW6BhXYqD16T2rwCdA4HNil3UMUgfIRCffJ82sYzCTslMxm7SjSgnwbJ+ckrm3
lnLawN/GelxvEqlfHRu/c6if3CeuLlj4Om1yVfkoThRl7hYA9gFgU9E19aoDVwdUBfa3TXWHc4/B
q/kgYDtySpvalObiIHHdxOAgxeBL7riOpAd6fPrO1p4y3BMJDJOeg7zKiFdDC8kQLqhpQ18lDef9
7Heo1pLUpfX6zz6jSe83LE+6J3Aj4qRtJaEcIPfN0MgTluE1l2d4R69ABkpbg/kbJ5IYnTtUFl/P
eFcRNlkE/WK3lBLEki0qmki/EdWOIM4R+nAw3dHq1NXowvwCwuvrdPKejlNDEI+ti4eGjddJsuDz
4wVwccqT8v0HnWPeYMvV9uSkNvkp9zrxrPb2UfAoZQxhgzz2GkfhpjHMaSKlRt41BYB+C6pMhY0h
K7+osLN1iuOJxSPPKAEnKp2TOgM9dkBH3L7OvHosGHkqeaK/vOZDydFPxiT2CXoR6EKuQF21jkoY
JyNGPHMry2sBSDoCjG9XHkvcs2n+ja+WMAw5/uOb47pa88XkrrbGT08Wi5X3O7SPy/YtkoEMY38V
OwjF+qkN5Xjpfdiz+xs/tYf+nXCCka4e6wTaQDGy7LUJhDYv1OsuVS/qVeBtFFaojWwWcLS+Tfle
7G8cZ6hSjl/5jYMOAK/8mg/k5k8MMgULTUT90ifaB9WQAqXdrxNVwV6mKyI4w9RHlI/0rWVvOMVT
7B1DTAjacV7HsTfj1uPYZTYNRLiWTYGWP2ydHiGefUtXIkAuHSldDGMvmKp28KOZicsAi+vOVag6
rG5QzTki5NQukKnwtMv7xt25UoXczTlR5LS26B3Kw4EB6Lfog/6oqkH7Wtqm/LI9YIfMSbw9medU
YngN41QXspwG4iBU5EfDxwwjohdc100SYUPHR8c+N0ZCnnSswUGcRchlD57sr9OeDTpXqfW7LhIM
NlQDaOLrGeQA5+cMRp9HHIlVxQm0jlqHfd/PojJjb5QPvzBxeQv9vaMRaUmWp/JwDbS1sfeiuEdl
gRB34Tzbo5gXbcCdyFdrELClfX+r18fnTOWV9+wLF/HHodq/0rKveN7VpxvGfTwpIkqtSi5Cf/g2
PUvybQ6wbBLHJ4HPtRZv5/b4y/b2YrUZ728RFXw8y99Jyp19L58CZOpz7qi5SnmVRxFrn21YC9lx
7g/rboP1bkzW63yeIMDCptudM7dMD52roziUgXRfDjseekglNjxVUA56H0yiaNcfINeRCtcXwxCz
ZYx8MFRMST/Kp+6RgzhN+ee7TXxbQ0YZNCVadcgv+PXpBt5q/3Vug4M31yDEjJs4uucyFikqbWUQ
wSlIjp8DpDEvUFxv8IeytyjVwpOuzOCx056CKxHkGWl+jUlTv5CWAOyIbb+AvmpMkPyzl0mCZrz6
MwIZnEbeHFO7+T6jfH+XeR+sztmsnQxjgRpO355XSguyb+xGYKM5NnI1RNwO94LGpIxbQQlhItGY
Kkqmvv6uIVA2bh+EnUaHc65oJf7FvhFVpuZesKlao+BdzAphSf1rTODEEv7gHEttTByGnGoT16KA
C17BLn6V3ifJJG235q/LTiaovtzRA2F7e7qCarcKn3bxhfXzci4o+DedUIG5la0XwLD0pPwvBhAn
93fL9wU4VJWLxrk4btdUJbgIt8INb8K/ejcfKTxvjqpZpX3aJUVVdJwvb6ZW0kCJG1WdlJsQdZab
BtJ877F22fCmxzZsDFVouMb1cWQhaEFJuTUeymhyJcjOzRcx7tWPJXBDZdWpimuj27CL8GuIZf6C
Dvzp1Za/UmtQA9jOkRf5KAx5ZhfzWf9tuE3YgY4oHfZ72Tt/pCVBlLx5sngFUs9igKiBUEwMosr0
TH3doid/itnjxwvjkj6MBYMVReT0qqh/ihQagGDau83/DPbbbG7Hnj/HBKSy8nS2zc5kymrzjmaR
+tWCV+s4s4KzlUzU2rv4AxDwQJWzrAZIVXfS1Nioze0kHxZNDca8lDy4Ss9AXcvqJc2Y9qQn3pD+
gNyEVK2lFlkDux2QNwlvqOVbXlosYSqqdsSoCduYob1AZ06bskb6KSiRVvIdeyTNo6kLJptBC3kP
UddEmslCDyw7ZrURli7QUiSH/EysuX1XsMTkhIXS5iqmCdae7nhjvHgF8WH2M5fAx4oKJMXskxE1
lHDyPOkuV5iec6OkM/okBHPRE2SRHXRYpHZeyxvvyHGDRvxpa6SNqdqQOP09ffjNCQbSj2S9ekvB
YN/LiwIXdzEdKzgT6yaYTLjCTH99URkSkaI4WSndDwWHL9YQS8oeWJcg1hEk4dj+4een3plmZlIP
o/wZUYTEBiR8rPqBtpwQT0XbzS5NVm/zyfWZN84W5B1yi5bPLoo/AUEVSIf8obwWNXUpdMPg3ICJ
t4opCwSMTrWUfNQQoanAT+ek+zqSYroLNdWdXQgm/vITkMAFMkk7m/NeWu1PY8R8iowkqc/EOkXK
/WNK4zB6wo79hx0PWXLFABbUi0UIOGK08V1Q5HKtnLmK9oV4NHjdz9TrUWW6cTRdCk/9eisjHw7b
Z1lmpbwAXnd3rE65ps+sEcH7S3y7s3xUiORY+ddat9fFuv+GTtpoZ1Vorx9VewyCMUzVVtZLdla6
g3QLfF08bJSq5kspyKzlZwqboZWfkNVT8YqQO8/e1hU7r3n81RdsxnfOwYhFo6k/ugdifd8E4/wi
gDV54bDTabpetyn1BMYOTSWm1ZTKrpSJFIvF/KfL5KcwMjPglkEkN3vx9U+lllpRUw5/dkR8EgQy
tZ+YD7NqdpJcHQkbTJv+e1x4kFBKGv5VxCmAARfTVvHYtADvpIh8iI6jZF4leM4I+HBLrZ4BtQ+a
aWDRrZ0nwfGXIkplPrxO40pVuecwb6Wq9sX77OoYbb9ui0UtH489jEEBRtzTdYh6i1ITrl+bUvcI
sQmdnZq4qCJOXyItOzHSRsqNh39cN+tjdBXCeJ4GtGNbWDPqw0F0Q8jnU/hLJUTLDQy80pEyop26
MVUaCDbagSpOAELNhgMXCHXn6KHjBFm26goqzg5onZON/6gJQB8wcyyyH9oqHZfy2Dol2OJJgzCD
T2l60jECfaRianGpZ0vfkSgEukqCpuNMpljki9iq5j4mrJGOgwcK/nP1e67NSr8ilAhXbRBBJr7s
8kHEbrgSlL6NmBx7YMbtRSqVIVLL/gEJLuw4e5wJT689U0MnUkOi+anAIXP2iSPh16OTXX6Cw1Br
tQwTL6aXXWvyfLjvJ2wJWPm2hBfUGv5DIatfs6ZrP8qEr78h2S5K+TMeAXYsWwjQO+czQInHFtk2
vcIDhmFSjI6FT53UE7uJT+e6k3P4gMegjjjMCtEp0aKmcuaQMKhiT77OYEeBy28y1EhwBKigmpaX
yPMDo6N8M0UFtZ8P63T4SNx2Vt6LZDGtF81lr1ALBQHe+Q3sR5w/pMadXZ1HDDpzWmNPrQMBmj9i
oKOSKToh9fOnCaAi/CxdaOHIrQFvhT0Z/QfvWHUyQ/T44jq9LbRQMTmsmRGFBU14KskzCCNTur4+
w+pQKqggizujdhgll3KDDyXcWOc7ryR3f6TnPrGYnEIFOl56MLan+hkvMLj88SPpPPYvZvXzgAsx
gM3pHnWi23oPOhNJvJMSmI0tIuoBQdzfAXAsrI3jDaTUVrIIPWXuHTT2jD7A3qum0zwclm5gVDrT
KZPZqdkkOU6H/mxylXq3ApkQk3ImKdLMINuNg4zWaTdLBKIeAH1JkYCu0pZBEGkI6k0zfXf74lDU
+GmSy8sx7O7b+OSGKz20Xfa7+Dai3dTsHWW6HdMbNgkT0/1WOAASzDGordLvEY71cUwz/Kcm63kR
MLeWTa5zGLD6RJIfuh/1awVHy7wos7iND7FVBBdcg/xkMHRL4iXApi6Bbz1VyvEYB8HkdVw62ohJ
t4KzRhMbZhqo+CW9Jdw7e9SNr6PInR4MfZpxQC8xPIfnA7asv4kCURHsEMIsbyCO8Tw7Z9ZApTtH
BLDnCrJbZdFdGIoOvxHTkuo1BRaQgnIc+oQuF2Tw974MEy5FnOx/aE4lTHczUGQq7kuwDUofgFNA
wXW/A9u6Yil03NnfJAfMIzFqx6r9k66oUasz0gjqEFBW8NFwZf2Zv8aZaYBkGMIzSnI2EIhqutlp
Ddgp81IxcrnoODd95RceWx300B3Mbin7vFH1KuJzT3a+EJ1hs31oakZ9vN5j2FT6Vp+vebYIkKKe
qbei9hNw0rFihNqJ37eSin/j3YZRZNARSy4t1hzYV7q0ZkSI8K3VbPnCmFM5UXKFWwx5GYspIFYA
znB/NOXcmBOkIVftS2A19kRAexZXEMBiBlBg53T4KUgeNxMYL/+pN+Esd+s2IFgjiLcbdY91AD+I
VNHdsfkmbToQdrUouoELllbF/fikiKZHPZt1RrK1TVnzDPkenpGsAZDFQXoxsa1gQ/CASEm0g5/v
Dyl75mwiCgx6UKUeje/UliY6ZMBiTJYCHEwKJbofrDukK7vbp9J4m/LhZ8Yqg4JROka2uGAd8yCz
u9HnJ7cRJwCJUda5MbY7tYAxo3NdkTYpsntMc44o28y8EWZt7TY5yk/Ecv8yULvwf0d2L+Y4iay+
idqQZHheUf7D49n3ON3soN2GSiYxJUT5sulAUDrMAp+o3/96+l4xLCwlNnegb9pPNwhXMF+0C+Ws
U2hhxWCYy6CI5sErDkJol/S1avhO/ekU+IzGeAlAQwFC4UlF6PWvXlAewPEaM0KZRgFSEzmr37ZK
2G7bOkqd2PyL3nGt6NPEIQn6RpQ3Qnq6QJy0tt0X73yGoSq4Wh/Z4hqVMW2FTOALtidJHaPEnnsU
LFfsk8Q6iHZEjuSNBkcvRGGtbjrssZ3yJfOB8wkZbgPmqzOh9Z+2AK1AFmz8g13ROQmZgbptRn8y
RNdUYs2Ovpcdd7mu8ABx2Yd5fd5tiB4tfFWHVOQLK1dIy3KOZRgNS99cPxx6N/DDM4gaVajhzCEV
cC4zx64Lo5hd0TKHy0F3YwZo/kigN28rRGd3l4VuXQ3RNxRfPkjKw+afyBjMBdqPKsyX/VPt4Glu
UTRLdMdXdDxMjim1Ah27kNL00Frmjb6yL0qd3GDUKV1+OBcxeG4BJKib1CiOL+o2ee4GVdvBNqEU
sfFnU4qhyl6BjpnFxJFL0FyBeAjLf6YUhlgxDmzUJ5LpR4usPcmKaeD3hzFRKtUvryCx0POasqqK
DY7NSIpUIBc4W+EW3kS3LiisVcR9Q8eSDQpMcxW7GCF9I/O9T774T3U1KMyGBcNrRte9ZqfXJ6F7
iBQiIE0+nXnN3araEuWP6evP8xAxt4eodXmlR8/uYW1DEUeVJjL9ays0COgTY8FSvhwcqQ7UWdDs
eGFvIHZlGnsRSc72gvnAen4qUUeWjiWAbg1jW2onG1Vxi9hbC3u8ipvG6iq2iT+2oZMYzaaYXTqY
NkQb1BzZPKBZ17+Vl5/8t7zy6p0alUBqwVPYxZfF09Ir7boS9JJERXe9Hv/My1tGVNyAmrXxr74W
voxUCqb6+ZZkDFl6vuK4ozJdusJUh75kBwNNTV+TA8aGJAzYuWoUKl9pFviaJ/ZbiseuxiGSL1EF
BdBcOgW1zwVf+BMbOfj9qRLDBEjMXjnVX9FapaT+6XeFeLI3mzQvc4Q/Y3QUyMgeITblImfAcYyU
19s76ezqHSwFbjWd/z5xIuf7QV5IKUKou2Qg4KxbwAz0P9IeSU8otqsZQPB5OzSc4aK8ZlTHdGyn
FR5H7m6dEtfP1nFDd3xbzqG/XlOdxVvcnre4AUYljiP3xJHIks72fDTauKXg3vUUskkHKnqDTgpV
7p0ORuXZcP8McGVtgFQPNRdpM7MqSo0B/BZMqn6ZuVOYG0OQypHOPlLxv9GYX5urgDcwFZ1Za+sF
pyHV6BAqy+7ZnawE6BPbeGZIR0fBeODMPPy1bc60wiAPTZ4ngWPFNsIq9YNQKTXvK0VY0hhbY362
t2nIl5uo2j9tsRA/DrT/2jqD74FAbIPM0O2O+7f0F/56kXSAOLKL7l/lACfD9a7nipfd6Gyqr0hF
b/QdbZerD3M75lh6IQBnK5+H/OoDtwe5U1/NhRI8rBfYMD77U096zTuCJ0yOJj32tLzRvFHZ0R1q
Xctv6hBxysfa/Q8Bw3GQf7o+76g2XpKGELWqej+nfxGHSsKJLSaYWEyOje8aYR7PDeOxbnDlIggC
rzkpLXOR7FHCGc9erQhl82krHDJMcz9pM53Tm6rEbFEloyf5s9nlgxjwjTsAydByGgPzr/S3uYaM
Cvl965Q/po27tuoHmNOhki/ylzw8mHKhl5VE75QnlPRowviqg7hXdRw10LdppxwNZkWM+VI5sdrh
Lfu1pK5A/QW2MudbFENpPj89aTw/PW1AOsxYoovwwnPdh7PKH28ItsL0axk2m7HwrhpGW8/pP2Wd
221uzxl8uDCJ443DVIPFzc37JM8CpzTV0hsYVmJxAr8NN2+Uu92d4ZAzlTzUIeJfSb4XBSojc4Ua
kWpVhOZ97EFpbCVdhK6tEU9BzxCG6q68RvWfk4UzRsSCYNWrWNrHUb4dISIwJCFb3dOzki3AQUuh
OiPAhjgJBT4lq+T51zqhP3KTRGZWtp1XAC8GLRZHSW/wI1xAR5CDSbj9wHOduNJXedKFbqxYkbu/
NZWgqX8XbbxZKa4dOMdBqXpvQY8LqqVlq3LiWRUsn+LFNBUBDjmo7ONcmspZy1yc9rkt2hKur1TY
Nr5vQamZInS6WRAXoSY9nLkzbZUbq3t99s9afNVoy1zbqO36ymi2Bzbje6W9MrBQtZT3g10ILVal
zSQ8msdOKpQeVnkaTefPQ0SD+6BEVjianBfslUVdUH4UmLf4pxlL7ihGCD0db96IgwmtuMIlIS62
NbkG7bVGzm7WjHO9a0GRsGqzONua1GBpgp8VSGjHqk97ivIUXUO+u1S5CnT9upZTW5UDgHCTtgGX
cZxdRcIFVybc7QDKA5R0DWy6nzgtfNkOWc2lgrcirIClQ6sXo7wtAtQvFA8qV6Mzu2zD+GveBY/O
IrrhBFQCTbQi8JVBHnVoCgpau7AaF37q3dLH1JsL9wKxhHdHPCOpl4kJx30NlDK82XGkt8wUaISq
wVohXjSdEoNk2JuHqv6oC9B93bX+CwaRS9Bud2jLysNS9CM3hzekvzPY1DXfOW6+6gk2F5FN+JAW
NmlRdIHVARJ40Mee0VW9mQpJuEtOymnEpxL50lqKYhzd4FHEFozQch8p1P6wgQ/N6wLQ2SMnOUWp
XDq9Hi6+HezFKrl+7McuTvxUdsKBXQyylJ82iPTWW6QkKSun2/BgkbT24GcNYEQOT0mFvRWhHZun
IyFz9dIzg6Zsp1pBNqWOuXOHMDbf8SYWOABUwKE6XwR+q8KzQlajnc+xuP+ewIJ8G0M7aFDIc6pX
DkYIcO5uW5nDmrp4lw9hxoTByshucDX5OkEr7L+ZQleRBlqjdLekv8gMIhURkJL/d99fnJ9gdWWI
9w05dQNO2KdDcOpwk4sd31dB/nhxG/OMlxSLnYEnnm0EnHC6VSZgKejAN1IRdPG/8Wx8tGBp0Bro
FaOrFrfylGUeNAGG58G29MoSz7ThiodGcwVdhLncQYQN5E8QfE+NpLWRPJuxsIaWOyHvVSFPDTKJ
TQN5NTxTzkcuSrroYOEE158HscO3UiRVCn7Z/Gh7OWxrr6UkBABAR1eIG3mkuYEerZh7obgMJ7TK
HDS+SVq0jY7Y6qQSV5Ffm2XL5fkXvsfRTQi9Xclxh5O+cwZtw1JjXEe1yUxsH9XaRyG+/XV0d3TP
azrv9SWmhFCEHOnvVatJrb6nxkxdcNU49kVrxbZtVBdCwh8CEPR1ooyDZOkaMiAJ6vo8QSDnt/NL
yt9+1UrOv7+LWz1sb/V8ypmXV24xGJvuu3yDxkODVEXPt3r9WBSWQzEoztEGF83yTmexJre25Vzs
0+eKp80aJyXJAf7ouGu3oTnY2fAorQ+mrCqm2zjG2GwadHUgxWg99FopZgG+qCofuikKJ08YwQpr
ebf1iFDbWYPNTehTo2Do5G163PhoOgTO/KXix81Y15EGx7Gs4gGrOjRpB3rSeLQvbrEhWhn9lQNw
DVJaCOEZm5BuztWN71qMvavyrZ0j8OgjORY8nrnktx3licCiEBk8Er81Tb5KC+YmHAfec0aguOLY
BzxnqF2tPb4Qk2FtyCezkMANubHShAn9lg5sMLm1EttwekzLdySZikC0RF1PwSNO7FJcaHtyOJ2W
wDD0UKBsq6yMQHWCxuhGsPLSrxgG6yNMOM7eYbI+P296Hbh8w8klFZZvrw51LqZWa2jpxGB5Xe+i
xh3nEX8W3Gr4ngz9W24K7EzUzhovr1286DvYQBu2SP7g4iaIqIQZNhiCeA2xB6SNKqfJ/7hnIsZv
XGm84xvW9gBsdRyoIZMLPx0MqOUgAgS0h5FJTklKLIB07tkb96AXkI9r75+Av5TsvB89UncVCeux
BPIqyAXH1D80GujlADNzdCE5Jo9E7YVCoSuI9zLcCfpdw8m5clefH4EKkGzVirH8XeVBrF0kDBRA
LdFxSzB0kUmZy3ybv+s3KWYkH4TeWf8Od1lmT/8FROevBytauMQqv6jYM8+wfITAiWwrq09J8yAm
R8Jmal4eOt8eG2wb1GMud/ulKuHebZgRFZOYcb4zTG8nr35IDw9OwuXQYkr3f5sF+Baet7ZBOrWQ
feAa6A0sX38L2yxdQ1H1DN+jl0MI1epYoB/fgsHdYWA5Li7LYNp8I7cDRXPc0B6tVO4Xkwfq3cjR
oK2ycyNz38DdDkFByIYfvuXHgnwPuKel4mce83fncYWRYUq9xzmKnPIAIAlnFKYBWqMhQ9HaH1ao
th31xt4tvCRkBmxov4uI7sKfJYGcRWCj4wYi5YD0040YaS094aOnr6Efqi7w9OAgI2ZC4sMmRhvj
6kQFh952UiAzKEQ3Bl419vW5FZi3sJOURjJT1Hw8kUnBccfk/r6pKUMmLN70NNZ3ZyHJsk/me9XW
vG04ORv8H0te6CmYqOJmk+NjQZwj4mGbqag3ADqV9HVVrQarboyJp3E51BTUxgAxKit2CiZwjkho
H7ka+Fi+ozsgq1/6FqlEaTD0Sj6dp9zKiNU3hJZt8LE7ls1g87KBf7o0KQ/iQoXxRuBDmiptjy1D
PJMu4QM+gjjmAQUQWlmN9BqK02R6TcVmWAcDrfZ3YTk50jUgFyJa2Io/vgS0XG2yAQoEz/m9w+Rz
/+WUOZxWLzIEE1OZ+UPe1sfiIhqq3hasA5eUeLLn0j3WGmpM+bUXsJKGBq8BqV0ba7d5rMlKgi9u
TJbTMA3cbo/Rwzk9e+kqxU5PJYP1ZnVolfLfqAy2uWz4Kbcngaz8/JwWCxeULyoWLBj/gE3QPezV
OJ863TTDChpRgRkY4OQoFK4L02nfygqJ9zb10ZivXaNdOrDrgqpKvHe2v7j0NJCftVQ0fxoE5OHx
qnCMbtOuyv85KLoxzoYqjkCT/jTZDjW719gLBKJWhVezq1SWzRuhez7WuQ02+KdrcaN4Aj2qEAYu
VkfwzVAR/L/mQ3cVqwqiywarkPGiNyavKvnkwjgiJ1Q6zJVxy52Eq/x4USnwuusIPbgyyECkEmz+
DdlOV74jO4BmuAF7sZvo3K7uEQVAAyyFCn+TaEkXJwBWsPD0Rpxj4c5d4WF3+/VUz0mTsaumISKr
ixmyPrXjjl+6fBd4LeJwzLetMwaGcUhc/TIuifF8GuZMYzRRzT5w4d1y74OToUJKOAsl2FHmOCq0
DEQSL9e8nGm6Cg+CNdxxue4Z0fI6y59qMvolyBA4pMFv1Szx3ENmZvmzwBZPczyduEQLoCLpbSt3
zQ8IahHewHsakE7Cj/8hzoHwxLK3o3Q9aVXuo7noNavlUUWBvuyjK/3xGaePolHtqgx1M3oFJADj
IEDh3185fUKRu4qbFcZWHuXDOTNbOwNsPWYhvhwUU4qddMJPvQ8yH+gYbH0FgPZndr0ooWNT7m+a
LbNqyPaviPVgbSm8GeaqrBlm8USNISKfa6nPftdJbr6dhQQgNp0XfmtgPVyipyPzoxmgktfAvyqb
T2VAlENoIC4DkacJ8H1FzF/ADoZ/WO35j+CY/8mZjbn5QhbWaK6+cAr0nlmILGDwPbzU2OwKrgKh
Qr94HMwA6stXImar/PZT9hGxse1UFbGiHeLkE1hGDajqqJP3BpNUdrevSD22o13p6mD76nxsl5F5
01sBztUqKb/v+4bYKT16KoVlwCByUH08ojnwAbpaiTKzrJ+khJdx1ewniVTDkJGoxIqfzk8VPdj8
xGVCYRUM2nXsjBDWiR/6bbQx055M2qAhy1x3r4WaP3ajpXRLpnxwhYS1Yo6DwDzFd/treZw3EURk
8OqljdbNbvh8qQHgDFEvDErgc1mMmR9bQKWGU7UWvg5Fq0w7Tv44u2AlQN/YqoGqgg8y8uYLYs3o
5e/bhje+hTHfOVYxm+ND6Y4fTk7zMgJ5ikhQfE/hMOILYATADF+QJFAjTjaZxB1RR+yl5JNX6wCo
ieTO1ymGmn0dGEC4jG0foXW6DwvT2rpAAKLFwIfCvAyjFiLrLewbnaA2Ezlrbc5bPeXDAZWlAcGk
8lEp0qKcvxEoBg9u0LPAxUsgIxnKWLeXOA0S0HJmrVA3vACinHkQoGc6vNxw+lTLfacrwtJia2dl
aSMHy/KAXBG7n8+886ZkCa3YCX4fpdOWOlvYEYlaPXiVDdJbWx9pv/q6eBEzuBMSskJCJz2917s7
LZq+uhBl5n37KJ1N3lxcV8Krh4epkB4vYe6StNjIYslJUVnO4zGF0b0quEGyqSAaYML3G96f0Zyl
Ra/m/vRUZ22+l16/T9CBsT9KScGnayq76RhHUcwe/K/XVFbATZLkYo2SPQgiTMJwb2fJ1YiC8UZr
p6f8eQkiV7AJHpWEdiYNAGvrT10LxpORWkMUDiMRAO80prfhQhbQQdQlvBTAvTcNwDfkfUvhvCQS
C3N597DAvL5hX9OSLyWYvtSIeJsDpSRzK7GkZ+M/ZuUBPCifM1YSTDd+eYFrNIQ7soRnATAtMObN
t+hE11EFDv8eQTESUhCF3ilR5RPpPVgP7uHNKahUM0jbPacCDK1OS0aMgpIl9i5B13hwCHIZinAq
Ux9G2RyO/YuJj6Sj07PtSdxlXIy6GlqO+6UJ/98xloqEelDYIR3UH35qvsoeMtKF5xMEKKSkYnyg
OeoE9BcLW9moTQQU6fAfmA4wQ8yIwTwuWS4W7Jj2t72pOMqTqACZvNi/IehNZKEyc+8DzcHQaHww
L2qikK4fd/pXRySxJhPmBFFFxKVjgE6tj7Nae7K1VaYWl+FOILoWvQUhJG316tJmoJW4kuC/e8eR
xt/0Khps1uVZt/xE+CzKXG56uFFzvV4AjSTB/VD9XBHfr9fmtTyxFbFA77eoMzs0SUBWHyDDDamI
TsBp0TfuCl+zN9LpIZtPqxHEv7TfECOUdaM1LGRRoZYUQAGKc96rLODI7GUFkxHyCWXIqLJcEUGm
MGaS5+a7OwVX3rV/+2cqFQj27x7pEDxae1mGUwfeq1ndDrkT66pwPPn/R1+JdTpnTOD3VXLyBXSS
y5vnQF+VZGYwif3QHWWFxLjlblYAM+9ONOmRb7OzOcm75/S4FE6Qr5FMxg6OcfnGz+tnYgfEqC7L
dMGPLZp4190/uu/aAxcCcNMrqi3rRiRKiIJCXqwNlSsceGs3ALTAf1mEHl4Ryk1QS3H9G/10POUQ
IQ2ion9uWmb/ma91sLNEG+bNTPNrvPw9kknyunX/w+EjMUfd3W8/2xv1LwF9nqDLtXiwFN1jI/Cw
pDIqj8d8kldskQJrtHtSGmpCSciu71xbc1KnfISPn8OkI7bKfmVqTDojNMNH4vFB5AJiK3aUXKfc
rlChKsC7wgm7xqm3lFIi35kjHfcOM2IkdBVN3DIIrW/wK6ThmFEWXC5biSn2A0xN+nqh0NhtK3xK
m8/NBgd+w+da+BvHJhiCqM0LzCG4lBMfjy/ZTh/8ASp1NolwXGzMUJjLsKwCtMbHVDk+ZjmnV/EC
F+sjhkJg03ZUQOVdq+rH7A3fcEDTrmgqdMBwzXzyfl+JVnZREWsGPJaOpb386J1L/hCjwLIMVfpJ
ACEWwIEOKTzP9xThBCbP1fFMrdVAJ5mhvXOmyTPZ6ynNNyIuv4DZLMTqq47u01IkNys1LWLI2W0+
Chj+jW5uUjR+msyaAXrew4E/+axwDwbYFi2RHB5j4wJWmlmZyTgnv3ZMtUn+BmWP7aMQyuKeXwu9
CZ/InLWrk67vzcWStNrC9C5eapeD0wTaC1jJhmZ8GaZTwYHhMJsBri2vFYtcvn3U2t45/3V/VeNF
rOAnRC9TLLhyDXP0otI0eqycoYcK8lgQIE/1uDFML+L8hcWQQwe7y84SSx8Y7FfBikMugtugdBb0
xvAdUeKGkFUlTvmAGNySydzA/I6g4lIng6L0/+Qvpf+wpXswI96qVxa7FfWNvXy34PbS0WJ7fe/j
LVobE8SdI8+4cEh98PgYn4Stqa/wHVpvkP2Jxaxa98pN36Jg2T7lLeBnv67cguGFEjkRCmvZ9/7w
WKSc2EnwsIuyGbmKhUJ4demNOQSJuWdKSzJzrkOJdD/rpQ1EqleJOHm0AiiDWdLu5QEzJLEzuvoG
zSRV2SWSUBRgcHj7AYHYOx1ZvapBsAtRyHObTHusmGOUmvd0ZPTOf+KyHPQpIC8Dv5vfYuFeCnlh
lqYyuJ3DwS7VW5ctxymBTf3q2fGUHm8i/Ae2L8I73kkHGkDQBr6KwZO+JCVcPyq0VMjXLsJ4tJ/t
XxrBnSgLbsaaDjnun+BelLBGEmntUVX04Uf73l77p/7dPsntLtl/D3P4ARAV0YF7bEVv1rn6YIzr
4v2TbKM/4BmbAZ0kz97saRLPdkFh4xqKIeCVRSzOeQ0Jl36yoRhYXX0xxgcl603oAmBreMGW6HCj
CVjasTFcnmKISBwyVrswDhel/LbwXSrn0DyZ/eHD9A55WVTbUde9jbssHcl6NJvdlmfoBATCFcQF
Ktr6uKAxg0D1EpFUgTUlEpaOCQRrKR5j6CRrE0fO8nQZlbc81Is2v61WaE4b3jV6NlmwTue9wOW1
IRMW2azUJrWJMFDHBWZiJXqHvpbk9iJ0Xrpm+1Y1NX1uR1MkIyXTPSeb3VTDspkqof3mZ+BQ09ZX
91xxts3gbSaF/GdwDzC7dVhuX4kJbdzGYFhJtrUgkHLBnLN6vpxHY+x+hZxbdJY850B1hm0EE1AW
tBlfpOmCa5G47O0GsTe4B1Qh1KeDWtcLHMVdbrLNYwO917m4gHo9d8T83h1x5cq0WjIYVT4Zeemu
CIbhJaA9uLB5JVMtMEf+f3pXlr5My4opoRAvluX5jx9JIQL3SWHuXIhoWjhzYcgC5u/NN3a91wOF
S7nwDgIR9JlW2/FE40r41fae3EBP1JQ6B8mlZsKbzfEBFgrfqkzvi/BQWTorsxERdZWsxUPippM5
W1KZbpxeMCwkdpqfmXbBUBvATR2qmLRX5U53XNM3xzOxNXdohYDQVxcCB/YSXsO0bRQm8V5XqZxT
IHgguqqdVAyD0UYDMqp/y92L+GWRYUNeVXiUjK581ceL5PrlKciE8kx+vWoVOe0rGQ3yMeDR4CgL
EZ89Zf8evLWF9dpDxsCIV0RyuP20SRql7f4wTCxlBu5oQEEKWRTRSFrTpopW2zHxZ+aSwJ062DR8
vvPjl4TDSUkJsuXHmxmRAPdbkK7z8RYX5TK0BtYhRSa6kzJjL3T3rAy5wZ4WHrSaNNE59MjsAroG
PbgsdntmNg+xlcEpEzEfgsCPj0A0HaoiEQVE0MAdUcoYG63o81f1m7c5dfpoYysNuPV6VcgG+FZM
OMjFlT6n68+C64Vu5rmljQc6Of3lcOfr/8Fqz0jitg62HxB9tBIuDkTralk8ZY9pYJpnJjnA81N9
W8x38qkET5cWg4amwwnZ4gwhi+l9f+gmCKMPrFf9Ds51VEikf65qo9sY3kFW1rVa31GM3KCwAha7
1V54oz7df1hMOuDWaWvztC+rENlUI6ms75FQguuQgirlvN6J2NldF2rpSPM6R+U4sHwQ9H52bUmN
8MjhO4Ybq1A9uEs42IUOz3ssuu9hWn5NNBOgJ1FNMgcXTwW01+SEUYKSzBTGH3MvLDPrItI4g2pu
cbTMJ7xqpxA6b7uVuLEu5W6kMl3iM0DGMyoEawoDHL3om/fDLD8ne59SCqzAmM8jcekw9K+/dhWH
izeoKd6F1HUEg+jJjM3ac5IViI0M1cDlvfzj9U7cXEAQ2PAmol0H5qNUesnxrmrGZi/wyo2S7S70
T40ssbXmhmN4hqFoAcvKsGW6USi2b0nT7pheJxzMFDcKaTuh0sT50axHLw1JiVpV4nVU4bAHunWv
7RCn3b8VTYr+t26SAcb/LPA9TSf5tLgicViUmbF7gNwNsY+EnNxCvhZBjLBdARSBPcCDvEkK8GOM
s65CDNlwpXL4R/3MSx20577ZJxXRaT3hsY/l/3KiJTPMjJ1z+U9fNy7R7jkWnW15ES56QRhibRjM
y+PqAjzq0hToHw0t0RHmpzE3DMj00AmucdWNTMuDv69pRrJzaBnFOaCw7mNV22+zXNG37AXosshQ
luX7FByFh5F82wf39vuE8E3TUoL7wNnG1g3k0MVZcuELNRcl30PIrsMbbVO4i1KzWsKrohpCOOPu
d7DDTRSiVUZuhsx+cHH/XgXAK7gAng6O7FS3JnU95BmJWKIeR9bdngt0xkyRMlvbn9r/YHEQA0R+
Lk6Jvaik4csiY4ELwBG8QmlYqa1Hce0TLg2XmsDy5SWNCw85tCCKcEeraM+EiSNOmH0LZrwSG/qy
9jwffKyaHtTINGmXQ2F6GOetbYveZYcBplta73xPi1BrLk7Dx4VwFkED3bfMkP+rPAbnYEh9krhA
CH1nKi4i4faBzzTbeoiVXnmIw4/oN/iSjc0AxEYS56+A7kIgsX3RDgg8N/TEjLr+f7KU4PjywBBl
XMyqNXo+RlAJ0t0inorAeX+QMXp65G/Vvbht6VdTHZSsfHaG9fOySrxfxeb0g7iVQ5jVPXEi+nyz
SHVYbwgAWS4nWYW017eWWPBcOKySRAjTR5L2niodCX2O5bxAn8CbX8suA1G7KwBTpS0Ey55ODhxd
2rIG/bc6ooc84Bq5WGnH6ftT9gBiQ/SIcO0snj817FhefA3o9/lIcDwYsUOtP2r0jKK5DxPFUxh7
t5Rm/iLnAaig9mauIesXPGwRF4oqpDtozNi69iJxtSYLGYhzwikJuktv65hG9wlgl0fqr1B9RjpJ
JjeheVpZChN3T5RBhKLIjrRtP95sdQN/u7pPWQio0H/zdRKdJMSgSCpHCFvOu4xtT2hR7UcFUCm3
lJ8bZbEpM444WZ3NFKZc2qhJUsmJVi+AW3Dlo+xTgZf3MZFgJIpAkoRSuQgiXG+4tdpcb1S2AK/U
oK3XtwPM3Ninr0xB9rmQpMRdcJY0fYpY7Zy7FvJ5fJ2ga8yJgH3qzK3tsvpWGW9UbiTcnwQVTLVm
985wopuHz/zbMKXIY9EPKt+z34F39d8OvmSW9K7Pv/jqGlHAos/7DwwUOyIRaDJDz8T1wT8NhxR2
K0A7n8mLW0PdMz82K3e/knAOIXw5o7plhJD5dxF788KFvKsEGkF34nz8a0CprWcHGGHu/fMcC2uw
VJ/LU8ilhset/+6uK45WC7gsD8jdDT7N6UkHg9he7IwPEXQY1HajJCQU+z9E4qO0pcZIgFbTHFX8
B0JUGJ5B1nDIuVvV8MYE/2DEoiEZ/Cw6/ozuEOPKSDX4kOGZBoTGiINKRxnLq5IJVPz2qdMl6HpM
j7kCEeEL0RWbHIVHTiXKXutP/iC1n3N7y6845C+CmA7tH+l9FsEACQcFB8EJIQcLdi0FvTY3E7d9
sqz8yt1mtn3v8x+F5pT1CwGxWXWJffY7EqaOiX0mWZBKDZSB27B9dJaHPMFWFikCc/hBto9tJBfa
LrdNV43vpca5DddAWGcEb7D1qpsH8jufHdstcpk6PtHPjiZOuPicqlcfdfTxOic8JiheKMDSDKSj
nXUMolq2/o+rE8HHgSWD/U55pIsEzbwb8nIBZnBjkcLWY1KdrTsoWscwuf2CvxAOKqY+eaSlKl5w
o65NU0wXIBbsS/rPEkWn+/2n3Gk+Ma4yOKvRDoTVvG5WIMXUc1YpDIiTmT4Jc0N0QzhFiddD6Co6
+omkdTboCIwhVLCOBVJBm0Pi4yFtV1ey55Wp9k1OdfD4+jk9AiltFfIY5FaWkpiVf7ZtEmp0hn7+
HY4cRij2vrmDP1IreDGjD6ASopoDjF2r8eKkvE4cgE3K0iQeSOwY+KOS5KwDqn84TD2gyfDCVkGQ
5cw3dtvsouh5H8rWw5/h76lqXcrGGzL42TMwr0bwQJCoFFwW8vO5JDjyR5w7qS59gnWMQYqHnONF
TrxHl1f9bGcvRwhfkhsWSS7YP1Ax++D/K6xKGkwgd8rCQ8drdpILsOGPnLVGbKzmJANr+ZN+R0UX
NLh4k/B4tNkms67+v8dfkosYnXQ/Q8hGNjEY4gDFkiNA6+HCEXd2xhOT3YXsRjTIf1ZKhkWQwIC1
XNBcRD+6IpUvx0cYFRT7sm3BjzfsJCl0mi3tbf1YnI9rEgyfe4G25tokSoUmAq2F86Qjm2i1r+FK
eTy7fOdWnZJJUvk28FnhZUJ0y7cr2dsxPXve856PI3HsP++AiBvFOteeHfIXRz8CUK7Y07HvwZ0C
ZyhH5I4DYFXMDJbJ0ESaGESkQhT+fkJVzs7RRwmBdMwJvoPzRGsCBdrpqNzZrsVgR1nGWPUq2tzH
ISm9ffoDbwqtSQOeJ7oJj92faxB1yQwOiDpZKOa4qT3vpvcP8T4cS62Q8vPcIVp4qA/e1IUVq5Si
wdRuP0MD8O+8KwYA0mXc/ueY8ukpQMjuNjkMU8zpLmAxyqRtUhW9yrR+1O9iU9mxD3+/k+YWW+rK
1o6PWAsNQBta1ax8fQEynFRX0nmQe1G9vDb7Qf5kj7mRnFcI7ALtUKTt3yR8VoIcM6F5ZyognUAt
kXNAjdddQjA/h5MVeLGd8vjBARSPTYlEvz+y3lU22t318NECqg8yPkDrqqo1on8zk0nk8JKshG04
+QZU+vgdEWvtG69xq3rYvIBe1pvduZuX6sxOxzfy4/qSpJb74i/+WiYLfKrOQgmJCt+9tVepcL5R
kU5pKiuCmR1/LahUXJ9Siy9MefiAoxAJAUMrRCLUolkL31BAxwFBUkj3dH76MvHr/GGCbORocM/k
vyK1Cm/EVuZx3/bUUT6On92/EzAvK3Cl9ROBT3V25GqnHTydfYzSZn9fV5HgPPOaGzogJoS5etPl
i7MdyONnE93QiLdZD9brZtCXov1d076DRE0Wj1UpQru8Zw8S5vSSDMAemRb17Ck27qnY/Z2TkyrB
vSsxGRWJcrlu09Ofc5wVTql8egODnh4BMQj9mQuM9/xIEERepgKeGh98YAvYSQnLjfYfW4Qb2QX2
mWOUUw9dnlixcugg3d2deHDL/c5CzCYAnf/N8DWKmi/JgiNhGrf1XtZa33zH0YM14K38p32n1ny6
R8JM4I9PRUrQun5273ghubg9reCHUiHNqKrKds12QglPe/5NcQ2ye/WVPTt9i0XK/Jmn3PGBbD4t
Gr7LhmnNbPx+YEJzVtXam9IOBQlXoYNp3IJZDlhaLJubultTtmcdyAT/h9CMM1jyERtUj0eNF9E7
Tfl6NxxeCpLt9Cybr6mWJv2xd8XJQXOY5k6I1ut3bzzksxMCubGxFwLaomMXAiq0gHjHl8PcgV3H
dDvZlC2K8oz6PoKuQ3ZMUY+m3EqcQ92WYXMJY/7qlDdla77yb9XDnS/yzE2oVGMqP/cSNsLu2VnV
hQusq2D/8AXROojOk2PwKvrtKImNvlHUfKu/GfLRDW2edbdyLGUtWE0R/atmJLFk4iGJGVGV7dTq
xPNpfTHfNR9bXOw5/Nc+4tYRAzXN0fWsiDki9NPHFn+cqSCJvZ4YCD6qfPnTAtQzXzcNvxYjxJFq
4qiWcD6Mhj++Dk7/Qf+de8RWOifjvXWbmXKXESxoi3huKos1NbG2ZbABDl79W78qqaYgzN4AuXuJ
1i9fExbEP21imrnc341hc2gfxAzk5NznAm4WUw6LgZur9A7KpVekINubcrbHARRuh7yeiCni1uhQ
6hHIlmlpelVhQph9OorAtR3A8gi9PdL58jAwiu8jCXKgvcmqSPuz1jBjYrPbduRZ2r8oDCSR8Atk
SCcAW+SEyDYWxp5bT43i/B+87KYyTDjCFNdHxlxqN3qFJbmPbbdhugvadNIJ+SycLRd/Vy1odkA3
YB/UGyKxAMvnT9jsgfvI+a0Gu81rhzeeRO7V9yKn5r7wuMBhSE4rQH9KiqJSu+HU+18OS5iOcXGI
ztzWsr4CHt59/QcET5Bb4iu87ZzeMkw1Oh7tnbUD0otzxVNJU/TeGzAhG4cxWIOQM+YcQxukZq0l
dE7WVOWhVp+LH31OeUsxeUNa3bL6VKlJacInIU4/xUmbo6/MEY9Q6weMCfn/gPOJTk3tTvlHmV3S
NQ0NE/5S1NYlokiR2TWRWVm+bjvnIUk/g8mWDI1ANwvU2I3VMuHFlsYLZjeaKFTFMRGrH68ttWI1
NHFjJXSy+b3MLwZGwT7jfJ+LE06wizFGq/gMnxTWYkZfDeQaXEmtd8cEIcMGtW3DxuKrnxvmddJa
yhwHqTaI6zNU6vbQ1zUnA8zXqMllhzLoYM84D2cAj/E65SQYND+EReA33BFzBzBY2j33wTqJ/n1g
pxtU1fS6UNprHspnfV78vdlRqmWDui9WyZwePcNa72+uO5nR1w6ArkDYFlkD67kP1QkwyxX5c3hE
/GrY6zj/G8YxK2kZoGBMEwy+eOTq1NQaV9/627d9p3c8RbgEyOXQFasgw+TRvAym4opIpfqjseBx
fGw7v5ZaA/Gis9zM1m8rKcK+3iFF36qQc7OpPV1HA0HeYVFBT6bh42RMmb1PbuEnrfucz9XdTDne
noWvXnP1uinUd/wgWuQEnHsiBRCMUOcol94Idp0ctrxXFeDlK+0hOfz2AGSHJ9UrlexeoJDTG5iZ
j8Vw8RHjdDHzohtBeavmtDwJhobrSWVbSrLL0EZd6XgYXgcfRo78/AC5aaR/KfL49euu0rOwb6kd
AHYQD8/SqhItyKMrMCA+Nf05g+xe5lb8Y8BFIJQ1hU5tFoKtIiJxSWoRhr5eEuHvPhi5YG47BZNe
zC8YZ0UPTc0TGRn60W2wA2YQsHd7QkPMZnNRn78mmtjqcOQLazPhIequqhgUlgsNuszQo1xq+Itp
146jr23IZWAMDzwqEJ1UlzLdAotkojM/UO2mBfSf2x7ri5Ey/mRZSkc1AYkvvsCEnATN3yXxTBlb
RYI0lbhXHkuMTp1P/R0o1Ghu3w3Eu/gnyshxz/SgZcFVTSCpUgEEzld+e+k4/2lJvSLyxu3xZp71
Fderr8msWwSspYALn8ZMgXqtm1mAt+RP1RpYOkmw9gamX8Ml6GnNvRYF9ho/E8brfCRtpitOXiUg
2e7yTql/I/MjrGalKSBV7YJwG703b05QXVesbBpsHVN41se3TsOTR/TgTGdIS3UZoWpcsTeVj1B/
nUzRjNPsWACJ7inEb3meEYuRkSMgEnRArqMHwZui83ER5qV557npXU9aRLjkoKRk+eXHpBDbT4kn
z74sxbVOLzpC0Pt2azF3wH9pPuKqpwIEnJreDzRUjjgElTMBdsu99a6KASNYn2r4/PfELLEYws9K
5vzU93KZxQ77jVOURsbpuOZqrkjdWhrO2b/kA0RXfz5f3mkKimcYFqN73oMDwB1cKdM9mWWfc57V
FdiLvt2PFMRO5ZlTju0UDvN29hEsQmuOkE9DPa904ZqwWjCN82yHZqXpf69JaigSbiQKGD13YMSd
aB9ay+rHu8HojsMiqbbxegTvqrp2Q3WMHYdNQDWAPT5Vqb2AvVLnn31EHoJ7NOhRVY1FHPN2qjQf
lpY3FIhgxOH++drtFJ0biJ8krlZ3WzAhmIw5PmmjPwlt9JDg1j7fv8Umvl/U2z6nn0Of1bN/CenC
XJ13nRJBiigoPem01LKrRcjj7bFCNtRjheYJk2CFGkTjlDV6OANRwze0TvKZgkOT0T7LU6VlaGDW
HfxJogKsnkajGpXkQFWKcLS5xOPR6UbdiQeKCHeyLNr+Ro5cTv7lQMqZHzy4YfBoNpllOarneRKM
/CKzNxt2idCcy5Qu64+wnoSHsvluQ6rk7aIwczl3Eo4lJ00j5R7bktLVfpa2iM1mUwwwuItTEmQ4
H8xi1fa8GLFMgFTmIXnDjF9jCFSQfC8hhY6IIQ+Ri2UpAgAmis2A6bAkaGawr/elV7UpptR9Vr0x
+ZAbmupWUJVCXHCgKMOzEFygbWHwAwPSK6BQBrOhyqZ8HDP+UdWM55ZK2WkiFevsPm4hFUm/drBB
bgq5UqVIs8rv6qbXw6sehHcePvCzamkgxA5PwZSQxqe9q+SLcqRHIzkKuHBKp4x5hoYv2KX5znY7
KD6bYu2vJhYzbgaI8/vKeju5j25XF8XvMXP7c37+/Fd95nR8XvESp/fx19uH1obc+yyoue+KkpP1
cKeLq9ciS159sTISIr7IzG9jO625ER4XnwC6WLdKvk/Md/+mHl27ia9ro+UYOUA8PBGU6SSChLKv
wwgaxMzGLlpovRhWZFSTBMCaHyGKi2NzcQNf2Ivpovn996qBWavQ4Tq03Su+4/zxPmek6iLEnB3y
xN0L8yuozUFuvcesxu0alhiVBVYzOTtw5lmhsjdVcg0Uq7RPdFX7kQu00iWBx8AXVjTK37YL825H
oWEday6nP3G3sl+dCun2qOHU1/1ZTejloiq8YgM5qxzDk4VqxO8AAy3VNHpCyr7UYIL6PhlgCsbC
zjqRtp24W6zvE1R/5/LqW3FLT4qML+He0VMklFqO5Su3piybG3e17mX8BBsnWnMuTJHfcWvglccT
eias11TPaI9EVPyz58ZJAD3j06v8rNxDSQ+16T7Il2cEmjIydHoKbVtX5sgc5cCs4A7hIYtCJ50V
KCVJotBuLXgQJTsAJONEuVh+7K0D5ubH7Ub5OVxMONpatkimIyRqc+YaqzsWcIRUpmlmt+Fbu7fv
l6nrdWFZGEBq+97dajaSm0IMe8TBEESirVC7jiD1rG3k8ran7JPeYl95oE+fBAp7VG3RgS2aj6F/
+HdklM8l5rHaNDP6xRuARyZq94GLRYdicqWj23Qf1mxZEDRs0ihfHIltVqIND4MJ7nLPGv2l2es4
tDqnxowDTjrqTyam708wZg4B7GP39XXjoKuacOhbTjNSp5Iai3FTTiw0nBDeGc7+47yEtBJ1kjWh
7QQ4I+2iVqK3QnyViVO+sC5S+kK2+6uluoIjYcX+kQ/ALAUBiFUkrTRrFQxPPxv9B3YatVNiPDQR
2aSyqYffqRJwYtJ7Vk2az4e9wxUFg33BIPLcuxOyVaYbLRIcQo0IjXmYxSXhqDJlQkJ+toVAdkJe
hM5Y/HZCvL3btnFU+aTpEfq2k0zTi2nAmYxHaVmwz1MWIU/Qa5xNjneITz1CIkjKpK8Oqqp3g+QB
5Fb7YaSsVx9KfMAfUFUDUqK3oOWIveYmdVyMy/x7a91+kRnr3gK4EDzuhzA+AS328niEfi2i9TK7
DWH/BOLpB3IxnkFsidNoCoVJuMGDqxVfiiwufKvH9T7uk4Cwf8z2MPn967TBKuG6Qd6FZbDivd88
NKEJBAcyiKta9M984AOfC0wfHNQN+QZEAkU5fSfA1PUTVpvzj7JwglScy229KD9k/VXluSsuLG1F
DsXNaxyP2Zp22VMSH2qujUSj62gFRS3UnKEAejRvh6DQ8cwSkX6uVEL+4QCcZTP/xaEODKQD1vTr
f2E9AlIC5/PyGQPOtOLcicTAMLV7SRIYvuAyascQEE3lBRMoMvRu1KV+nb627iM+T24SuovjuY08
UBgEReJNiWkMsBrsb89refqn27abBxjwFCz+X24bb/NbFg+68CvCt6yVSTkH47dzq4AjHkHtzeXk
Yf0c9CXTQ5XzvlDF7N0Nu6f1KTHAckOqgbSBdLF13EjhKsLLP1ayLI5Ms4IlShu0xdQfqorqFtUD
xyPom/kgf3FVcstFiTCHsICZcV3/kGB89tk2yLDHWGXa/9UmmG1pmMBGtT7npnH9jdSuwPHTc7Fg
+nkgE3iWiKrYMT2NKepNrguxORjNiS8AMM0yKS/wBcHQeywNawm7FKctVYHiM7ILG6kwf3z45Mwn
dTUcdVrCWlC8p1i8V0Ipa0IGTw8J6yB9sXRXMQA7h9Qj7LK312eLaV43d60K19TWyukch/pYOL+B
Zjx3CSgZwsYUyMhSahy0aiChB8ubHeYFpWkhKe+GrJMG3sF3+dXkuYVH6UTtwdNqSiizKy62BO01
jY3RuJ0TKthTXSh0L2MnZVMM+ShAFX7TW/UBi1iIIQPAGbgaJNewFb+E+SiDp4bLAn5fyaz4MvSF
U/wh0DNoExauNa4uMWyMGIzXpNL52IshOYVPxy+O5yj4/hPH1BpJB9BlJNyV1e2urtqIifTOdF0/
ZQDgNruLudMFEXASZMov2L+S6G1SFmyECNONWWZKX+rFw7trvcQT9gjlttWE6m7rW0knFtjLhXwO
PMtddbM357jne3SGu9GM2t8JYt98GhYXIM8cURSEyDJahn9hG7pgGKCEBIQUOvgqtevQKDHhtjbP
P/4Ubvetu9Drm7+k9vQQiD/LDSaxS/oHvqd55W5JTloDtUa7fGkudj+tyov1yseHtQvegNBFPuO7
HIoIiFVWlZ0z0PlxenLM4usUpSigfmdMLrD9yQSG3+kw0S7MUIjG4dlP0k3RK1YyDjadjgU+53e2
ihx9lnp+Pmz6minEom/ttBbZJQfREztOIs3wyefIE3Pjz/0krWpIxlNU2vN7VtoEWQB5rfVZ2bTc
+HD/ebYg66+EHqGBYEFg5xmR3cl9NQbEDHbfLAxWwwtAEbY+n8mk3WG9LzRzIlOfiI8CxL4y3LcV
8//MHl+ndFiCx0yw5oSNnaMXq4BCwcG6T7QuUcm2hiFbE//M+hUgdBakOR+La4oIG3Ka+PH9Xwo6
jk45T6TviNh1B3Jb4tfo3MnRtZGkGYBoPhp4znsWoce8OCmUAdU4Y6UiATFAPtQKcVR8QY/07QLe
meL1rsVnCn6kYTgMDGQjRyqFyWj71qCDfPevIZPa7mt3QdMhq3sbPAqFhhSkDPkYbpiXoS8afdPS
TEVAwulBNNK6ka/g6ipSMJYngpe7ndvH0NQiIxdNlazdj3u2QwnQTc1RQH5C7LwzdEGsrW1oxYc/
FB6pdDHfTrkEl53NZh+9n1o+Am81NvHuRNQxIw1QgRHz0YlOwo6UmWA8QJ02philiSlhmPPfV20s
vuLRQ7owISlgcuIWXOuSyI/u8maXkOhN3l79LmSXqTv8JsluBKeZD2YSO/gBPckuTmUKLaNy9NRG
dP0IChM0niNyZ7fA+mu5ht4f4PUqrFfk1u+6DO1z9a1sSlyFMWvSIpPeQ/u31FaWs7KZzmj+81Ey
IKLERfbk3wlizTHdHDMfExRFB5r9JfiUBjGQxX/TqjWRQM/Khm2vOdWNdDMhOhPZ0uGyoLxJx+lb
zZoFjtW95T7bNs1tQbvbAmpqX/TLOcAjBGxYz5dKR4r+z7K2/osEqzItYR8ATkygEKgVafbjsBIy
WNAh9z/+rkxXM1xT0jD6VqGAZgVXsyBXnAGwLklTY6J5J47dy/LLPA284DlK1B9dRpJ0r2VkvqxB
5VUm21tWx6eK3d9VYlzB9+9C8LMKX9jFPUedTFh5qUaaUSp+AB8/kVV4pFggscr+5+OYCzC1b5FP
Y+HTcV+ltkLqmu0Dqp4DJ/rWWvwgHE0uQ5pNpybMBjt/InQK8kJofGGYkdXIZr2xuEDuAEaLDVVb
CZgLDC5axNpSK9McQVDLtH/2ShtAI1V1NUnhpGEfUtuUQGDCjvGbIo4Ukqr/15phbm9Uug/vwYyT
tvXuEg0FUjexxunr+WbN1AhJNzUtBFdNuu/niP30tsy3/mRreon1Fa86H48b6tC1hK9nyOy/KJ2m
p/v0H0617qJx3/TTsCfCJv/plnta46Yv5HYQiRp0BORiz7wSkq35zMkTIJqeDD2ZBv2W77c9PWg4
0m4rpdTuF6LtYrlpKSjAblIu5sZ3/36MwELOF7hhKUdr3CGErdcNCuyv4zOXgFbJ6UXvrr2kC2bb
AUlAUTGF/+MnpS7/uYIXQCiRlt6R+9mT09NyvNUA+TSZTHK9VoM+rIHKPo3Z4d83tSSlXq8n+gKo
T5oeeUY4syEl5osZBRZCYkFk2PBToHUFrnr8NSgMZljpxq3gE7OGlRIwasJ4pOwnIPlOsEPByzgu
HNSk/iGOJroTRo/YinJNwVgvvZAxU0vQoBqdzOrV0cDIpUfGzSW3I+W93yaUvEYnNVSpWu8C1VnF
/Y65M50T+Bxws6VIcWECrlzCK8YwwwAkaCqzEjpo4DF7bUbbFDBlNJDmmGMd/lXDlxQo75qhtfT5
S2wcJmY0LKIPowailquGivHkyx1narsqhUoutuxJPCoA8IVjkpK1R8QaBGzQH2MCJnQHWcp21Im8
QV4Uq/aYnz6KDjjL1keNCD1k7kciiy0Z4xPPpy0xmSl6CPM/+gK42BkFAH+auMIrWL53F0nuW5w9
WL+QlDtRGeIaQmQvGZNA8MsEDKVRwiCkZLQZcI8/RGAVDzHbW+YM8IvalU3tCY9ePWvVFp01FGyW
eag0z0YvvcTQL9Vduu/emZBRzN1Q0ar03vjfS0lVOGM/cJrnGqwbfVLbvXYAQcVMPE2pN+zSGC01
RyhhhSgJqerJZgD7nShKaXm8cRhrBcazBiC/IBZAjurn/AiGOwNcT/Zgx0IjwiJQUH/CnvOX3klT
CvEeyV19NQyF0Y2XmEpLylIrH6p6KnbaEhenG953hn638MExHIMJ6IUskZbZTXTVtnPzjnieQDj+
ko5h+z8xhi3E1ghycNTCzNNJ1dgXmtiG62/YFDiHGZxjm2/SnIFmY1ohSZUN7ARo/ZJueGyykPPj
IP7GGWuOe3Xdzu5tWl7zQ59aOSOPYUROz+moQHs1dEtJ5PPKTBvwL+c1FneSGyuLmmBrcXJzTyMC
A9lqy1tE+Tk0cZGSpVK3Hgu3r4Pt2OJcUni54zWrrKAIaCFa/xQEb+GbuKKALujVe+EcgUhy+eq4
Fwx3WzH+QZfOtqBIMGDSsdffBvGdDNxKZ6dXMIT8ZPjsHTgm+GR0KuGs3HNFlIsj0Awp49+B5+0q
igfYWKl15Y5YWto16qE0ZAx9HkocpD0P+lGg23tTE1/QL5iL1HpGVFIDXW0Qz9Z5CsGlZOM7pmWk
wS4FXXeOB9KwpLWbxzIP12o6dv4YXb0fd5Ka6Jr5xHyPueCuaWgQfAOPLc1DuZcjUHpneKwnPe1o
nxKNwMZf64n0E5FUpvDN2z5roMIF6Tzl5L83g95CX9MPpVHZfgVKD8GL2UfzGfKrrkwwPM+228uD
u9lH4XWEKpWoRx8yL8BgUbFC8wTleFRMx7VsE+U5YL/QkeHG1kwtS3navbbSRXzxmbMlGugLY+C7
CITXfZE1Utu9owfsClXO/P599DC8SSifjkXzVKn+GzVdp4K5qOpAiB27acan6C92rX5z722MfW+A
/gbix0LVdvWepSv5YUv0sSFbBB4xGZ53GYUql1VaVDB1pJL4DRztSC6lKvq29Y5UBemGj9keN/GR
DZ4EZ00+LdERGhX/QLRy8ouyBLKJonOIL5WKccDj17KuqjECXIblqyOC/4C+yAd/oBxO7bJToiVM
csBtVlEy1x8CUGQZtN5cJ22uYmgiGczbEU499s6piNwm9qlQ+Xcwb1QcYTj43TFQGTTYm0sOlB9H
8QS51WLoaMIImUkCYIZzZQkgeahd6IK1lLLrDQyXiLCvp9lroMm/rtKOdVRkVpuLoy6EkLj10O7h
95H1cKzNry7XD1RV2+4HFMEBEB2R+Jf6k5xyJ5VZRZfdDPxO7GQdRT4AjjZCf8U7s1xnSHW98Yiu
Xwx4CKHuOkbzB0uOWx9KWAKmGvkzeS7Pe1uQ5suaiYTcrBAorBkoAanRjttCN6Fra3CKiLgCXMZN
OUxx6ODdzTvBcDkDExzn+iacGNxtPTvpO7QbHTHdhVwfS+lfstA5f58qlM4O0d5adRdXzggVxex6
7vf7wFvmCNADZ6ogfo+Gnjp+KPI6u7rYbN9L07boyDZoYpL1p6ZgarBJMMpLTnOftoNwqoBqsmyV
BG9APW4MMP3ySRlVOU91t0KJ6dWahVlX/7z6f9UqDOlsa0fOFiA+MHwdlecb+CMLLGaTU1Ir3DGW
YtfO1EL7G72nGVN2vg/upzlvzugKOG2BHF3pAt3Ce1yIPKfcdzgshKzsJmUZ5K4a4w1fD6KvP2a5
7WanbaLBetWcnZwP+Ofzv7BN78j7a57f/YCpkdz1/YB7hW6Ntz7CiRE+eyd2rKkGdcE1fZdbHlgx
LHcDmuM05EV+pJOHZJ5MScnGZjuiLfSP9FQ3ONRNVJe5oAmUIUwHdFb9VhRK8UjGJywUWunszv4m
t/mCn7c1duO19phMPjCq1Zy+zFk8O/7U3A2efxBI/j/fi64vAeq2xd93e8oFuG2AA8X8x6yQGH1H
H3F29fLkmiYw/0VYY4YVT/nxMvVy3TaoUCrpP1uLJG8W3LqBddlWBrbVScC75KlmkUf61tNcl4QP
nvlZyMoI3CnJ/zVx/MRykTAAmPBjki9PY/eB9LoFcN4HK/fBxeOiiN4Zu4HzqXEmmALFa9WwizRQ
4PcEkgn6LKgP3sBwFZm+7oMeGlVyj6K2ahaXa+FJSJSMlGKKmSm8+EbCeqyA/gF/DU7nKvmllUKl
8HvUL+wnFtnMrCXec+fkohyOHxMiA8JNVEnk8NrLu6Wc1cYrtnow9HcGFXGlDg/hf76u98PnL/BZ
YPCLutg8Q1my2DjtBhIufL5ZX5MVc+rxMWCzui0cM9SgE7Z9INumiioU8h55jgETT331+edF2yUi
4y2HFcvN7Hw3iZQYx269dBZIrYfxZMpwpNC8ZYzh8hYbvfIQ6U8I+MKopbNfSsOlettVv86CP3AD
1tjb08gT40cp9Qc22+j8M6W+yuDOB87rFlKZu2A1XMnbqAPWhbq9NXvCw4l5FkZ3g30JaBb7ilib
Lf3CKTVPSQFLS6A84/55AjPEQlRSmuuGWqRWg/Kf3fgdagx1ShyOGcsOXlTnVu2jqCcNz+iy4/3O
MhBjC+z4XrsaDPhIi72idR27YEpITwMJPtisUBqmJZnWfrYQhg28Sc5jA3w3gJTngT1b1T9zMqin
bSl9OJFFAsrx5ArUm6jnXw9QiIDvVMkgJPfeUvH81Ll6GqsAmbhGVzZ0pXmsheCxZZ7SS0wbqHmX
swrwPtflxCIk+GR0E+g0O2gcdGoXotMGzt40fWUEPgzfbCKVjMf142AQ05z1GHsVoOyN6FFj3vMv
lhj8nZuukjPx/DAqAFcMRAH3ozz8yksdq71P9najfl9tfc6zYmcSB/tgAk+6ziZegI/GpcIexQju
DytGgBFKEt24XgCV3GatXZa46OXqJoYNuWdaFUNG16zhJHxugcbF+I3ZWU+2JGC9Yu6egenqx7Nk
pMrSOXhEYc0J6NLD8Aiq3Ldqf6E11af+akW7s/VMk7PHgwSim5GeFy8zw0kJvngHvcnPVfU5A8b1
AXfzylOPouRqX81JwV3jKzPtJgpo4wdHCUaWbSRi939ew5mPs3SphGmLAY1iX3wcTCHTgrimhrI9
VS7eg7BoTmEMcYF9RfsQaJCQgB4f0c77faTuxToIRwxrnSbO9aJyoFDuFkaAZI2f8zYiShI3z0wM
NriQDK+k0FECT7M29qL6O4E3duRWsPjVFPWleKfxF6y/xdY15Ua9Xpoiuq+7depX1qe8XUvO390M
eJa2p/R3U5wAKXjB4cBIfl3ernMJ9LFVJ0//7bilVZ2cxYdZxrKheqQZoejOTzZpiNwJivW202W/
tioKExL/ELT9HfUHU/HCoGIWXU+RcjgxrNySdT3mv8v82MyH90Umf4CyjKy0QbwzbslhXabMiWLt
eAI6O9AwW+MjjPrMdgVHfvz2v1g8t2Aed1yZhUzrnQ4Jq4yZEqVKC5oBdE06HF5rrByIF/PPS/1F
Ra8NUsNNGUGhVeXkOZ881tRrba7xsXX/6J3pbtR0w8OyvChiu58fZd2qSJDFED0SNKe5V71oupwM
ltwHTsurjcY1uSZyotNn+o6mTCh5xlXOEE9YbxPBxHd3u5t0VrkS4uVkwsDr3h7I4Dzkysq4dkgj
9ytrVcaHBTVzRk6H3nfaoRyu2HwoWXe6lh5iR/A3PEglZG/qvSXKo6uY+dvDdv4NugwZEuMdm5Mr
fU40FLT0A8PDS4uKKwqYk+cc+Wv55yC14cwtyS7CXAb6bH3aJGXZiTv+pcB41XcaqsYY/VKknPyQ
nrSadE11egVs44AmhjkWHLeB7ziuDDQsQYbiFc4h2gNIU9n+YBWOy2jfUMYS8TEa87udVWOg7uh3
MlveciDPdaLgqbo6+BA9XXDf/gDiwvoyYtqDYhx2bpZ0+zTl/MT35+zBzTLJ/kvCDGRv1mq5IiFo
0UxE2PfXZrys19sYalP9GqeS3DkY0ik8d2C5TADulzN6DnE7exjbWKFHfIiS/innUY+Oe9NMW1w+
YZ9T6qalUtuJZO/PWYJ9zXi5LvD0/vrw597lXz36hQDWYcWtsVy5f+ZPLSA0cCEISM45OMLlILsz
rfJjTJAjD6k4mOOHP+lrfe5ccQCMYevb6O5HGRZ/aE66swlsyDDSpE2WTEcbNt2iGL5O8oNAFSne
xvWL2NaCVEmpn9M9pUhzX/szJuPG4SH1FvKN0lnmiUPpFgnd7uZRmCdf3f/tV1E3KO71fsGd7iny
2hU6GSWGkK+/ykIxxOJFl1zBeZ44MdHXC/gg2X7CgS/99VFaLpqGK5jXCB1xPnwG04wsAtEE7ubX
iFAXGh0HgFCBBBGLhQDFEbHULjaDdTqTXdXv5jpKSMzfTZVV72O4Lmq76aMDpJsKDsW1C4Q0Y0oV
/SJnD4x7TqhGYzp5Kjl3VDlx04GA6cMWyuzMqbVO6I5l5ch14T90lANLf14pe9Fu0MFsK33SKFed
Mk5T6dnltZvW7uhCPsMgnrtgXdTLtnH+akpkyD84N7ICGMnihXa1AVBPlJ643/kUdmZj021zhP/Q
WHPryb9ER9JOImm452p1C47DKRTYBPx53ShOTfbpZM8q9UAqF+EI5jD9uGd2L25T8QMIZOaXP+WI
8iof95jtyC5Zjrza4ugxPgC07g6VMzyYes9GpOBe33Fuy/gC7+MwZteqm9L8pHjk90Spwb22e0ry
ok6nBmwt8uA12z3D0qu3XVrkmHTU8O5uGKqG5svxHjusMI5YaXthBvoF/W8FrHrIMDN2GNzKBLWl
CPM8XjiS7HJTE3tSxHKgQlMAPKdovwmeHI2vB6fbho1JHKeBNR8O6ND/AwtiZL/MV6Cwsfh3KEzz
WhgC0HmEbd591MgaBud1vDeh8JsGJSzkJtlmIs5qne6Ifi9GQTZIAJL6fxmmwpMsZwoormnCLYOX
yTdzS2s35MlmmIi5fG7f5yZOwohSRDXgjI3j/ji0vXzFg9PiHOLJ1jDlTbBVXO75OR/ML0UFmght
9S8so/MUPrTLri6pUtw/ib1qw6uQUobReeJM7n8TXJnE4LLEhK8JTTBA95VVREEM0wkTCk/RWyCv
szWB/dKDw5JZjYINagvOeoODIpbERh07LdyipvDh/v8heMQCov11LLzQb/MMYeRsYzqQ8mPbEqes
dETpphbDxV240LhSYCDc2c8L6ZAZs3rvyqX9G26sIvnXP8e02njtTLd3uIN2TxA8I/h6P/ozhDyB
22EiNVHs2/WlskWcwwS2CGLGRGzF93v1hHEvjVjRiMDG98GO33vMQ3U5olnLupDcFyKiREpmnQvN
dgrJsYC6YByoM3cLG8SixVSBFlMb/HTqWR6mxt0eB5uC4MUALbIrR4TnJyThcI+McwszqkQwzHfY
4ErqmXRrzf2K521CXaAxEjpgIkK5N1fVx53OLzHQI0Y2lwKc44MzIoK2iRkbPmbFTkt1ybxm7qnh
YD9A8BY2uEJcNBLroxlWPm0ANCjVKnQjtqZ99j3FSBaTrDxXTv+AyvwyvwoCAy95ZKD+9SqyQQuQ
VyCqZ0sR0LAf1VqvPHS1g7ynZe0MDnyZRoLDN3H2q1IStIUdW0r2BcEz3CKeFU57JmwmM53Sb/q3
uKBH6okZ6nltUNvKiNHoTFhWLqP+CojmYW9ogHQOx2DjIfKTElm0jcUe/10+uOOgBTa0Sk4B7lU3
HCTUlJHroKDPcVKt1MXGYSpsNHII4dNdfyA0xoFOA14EZZUE+BucBxjPCK5DS0t6wVmNcNih7aaP
O4siqVlVcAL6uEoQML+ofnrB6zuXyq12MgAvCgu2rB/hUeaBX5Dfva0jM/FWpORTRzUmQ/ld9cc0
5JymMgRr1o4q7eU7fcCZPKVnEnVFnocJWYc68aCj/gXE73+uO6NEvXDmUht6NXwnT/fVeTgux18j
79FuCLzlK0rVU+b/2KQXyO+jmBF82EUr8wW6vJBERH/6/IvpDQ/LUdAZ2MX1tSUpWPcLpRnoCURo
seS4TkuY7RiO2CrSexWR8Eq12tfWlrRO297htJdkIhC9ukBb6eNjY4nMBjhzxMWM5AB/31Je+beT
VfLLXMBxQxBkeZYRe1MP/aYMxwoRKpx1xct5f/PMFDDZw0cRRcgHlO1Mt7xOvzxX0LYYjvuFILqZ
SnAYxF4ZN8pW3wHMWUuY/jJ9XMBcc++so7Bf3VOLo54E3wK98CzERVuReY2i51DEA1mITcdcuqun
0IBrWlP87bC+E7xHyX86Q9cZjkNAFPYMmBiGRjS5MnE3xqfTO1kMWDkCQsNGWjSrNhf51Xp7RoHx
A9U1t1Lm2fN9OS5C4GHlgvgyf3PdyQ5sOc/Y3xewIZKcc98CsriyM5cfOarRpazUtLtviYPejOQI
Imwavc1jP61WalNU4113M+nrz4sjh+VRtZELkWfl5gco6dkU1GKoMlDtjlxI1clpa9N3NzvSLKR7
c2X6cVI3a+bf12LGXZpImHGaDklx2plr96YmjfGCxNRSWQ3STyc5TsNEdZM01WrA9tCr0qCSwd+O
PY+VpwsqICZ8Ai1+M6ivH3wNOThAEktEB2byyoYf6noVqOHXAOlEsGtwQT6wNN8G+Z2B082QEL7S
GBlXR8IFqs1u6Fa2GvDMizM/BCk22TqCX29NoA3QbyChQy1Zu0W/rjXrzkR7vbO9kzLorSDYsam9
Va4V6Ivs0L5vdravYZdgQfhYjsLr8pCtEQ3oAJ2hgJ8Bw5jDi0t9r2nWd9PSH9N/bRs8OeGxYblv
g5PsW4vxQeDJIGvU6IA38Bvuqov69JnaRfBc5yz2U399cNbXeX07gWPtkqafQ85o69/pFTY+PcFf
WdPIbpY6myRf1ox+4nweZCMWq3y8XK0XnWx35H7kTYrHMDrDh6sfVKYyE7mXSyv29viv/5BDv+Tk
jmxPdBUFLHixow/ANcwKDNzTfR8AxOXO8nlJR9sMwEjaJHLC7+EE7Cv0JxfORF4pver8wamyAVwb
s6c5bTKzwlW/6IFuuoqxM0BJwLBcUMc1SQQQ/3wWjPY2IxM5Q8w29ui9vSz1RKiBOzm8Y/tN1alz
qI7fir5wOzXCLvii1gYJm6v0djJ8xBKav5bsknl+81XZCCdOIdssbOMMDj1dJcElgbB8v5iI3wwC
/qBZpEysiFP616fq4RZGAI0rUCRUab24qLnG/BiwwG915LQc130R+cUGOjwNHmODI6jUNd8+wiva
24g4rfJugyLmt+cLHIehBlYrNXz769K4b1Z0kHiB+4yLOhzY5cgqggZL8co+WjgQTOF8p+5lv9IX
Is4WeK6FIfWR+lIEdpgMymmmJkvPja96xkJBgWs1KFGMbi5tVp2crvISCWnfu1PeK8HskghNjDyo
xwdQ0ZODj8D+OdTj0n694xvAlh3EcLSi/2G5BD1kHmPfARzcRO31njUaDnr124dGB1IeihDsfzXI
6YIA4RnLFWNsDjwN22tkKO5MugmH25F1jD0i521NuOzgr/VTcBzhReMUPJsKl7o/AOa8DAjkDV/Z
cfMt/VzZwDuOCut+N2G/KxJJfPQV9xAuD1DDWXxx0ybcmmnFv7jB7MqBeMALFswMgL22how/4nB9
dHvkJ73fksQQGIIS5wB+02d/bjXwt/ooWbU765FcuXojXXj3AJTVjNbAY73vHELgjioYRPsR7Oyh
DM4k4n4uBACHLf55md+z/UR+M/uiYl9/P8hYmJE55xpfnbBPDqZ6UQMKa9VABYtUIpNlPktj1oJU
vvxQ0/tl4ubfD/YDh0fhZIbo0QNtg/Lw7vFLSIwxWy5fTq8jHRA8ioHo6DKA9mZwCfDGNwfez5Qj
+rAWnnROEvF1P0j8kjr+n3t3IpbDthYuSUo5GtyK3S1Mu/Fb8w4+u6PNXR5slcpDq7OiiDP6Cg7k
Fo65l+DoG/8oPjrtvctmxIEsqwqS5hnzpH0MHj1LzZJ3GIETt8sMSODJG2QE8e5E7oq0ixE/HPjD
GaA+Q9tsxflV5fzCnSxa7iIK2H8q1MwVe+A3ko4mQukQEdsZgaCCLIdE1UmB84eRtojV1a7o33JW
3WpNxbAwb1dLUd6w6mxAvk0bbjz0Cuxbpo3gWz5vnP9NUyi0lxZk4qYNUxFaXOXVSRLCcSYYhb71
+kYHGQEXiTj/HgI4waJKDf2O7n+wJordvMwF/v/GtODyOPgWy1Sn9ydB2OlaKPRKkVmGZ7YuzEv0
e1zxScSqSsRu7jKehckd1LB+Wh+kzRlM/B30f6yIHPFGtkrYsmJOttfeHixSOm5NU1+ilRyRhKQg
pH0NcTlIvr8y6Y4GjitsMv+8R2V7zOx4GCj3stRGqVezcpJvpHifSypLTpW5mJCggGVigPVKgReO
aOvf9p5JqDcj9W1dGG/6DTc7p1lQojMT5HGLNCqbFl7PqHaWCjwHTT/JIAG/aRgz4SJEbuiIPeRi
/smr4gtI9wOSq2Q5Kads1CSthtx99ppOaSoT/nr/Ogo7cWXv7lE1jm6W+oLgVXTEmknk2vK6Dkeb
5Mjma9HvzS3AZFkT0/wIzGepbIRwqGePd3RcIoBNQ1vmsVfOeMSeNKYCWZpKngCUBMVlW/yZiaiv
nC/SQlh9edAZdVeHcZWHD+XyNnFAaWkSrI13kL/+h5I1r27UwYKYW0wJIRCZ3tFyIMyl34Qyt47V
X/rDb5w/Pcqubt+7eIoNwTPDsRHt1k4eNPOM1IjbZPsbCJUMWpbcdujyhMSD66rjbx0sC//7VI9t
ll0lFw2T/WGbfNt6lQKss7tcd1weQEvBwVWBuZ+4i+CXx9p7m2GkhXncq0yHjooqseH42YbbxGrx
2lQWOqdHuwo/fpwDxYecEZFQ6iaNFXoPGL5/Pqbttrphx4VLQOumccOfBIt/0dV9P+zxZim5xXuF
MRFwGRdDO0OdORRV6Tyr0ULN/jduRYY2alXRWYurfWqilMS8D1jUcFBcm5xWf+semsBTI/qOUO2i
wUSn7oldA3VY7wPjt205C8NZXGMkv9b7R29hbDYHb6sR072T0uLEBA/9KkNWobSDtkp/GpbnEree
QUGI5w6otpmrhDlm71S5OHuKko7jPJQKbhFEr6913qk8E2yKcr+XEyiW6JyXrO5X1GkUKe+bg8jt
ZNwig2/U33WWGHDZcj7b2oVrOTi4pR7B2thzlwRM909nXCAZMRKQmR9mO+hdy83iA7LuixLHqxUS
yhGR3rIrrqZ/utB/MwybH7xXN9paIgOUmhWyMEbIyyY6p0dWwQxwMs9kzuYTtDOG38rH72g9fEs5
9yJ075dTM8adv3tVBAqRYOFZma0OaSNgKIL+TBnJ6FejfM89+Jr0Jz8QNtuXYuKp1ryJKepMGm7X
fhj8JjJ/7ufM3gdRV/wn7Uwv9mnp+aS3r99ghpLPfPX0HwsnIpS7Y6zi8nEUY980DR12DPOokf4d
czDx25u0G1FJDyKoG0m8OYi2ACk9clfM/9R193rjMDhgge7wH2tM9Zp1Q17EfhqRMWHOT2l16kDd
FTnMx6v1O9k2KpojJA51+gzey4yreahHrvXdLkp1XBPuEXYFuINzp8OGIS3jfHwUhU0u+tTylDgl
97W2GFSNvxKFOvf2yy+/eY+/MceZ5sV8NhbO9deAKRVRfEvFZV1QCE/Bc05BXg3B1YpiXc3KsxUP
pQPCBGbiqi9rEEnmJYIzSDuLXRnDPsmsm+EOw7Z1NAE4UsFJ4Vhj555UzoajnXWIIUOLtx3k8qFJ
6PyrtSaqZSwx68n5gThD0lQbPGtKZw6iQlxlC/Gg3UisfkJ8eeJ9YFeYqLMTBmco30aETMXrT6zq
r8zGp4+/N7zgIgCj++IP+kDIRGc3T1n71EKwisyqIvhsdOGW9l6bcog4laJPqp+NGgBjXZBrdI+G
I3sSFvYFtGxlvSwykTZklcKEvwj13PVgAt+fHFORaSCEJ5/KaKOvMDcUEBcZPDct9x4mf0RX0wGc
f2uj/4azP0UvmAUTOYwTy8FNWPBiCkLTacpCh9/pTZYbvzrMOlYe+7nJIVEPdpz3iW6t3Uhvhji1
Zt+3Hk+xxRah/fkh84Qe66URj7FpQJtsiUmuDWCfP7Zdx05ID9lFGYdiDclzUAx/MVJniiTzDM+A
si0s1Vgslbq5d3fYCBUoADEgbXZayw6IDn/whiu96MO7TwcfnU7pc8QeV39tmQo2iCqLhRJi2Qsq
8iS9ecliQYlRWc2/+BjhJrrzbrso41TdrtWBLA8TwgtEee9LVm1k0TRs0DvX6WCgT/2nh1W+zBvj
2GTgkA0dmH/zd82Gw3jFa6yTtfcjo24e4+JTXStA4R2PR0oYGYaA3VuONi5WgA5yukrNB6RJZi1o
+GZO7+U+C9m5zfwJZ7qC4rEDwczOoef1JC54h5/IsaWFqYAXzPszyob2iTe0SG778+dIfT7iZPA/
y20azH4ETuTDL340q2JmZCBTH/8KZrOwwAMtD9S903kc6yWRMT2vt4JNSSLnlDRVG5xrw98l8uO3
5oDtdKVgpjprB53aNCDTyIugpFwJp9b6+HbZ6MKowNa4oF/IZYK6yOcfJSs9bybqBsj6dS0VLdzd
VcuhxJ9uxKO3Ul287k8MCKwEOOR1F6QCKNJYmx1P2UChXK6r3BxVgDy6YLHTm2gY9HcWSQ+vQpt0
3DnrmtIgtv04ymfUZpK8L8Xa29ucFLmVDFekO9zH5UD3Hx2a8Ns52pX/chqW0GCmFN4RtKdlq+eb
O9HUNKLIgtPUcd9pykOhsu4uTQGGWP6E3OnTfyL9RUkjX4P3AofodCQ2qlkVDOLbFQvNHS/elp5p
pX4c2YX5r6qAlvZWwwVxRZtwYBryhUJKciponH4PDlPCg/9uqRA4Q5FU6Jfoj0bygyDY81NEYSms
p00lufujrkmcPye5+n6qLrWmC7D9fEhfw/incBhPNtj+6JzcUxR5+Ynl10hNeSWpyVT2OnItcw5X
PbbipYLrhjYOU7uJ6wNnyBLEVLAx8Y47YfOKcZ3Wk/JKWAVpTNNG2R/E76Xsw9gv2YyL06/gsMdJ
ubv5zKA5Zsv66OmiMxKRtMLKUiwqCqhdra9DlOv8Cv702Af6z98FnETHpMNgVSRn0fIcoc8jo4ij
FyDtpc64K+ZduJUGMWGzJ2zopK3zMYA2nfCEW8FH7sYpVdGCznhCdAN+peMfH6UiLdLl/SKUUeaW
6jtxYhBDdUVMVas/o1R30CdPN5wTYkEGUe7hU8PZdG36bvkO9y84YN6NxiVXtocy4YIaToXukulN
Y/dpUZxNHsINnJ2qmvzh5nVKRhYenfRyor4wvZIJpf2MmTfg4H6sI77vIX+DBvNvW2hAT6wdYV6Z
dOPEis9c503g0o2dKrgRG5XEG7BP04MBw6j88vCpvCFo2GgsVVMnc45aL4pQWnK5Ghgu1n5t/7yc
MBiHsrHE5MAXsTst6StuHR7SmqNpd8VMTzx5gvv8W4X5G4bGl3wgzr5XnrBP+s4PAFmfkndFQuAO
qLNijtzIepnz+QSajS4i+ETsgjd9hYkzR13zeegqnwMyBFkv5mH1d9tmotghomfXdVeWpV8SXuI4
8OKJyNxp4wPoEzirTVjye7krEze6cRc1x/dSdDYFvcJJXFyR/dohDdBKo4rb0HvG4Bz8EYRupVKb
wUGw4IObMF52XOk14C3iUTB6u5CzFm+GKZY4ambkAJMBkrYuuNULNrwX2s5JAcb9svc9vWj9rVK6
u+BWA331siqiGTwU7bs3P6ilGcG4IpRe5EtdPJPMe2tzfpPl1tO3k8Fb56mOhK/9PPL9iqkvborc
RmUMuUXxNmKe5C+45mVeota0wIP/WQCiKuPN2gvRgIPX7SVqa7GA0y6VzpPGR/OkFpcRAeJc8soV
/QdgrABjxo29jXiDjYcGR292xsNgOj8/Tv7qkyRyWseETvXMlg3ziHylLYEpouQCXcyP3mK18UMq
o5PCEo70tG+Bgrx0Ew65YwykzET7UjWmKBkTer2Ogv/dHs939amSfLrYcmTNezrffO1D4FI1ocHy
c7PvsjLenSZKpXGQDH6mb0tjqXeP8a+jQ1uB61jt+hY0LJKzgY0GVzRgcB7lib4mIC493mS7hi+Y
58ZgbUn1OOicFzVrsPC10W3tKRqtpgx6FBaaCiftYSxVbqzhLto03iasjebUen+ums7EqJjAMtQT
UnipMgYAvKFGDzvRzXAaTjDl5/m/QuaUNIAdtGgS/bPghsK+GDiuGlJCQF/ezTnrtfuVnBLds1wk
wz49tpZTw6zEIyVddUIosz1bIEgHLhadZRaEDfdIL01GzaI5HtryK8NgC2RMMX7L13TDRNSdZWSq
aHm34TIGjo2F9S+FIHFHrOfBsQo3bPcIuI5zDOheeiM9shP6LH22eeEJCrd34VcwrdpajpIHs6Ur
jUcGJ/Wd5u1KFldFMx+UyMes7o1DaKJsF+6qYaDHyyhgIhhVLzyuI/3ZGTbjlcnJPpWRAYNM+cfl
+PqizG4IkwMSD/vC6+Ru0fkuq4EmaziNLdAPUYSwcglfolsUKLcCI5AG4CMhzmVFI5I3+H5fCbDW
6Y2clNSnNSYMkAI+RsbMFdnAlIJQhn4UjPG10T6yRmgdwdlIRFCqA3zaYkdTJaSnb0lelDAQfDuh
qmsqURuQ7i5C6kkY59ueVV8w+Q9fvRkPyER/VEcjdreuM0GkLD6G3z1yFwS6WrGlTgAlKkaRatMA
tTa2fZxHIdGX56z8dcVOcWvNBHV9hmN/EcAphWtRFaSE3bYJn7y/KscL94HMMgaF3ACeQ9hheWap
Wfm7G0RGWdVbxI/A1ZfDT89ga+6FddhrcYk0yjsweKFCqoOrC6iuAGxOjxrXhQQ//1PMvxvOBsN6
3VytRmQesGlwv2ZrTf8bzmjd2FDyUawY12FzvU3alRTLzJmLVgl8dqoPt72JUr6G7JPZQtzcFiJv
3UAtvuO9eJJQ+eZvhPqZWtapMPsSHg8LvL+jFcf0YDZf8sWFfXq/dgbInPSABziyDGo0VyT/PGhQ
qBTQs5cL2v5omGVe9+nB+dgcUaq6J2DwdTxIkXvb1Oo8PmSZrLjvgauTcOqNT7d4we96S7NuSsF0
bRe2Zqtyj7hQy+FvL9eKq54b5np6OyhQWqGA8I/+LWdcYArjYRjUyk3lGLBC31PFv6RzgKH+Gbnz
CzvCfvIEe/B39CvpJ5Cn3N8QXiHSO84RQtV5jwibFsO6kqim96+HJNzN+8EK9gXBJ8Lrwl1Hw+D6
cqxfJWDBQx2Gd0G2yKBOYJwK8d/WXdm0tIZkYD8tbzxKWnJpnW9HSDMP+kfN9QVt5a7gsIu7K/pT
QbKDvZ2mlS5C1ZAK4OK8YHSr/fhYari1g4Qn5BKFwK5ABlHf054wqluU29RLm1SlJigcWuTGv8/s
b9mzASK1aorcBG1ltfnErnzf7hPU/8129PxFqSpAV93+Zj8vnnfLOle/L7XCFeztZyJzbJpV3KkF
eTorOh6/MrJRpyEHQQ4p5aC3qMlmjLvXARwwpcnc/iM9Lh+gi6MbJ36uyGjt4eQrNbEjC0q12Ht8
yW7yK3IFhKxyYpGRdzD5NK8ZTH8qxXSzqP8L1/m4gUgFKB2Psp8JswQoqy9fJevTFcZ+TnpJqA2O
Wug/MIcKvA1R/hTUvrzH5REfXGsHzOCr7JBnZ0WQKgsfG0KjEQTbyJ/KZxGAmOIWgOO8wI/Dlj9y
uCy3UnqN64VnoqPmHSg0XezgCd7X6v2TcKSARA6uSPuOnIQT1w+MYxvn22dIBpUe3tfOh5AFCGwd
3K2eh6NmYy58ILq4F+sTg7T3XBo3G3qu+l+Et9R2lN852CCzhvbmrKcHq9EoHaEupC5fD6W0NGXf
DKo6uAIyF54x7wrpF4QAQqeNKhnbRGDORCAopOiQOUf/fdst3dcaVzvkNod2lZkQHUaAwfuKEHcx
aKSZeUus9UeWLSf02w75R4Qa5cjCQ+crLUkp7PNtcu8puOx4CuQVr1EQGR6ex5Q+eTrHTGq/lgOu
uy5NR66GEqKA2gtIv65kZ71q1krhBOf3gs/tJpvmgHXHZg2k5DatXIP2lLOmUwCEErXMdmdYTjRl
/VYV4p4tvVPj4HiJ+NtAPncxN5Nn7706KfcjnQYYFIuT0y7IgGSE3u3uMRYvoh9OrLcsNtGPMzzd
7nIWwBkfz/KmG2CAwQbDApHN3cDeP9dUounBrFNG3mEKEcunCm6n1v45VonqlhOfIdynZW8UV6W9
MuRzAiWxZa0o2+8KmjWnzvQ4H+B+nss9bZ3KZX9iKCi/J6wTOExAQDHSwKpaJnNbDJwCDhbizsca
TzgAQ6HwysSWQDl8ZX1KsNTe3NRG6q/uIKozzIymjpyTdRq22V67Ys5AgQK1LzeBxlu73vz2k7kC
4fnuv55IOQnVHVjOBzYKb8PheA8zojf5eBOH8cumcKqqicEs6LfiXxzItCC6fhBJLIbVbTM3Zp/+
ewi2TlHTxWD/hRWcHc9Mj58X7pEIq3rZ3HC/BBsNz4iTFxDdC92Lbm9USdktdhN9/Zj0PRTwXt4U
2LVKPxz2pxQ1HQ3LOkNqv3SJ5XxMonp2YYLuRJ857Ix7TQL2lhMdb85dcDAZEfA5nSuK1t8KqS2O
LSF2/V6FZA+oCfscbCvc4l2Cr+OIk4AheC6Y4g4J9QxjCV+oX1ro3w7dTOLrmkHnRr/YvY3cSYfa
Y+2PQX+xgvrTPm/OQtaO+Nzm+ugS+dQPCPRrsy1KIrz2ZhJ/36Flj+sXEdmALnD63jScxoDVcNSy
E8oNOydseWIx/wX28vdb5+7NVXXPbVPKNT9Vd/rsqDC5f6h1+XOIuc16G0rXczN6WmyKSgZMhFj/
bPeSb4M5oVc59xd5F7+d2PqZGdpNkyg485gS5XIBmNSl5NTokMdO5ewjAbhPXD+jD90P5u6/MckR
QUXLlhHcJqBHiwMu6a4YFg2zqqiwTuVCOyjdVtoeoPvWrQuM4snQvSXUE8Hv0Er2TSlWVbp/QWjs
4lXeoVuthP5fYgWbYUyRUXsg5jSVkr0iu3RP1Z0Sin65QLacqEXjNWVWE44vsX86InC9IjjyPerX
uUhRvcoBrtg6ANrqzNwhSJ2nZtQD1NpcsO7PO97RgzBqTMAy2OUVrKvPX8HYyfQiwPBqhLX16+9I
pOBhVDvRzTmRO0SetmV/8qWwt6ssFO22NQTD1aHOqLc8cm9aG4cR/zq4Hg5GsuuPbk63oJKxYnMF
pKJErSIHqO5hJ/ZCRPGbzHFzXvWgVAdnLZ3sSd7uE3Lhz81JpqGcbVjv4j2/499rM/CljkBQnHRT
IMqDjMmgYioj/jwmjGnPSdPR11jCtvnY3t2Paf3LVvERKPMJhzTBryYktYCNhxcenCa8qem3IU0j
6dUODngUeGPK2oTBthelRj8OKr6TVEARcUBxCy0xz79/6sH1a0ZmrRETEHsJcB+RyRbXbh45DcAI
pkHrBYP7VAHr/Jzk5CS7HzeapiCIAoKpydfJLfBCdp1OK1wI1v40AHmLxz135hBA5AlW0xmr1OtP
Bjc9b8FJq+mmn+zD01q1MIglAQBeCRF9igux/mNdcoE3FnvwWwJO4XLitBxeoGc1sLMZ/oS4W0TQ
i7Ju2xmUFTY+j8UBbY08oO61ZIfLfZ4n6GywFwA4HM6MUb8xCrr8sFrJvT6OCOJiuxaDmyIS0Hdu
Ne/bAX50t9jF7XZUEp5KY5PyqHx5umHx3Jc3th56CAIhoHleQ8dnIBIHfJIj+jEVIbv04KBJqTeO
G/sImhuWN1WAgOvUj/W5c78DPRh9NwcXp02AjieBOhVgOIIxUT9FVlRs5iByugpPaUpkVHqE+AQj
FJY3yQIYOCUoX83hxSfVEBJgHbAMTU5VuOARN2upa9udG0T/loJORH5ojLtnOnfUeQrSV66mDx6c
1wYOxaljZqZv+mySmY9/2Dp0VqbaC99JxltFg2ox+/ZU5hpvUFo2tJRtW96Fy1LoPVY8hwgwATd8
0pK/HyFDpsyvrcH6sUBH51fwtzf2auHYvbiMrvKV34D4RSNnYo6MBmIa8OZBXVUZE7Cu8xHqdkA+
h4pa8PshV3hEB1+KGYDpJ1uCgZ6jcYeC5d4F9rudeLQmcE7EEZ9cfsfvjA8nbbTH1IR0sVCAHuOY
IwwaFzRrgps6LPVod/lLrZL7nXJV6WtKAKc0NToD2mAnbn3N//UHQnyJhuky3qFvKedt8BqSWqDA
Au/endTjKxJGqazKYF4EnaaSTJN0QQPnfxY/unnfhKOVO2G9VDb4wmUf4mSHFqVanCkIvewzCvVA
anf7WNpV/NOap2KoRAchTsvX3B244+eUiRQGr5qX6KlKITnwcxRIEBdloHkL8TKlmKSfkULFqm1Q
O05IBV4MPPfA+Ptm2sC5LK1/g9wpfEw9iBK0wFIjLZJufUBI537MtQuWXKWCRh6a/d36uVVaul2i
0pC9HLAaTe22rIPKLs57wgdNddeCTc1pdHU5F3gcoPomd2DKP4g9syn3DmTQEOWe3MSTRgOge5RU
8xgwj6tomyTwl8EYeeqqqK41Ptc7JW7qXp1ZOzOLmbKeqcFKG8zIq2a4ZxumY9caQaWagfMRPLCS
RJeFVpKQiYEZF8sLTaYGsUDpnWawWlpQDZ8ugwAGOx/uxNkcMkuyfLpGgrG4OrBG8dn5okh7e9dz
eW5LsPlSG7gajXH42uxoXosveKWxR9di4PEHNvsn5P83MK27yDBuEly9uFQaXtTWKe8G8wN9GXlQ
B2UB6qDbqu0yfdvy8jH7T7lQMoAOHQQu5GBrgz0ZYi5HJWmqpQJqUavO7lV6wRkl3E1Ag1bW4kfz
/z52OZW2UXBg+jYeBfraUMHJatlv0UT/t3E6mB4v+TuqKs/3kP7V6Qy+UikoFUHf1ddgtwoEiU54
NU8n+ZtqT55D4tHS2Q3uzdLTpb63D1z+FFrrwPENUB97QROjyzg85brgMZrttULwLhRZULiSN044
4WlwF8Xoflje5pgGwEmaz/0+gqO0ZRAfJzcy1l5FSmnQqFRaQy8tXD2aOURdA6ZkXxGCPn3hZAuc
WV1o0u3SRBLGulO3IcFuqaA266sgtjnu/rUe33jsXK+D17UjgPHw7xe4NG7whKliOtmwubIAMB61
5Fe23dXSb6zhVs34pQ39n2jz1DiDOFR/h8bcdNuFtgSPgICCZgsS1xZVORnxetpCz9TSSbuZn9vC
m8Z8aM7bWsp41BgilJlKE4zEgV+LOhAQHolZWDpdBA+RhxAi2HrWlTSRJ6K3u5oyJKqxcND9eSOO
dtJuQc6EprYng1LCBjgi9Vzh2S9ZHUSZBLkUQjEXPLbORhDTrNcjAgPNQuyWg33e9V1FRZlBBgXd
IsyvIicGSvgQUI37B60aKJb3Rq/nTUGuYIsPqIHecTvHPEgzpKm8iu5oXp1DKZAWBCzLEyd6oOe+
cEvtXd9hKulSGWW6Ek9Ct2Ue6Rt2Y/U/8W3amBJME400WFzS1Uk/9cat0si9mbFIAs9gqcZjwGok
s5o4DWygFBtLZoktrviZl1UwVqHN5etHElT9jASb2q1s7sfkDGGkIcL+SlCMinrCWB/N2/MG0Wo2
RiEAI21SWkY9S/b6bTaKiIa7kCCO4sEtJmR9irPHoeI003c/88L1evz4lwWWkYqAYncaUX7l/htH
9ooj+4EJoVcx6xcTTT9wpMj8WLbgU+j4RiERgchHKpVOVYXJ3rl5mZZXmmZqqx80Gin5YoObcIDA
KQVOMjbDHAshO/ACJ2LGi6djm8LeQiCWlQPjrbqhWL2kjZJVwcIAVfT0vQI3AMhLM4U/R28zwUnt
vVIltMqxuThX5GoB/gR8T5EiK7A8CdQE9MS/SAsJSl5JPftllS0JaV/+jkTSq17kaiPT0P4sNp3i
/MhW7IqnfutsAATozFsZAFKdWe9sLSyD8oJckUXR1TTgQDWVpLSLO8wZe59ElQtgVo09JINCZXGD
YaeCm6J9wgTk9u37d4ETxZmD3CN5qTfzhkUXI9NN7zQ9zi3/5tPaYhbLpgTbTeEHmkRHA63JzCKa
JqUqBZTzwN8W/imbneu3faIm6V4jZ65fAygmZkeQiiSJfvp4YRCkooIn90xONA7zbG6nLOtZgH5w
C2pxBIKI8IndclsFalQB21g9uynNB08igITKJERXrE68XiRL59C2/dHZFUc0IIg1A4KxPQwmuPsu
GoWEnbrsT2LJDNsi4xC14LtLcEmDTrsM5buCCVBa17L6XTv4XV8iMx92p5t5aeAlRNkw0eOVhPrR
qK9i6Q1o37Zozkaenk+aLjZqrKqnxDm/DaoFk5ehHb/dwxeLmbk9P0Y609jvNII5igEYa9Gx2LNH
gImB25lO9uYnhLkUsDOIEmy//THS8wIiY/YSyHeGraLgSiG+YUgmoaG+xLFSa7ELwHrj7kc9Da73
HnEt7EJ4kasimKxjHd8RQmNeIcPTx0IKn9SVCqqt+DAezchEU8aGvBHPJSn+ht3Bqqdhv3oDn3IN
64hjFP466+TrymFb6zgnsyy/QujQjrJjUGvZDYQaiUZUyTgS55KtIAsEMb44uOEKLoa5uFBnrGLz
RPHHqTQ/A1U5dFpih7sjCmfD793tM+BvflRv+Rq/5W5WnPGHLJpqz9pX4XIFzCCmOmlYwLp3Upee
cORg29BSFE3IvFFjlCcICTsD1XQKpcK1qIjFPPEtli/FwnmvFSgMlsT5BR7vVVKCzkT5S/mLv5yJ
EfmBYHw/s0Ol6jZeyC096iFxnhjLtAzxXTVWaH/SoXWkudbZZqTrK8ULcCX93a7o6MgWStKhElAe
ayuaukwj4wobUE0jigGJX2uFoRNVc89NqPcxxLf15HsBhvdHFwqt+K2lzpe+k2c+0syWiR5yp2IU
KtLx1+y5YWBPojH+onZeTjusAYMgo5YJxhBlToSx/FqMA3WXKw4E6c99RJVdGLZQx0QGopjw1nvn
VYl+UhzURipucVI37u+1gnx1RUfSuEjTzPSXrTNUS2AJK0rcvB7nB8ttvBIMEK3pb4+9NhaHkv+P
GYwFSsjrdY4v6d4wFqpc6PyM0RaTlsEsl9TIDiLL3yty8Lu2x03YB/63dyObl41xA6UdoP6nRVVF
t2oliwqj7zPoNZSCmwaHUsPQtGq9tvhqb1Nr9jQoEC274zrqlJQU47+IfhWxfyJfM4OTj/qSwP7c
LHKfD3Ka86ZvFA0JXhQ40HZsKDKEDwzxWZknxwZZCcm0aSxR+uSIxJ3GJFJ6fB1SWG0WnXgapFTE
61dMQIdfKUs4VB52O4ukVIz2GlgiCcvjggafFF9ywc4L8xFqR7BQZr7CNbInfmSVDuLwpC+XDgiI
t2jztH+AMUQsYWRCV/ERw5vBuFfh806X2YY4Z2Vea5sZxeH1OqrUTM84gsDdanssVfQ4szK2gVae
xBmdC011KUVKa4mUxUXh0x5t3rWYKTRJqpN8YSI5xj3H/LRcLMCspal5YO/26nOK79fRiRzZDaFl
BuXlx9uYJVh9bxKJkIxAm+FwyjWZF+YIjzn3lPkyYDxCJ6QI94WDOsZ8u+EIpgt2eDDtkWtsZu3T
5865uXwwm9mRkcXaR0SofRIDOBSVORJKDY/U93uIrznmdZWHdlN5j4fHqEDLBhqJKoaFSUXbi0R2
ad/KHUWc5dkTl8a2ffJU0VP24vP1tGCuaZ2L9wq4GWdbSdtLR8SpBxTPBMo4BwV5xZT52nj4Ex+1
VH1/AJ3leEAwXDU0KANuvOjBOqQLviKhhuJ8K65qe6H6awcJBkLNCf7NeqfpAt6wK3JwC6Wc6D+Q
TDd9YkDwud3N2/Lzyf9JIpi3nOtQd6IyQRW3o2lDjhI2lSGmjQ7URW/NvdQihU0T9aanLbb01PbX
ZTLvgTAZKJ9dr+QsPpqXbUy1Sefp8hFPnHTiywXRISn0+gi0YDZBmIF0h4Wl4pEudlcPZiO7eyKO
d6sxGc0a6jV7DISz8oSNUrt6s7ZYo6/uqR0dX7JI6fyalYvuiVUbWhx/W8KgnARbTtdfVqeYSJCZ
p0mu9ALioBCvsQ+RYz4guey5X9rZukpfhTdh2bzTyt8j3cdYHoURKxbshf0i7SomZieppIZbMLKY
NZYKUdtGONG9MuWz5jVtXcK+3cFWonE0PdByQgBDJrcBLMRcXI2tTNyfpIXL4sME7Ir2OXjzOu6l
I0hMNC8luQxOFUxIcuziPJ9TMnQm1S9GN0VrLoz15nhMlFbL8lAazA7MC5RIkIi4pNLRe0R8qvB7
fPPTwcMi/4dfZpV3TuSfPFlJhPQPOELgrRo6rbF4lRl6DlirvlLoV6PPlJdQjp+XaZFChDJY6j38
zyc6sbfAGKnWM+C2N1aM60fgqA0IC179LV6NXF3NjOFlWTyTNRKhDaLWdRxF68GUJybEOk0g1/vU
MpvtpD/vKumGL+5nWxX7ufCf+kenCUGvD2DXv7ccGDiniBDJNXGn4HnGGV3BNh07bwW6GIknB2E5
Y3dGe19ZaQqY2y+NRvDsGkM8n3ayIMosqzevshhkOzWC3+1XWmqRL+OhRtrt0bIGctDSWB+sJdhR
SXmy7VWFuPvG6KMO6TMWijBUElrPMcpKXulvNOkFC/2Xqmq3hSOvKnQF75st2DgnGzlQbJADxkk2
NSJulQm3d7LFdROkh00wt/BK9YtlTQr+cbdOd3SHszIh6TW8rDr4lMG3RviXCY2fMLZuybWPJEMV
jhqhJ/2u9sqjnd6Tx1R5peE+WdaZxfmOcR+XXVCTX4PjQynpeaScfb1zAbb3X6Wc1y86pPBgGMqg
iYr7ozkhii3sVFMZqjujT82i0lcKgDalJiLFiTxR8UWjvS4fFrLDAUTr5dvhYJvHzHhUmeZJL7q9
eWkZilmaFPWUV7NiDTXNG/HpjEi62OWhOsflinJeo9JXfKfeQ2rIfp58stpvgrNB95o2zT3/d6Vi
gt7Ef4Gm7gbdfB65NvrS/CoToPfVHziwoMoT1vHoy7RWjJXZDhbKjFNA8AwCHk5isR/8fSM39JTt
xIsqeq2vMubxa68B80RegMZjmuGrYhFvi7TViNAk95HVczHIYnjLeIz7yigYE6h5RVHPTPet34lI
PgZBItQf2vSakooQCK7MvScn8NpawKrtpwV06/4FORAhz0xTDrP/DU6zaHzrlDKBO7lhYNOHpwyn
f5X09d3tzOWniTOYP1SxrsP2YgQJX1B+d4fXMdGCSRUpBUYKD66TyH/zgGIlv09jk3Psvvsr9nNM
g4dETZaimV9d0YcqQrXIL2v1C0Hseho+W3B8gXNPQWLfE9wxGRcATmbV+Siq1ceZ8CuvrGqdq76y
48wH2JkwesKiXClYoSxewB54b+onL/ISFrQoMG+pkKBUn8K7nWHGSEV5Bao6KgqcYfX0wyMqTksO
xQ8NUphlThisWwWr9SUqEo+icEGLMaH8NIaPrPn6OJQBRzajkd8SdjnF7ffnadLy6QmxJe2D0bpN
Iw0C8Js/l4Jpts4/YgpMEeRlZtobFY491LkKtGCqRDs47Kj03KnG6V/vqCpYbDu3T/aRL/ewbr3S
/iAwB+r7lgqJ28BvB4P5lkyndtZ/J//olRqB6DltLmav1KCoXBPr8m6Lx5Yz5YwwxYtQOsKDTOJz
K7XvQG/78cRMdcloYaH5GN/Ut6Fkfg5yHugGk96VU+EKurKXJpg62X7vuFQ8a01C2jGyO73u0IxF
0P40IMusqOGxJQaeJSwpehy0pZJ3lYk0r9uNJF4yS+S5wNRsR0OWe2aTZLEX9tw737Tc/pSaMAr5
dq5IP7Gfsg6CjRRLghB7RnCaed3UxS+IyopltNejoqqcCiAESr8A5Muj0uow9zbN3/57VtMpoQxq
mL6JEpMuyX1qosRKaLleH3FbiticT6tdkymly49L4wlFoFtHWHNYpjpSjKR5JGkn3IEhKivyJDTb
zZY7o7Zykrm1HiIjmZnO05LyIE8fMSoUgdCzjKgh793z9CfdqBEU+aoPBSxJit1lKjc0ZSVkEWE5
RzcIdv7W+IVnufMUkoFidDgM1WwsAo1kl+FcNsWkmNMZXZropD5yNJvBqaqn9t75oYPKT0oLH4YQ
EuQhti9TXYOKQop5Y8CPXApTt+NijESSLy8h4tnUONSBocpaGUDSTYFDGxFl+irieS4B916VOCkM
d1IRHApF5Pi4zkSLtwV/Ww5dFLm9WBFA3Ww6eoP1VAKPY1c7PmGdV7NIhpo8Pa5WnkqAF9Yoi0XE
8K0/ihUWK88pvXpc+/aAkYR9HvgoIpCqjhiKX5YV2ue6nIemlpOoeXg0cioIGfelXMtXlpd+KJE7
8NJP37Op15dnZQe0Pyzw5TOfQKNeCBhuZA9Fsn/dK3S29HLQwhLE2vOKLm+9lD6Mp9ibJg/SrPZs
woJIa5UinYfWyeCAF9LoPCOvGaQ/26JQfuhuBHmw+W3v64AtZ2BaEdtYLXXQWuy6DYAPYKfdP+MY
bAb2eZFCmOA4I070sLcvucY0IvlUG+ZG1PTkG8M81lp1D9uleeYqH+Amlp8NdNPJaNAuHnqogTa6
zLYn7Xz+dNM0N1eUbBnIBQXl6NfZABN5AZ8/HLFJrBu0UpeE7HWNgZtCPcM7DBBUEBIb9i3iCYMU
VER+QQZor5gB8f8TpTql3ezOMcT9rinHhXFjNsohCn7Xd9Z7nApbk/lK9y/IubhH0dtVkP2H0Hs4
5XcsqXhuCswES3YTMgyzUwtDbkcj6U/L8PAN7+aOdEzy/ZFduPh2hLhVZcCNPXwjUfIIwoDX4Ona
vbygrrGAby+0jYEpgQgwr6vaynhWpWWIAw7pS0ydYKIhDzGjfxERIrdUreVGxOH7bx5XVOIi53II
nwwVGvVyWdhk9eiN6zkxXz9ZlMKd9myQ4CQWv0V+uhMcQEgbKG3OlNFWtv0a6zA6qx2/TQgdLbn8
9IKUlAw5D48a79K4YyNOzBmG/f5UIkM0hel5jTfZqs78QpSfpjdulkRSVuh8R55kbTFAsrxVgRU/
6gZPg11pB82L5Cit01kWHtnSKyV/xvHcjlw+bPm8lnnRBr+kjUO5jYjN6Niq2KbLjZZtQWDabA/T
6CyuQf1YJj4Ytgp2iG3PrrKB2CLbEyEia8PCwz0CvnMnT768ZMDtOfyEWgzS82NWHT4AHvMaCSa9
HfvV5z/r83QO4qioNw96un3y3vXa5t2BssOVMFfYYPsB7dMH0TneNRYj9MhYzgDN6dZ3fJmX+Ed0
szn7IJgVZQ0i+T1xxF8k9iyl2msn2xA9AuSWMiwZVLC1lOJSDBR4juy7YGk3ULPUZxQgfpCEOQWm
gWgOkHvzzs45mT7fqkmzYc0vwtxz5vskFZtvv9OxdCimxQ0Zbejxw2vbjknk7NUc1S6ilqWlo2Ji
bfethsOs0TAI1lvlxIR9+J152+qlGTU9Wymn8QYpgNGQERRBShFDZDjKxHuflpTbo5Qabl7iZ1gq
hT5M+whGh2zxc4uTlhLUWnDSwZJOySO3+Vjnr6RS/w+0U1fVnFQto+kX7GuKADKu3zpbNK5Jb47o
Y9TpipnGWl1l1kVk3W+s2PUnUEGdYSNUQDxqjTUu6Oi6AqHlIDCmGtR1MEiGHtCaf/+QPsU+9/od
OwwQyWoHSW6Nw5IpJMTmlg2mpFpM8GTg7nnwnc53l9K9N59fF+70yVxm1fIPI69zez9qIIqpmv49
3q1VoUnM/zUqtr9NGve5ugEnqxHUraPfX3moEHlay1nDiKRES7QB1E+LBYABNpllpnSzs1Hjsozh
i5QuX4zWjNpa4vdDyPFEE20WosYc1vNkYiVepVUwvQ2PefxhawxFcfcp+XtByj6HruUQMDJki5BH
qtaeSYdwL+rex9/xCI/HgDILQCBPVhLs3icrdCAwJG3Qa68gHfSk3V66fhb61wICp8GYqHX9zRy2
J6poK0YhRRhgXOz+IWIlQMAHPIPDYZHVHNm5FKC4ofYHkCVJEnnAyqPFUIVgt3dlx780elbBSwBM
/xVoRfKIxdQSqLIgL0nc+niJdFZTC0EH8YuFtwhY8B0LmWiTRWDJU1dg0jS4sV9O1gx7vPSaTJKt
2BggbUxwDrTV1nU2rpA11epMMBNONuNzy+h1M2uIuiV5alt9z4dkw2IljHkuAfwXXpvDF5wR68ZI
sBA7N1hWsaAsk4OvytjqQ+VOvZxkWUFzEvFOpvKs0VWF7RQ2Uhz11IxRTN+btFtqykKg7EjfoIIA
u8sQJBoVA2Dneu/0qf7WWSHYYUXEJT+Z5AHiXcmxucwlPT5awwHmPK4fohNy+yHiXQk0b4DtnT/d
orGxyAJr1pGnPYVlfyXV4HnZ3Mfth9TOdPZlDd5qUyXCroK1vbPaR/am7hA8muMGzu/1ZBEsmtEb
QZrNDbnVmt+uBbDOYoQJe9gzvrYmsHx7QMmpHpgrM1dKZPBkSGcr5XkaqlgXnCmhMWuOIFJ+tP0N
gljN+ALBrH5dqdSsONCB3GsOITm9DIp0o8D3Z1UE+U/aNDFZR8lUh8iRNwTTRtGA1TcqTZ3iKo5Q
/5S1//fkMdnF1qPZ7fQ3ZzP8IIKn3Tbg2wLALxWzTVkRyz9K+JyKZHKQ8BbdY2jtGqbA1VJqj4Ap
YQYrRJ3BS7j9XXIMOrfaLREXJs1O6giUyK6NkZw9VAGgPZZ2GrM9fmW/VnOYqjoBd5xFkX3LnhMP
KL+eqdNHV2B7cpor/WcAF3oFLQRfrSffEc8gw1SHbaVENb1vQMxB7xxtBE6U+euI1u3eOgaDJ2LH
tbcVSTPTv+i+W3yYhK0oxFdsMQ+44bbDol3N9mAEMV2hriLdAR32Gq65R5yv3kH/YhiIEv0AaKaw
KPPJZ3LHPg11I3IL4foTDZjTyHHHivadY987cbbRKkah5GTh+PfKEGI9lFHL4djVeBjMxE+Jj1xu
CM0z8ZO1//xIAZhFyazm48uwf8Ws2H03sLtnhN2mbDcbpTzhroIRrMVnbqIEyHYdkdVZH84M9pUm
n47745GGOI1STVpvWUReZqO3DKsAYNyK6pzMYPSzF8RCeWkw4b7oiluCDyI4HWr8djtblWOmHGKB
YhzyndBBrFqurV6AU4z4N5g6LFQHhyzBYjgRnWMrLS3iaaa3y9gLv6UZOgLaRkk+GM/2jFPDDdgj
FO7n0pql5Aa/KSsTAxul41I2wJzB70zWukfRsV+s1vy1Q2N5gDzEclSJuenAw7C9eLxsgfNMMd5E
GJfGWwLmIK9J2HrqyC/f7ohFiijo/e3Zp+qo2y9NUR+WxlOgaf8D0lj7OH6otmRn5/3gCxGUT053
c03a9vymW+rDbDdcmw06qH3G8tgiaDzO8PsXUpSFdjooZphWTNKWC/4FcMbrIxxpvNARwWmvQ29C
vEyIRKycS4YtqYwl6iITyWXHOaZ6CFEmiVuj7pUIVX2ZUbBJ+nYa9LtJd8o8k2s+AGpPxqK7GgN3
7X9BF9A7+m+yfHSaPDAdhW1Fm3yX/hryQBm6UQybTSQ1C18EbaRJbuztcIgkb0h7k8iHwAGLJopb
tSk/vJ4h1y8TcqFeK1PD+MhW/SANny0EUBZKBbF7VZrkSi603LOS+WMufITbUVzxiWvQvbSX4m+m
QgnLMbXTzBI0AU72C8aJWZOQN/SigPYpb6s55CpJ+0kFc5jvxvPyEaHMBxFIscaPXrVRqqSt6Mjq
qE8cmcAIlS3BVF3Uo42TOoFj+6sHha+UlwUkAPuq6FBpChpqKWGImQDOWppdX99vYu8mDUG3NJ1Z
UjxX8e8GYQk2K7UpSheYzGBzSFCI4F9Id7qZdbfcvGKdImafIn8VRO0WDnolkbG3Y+zWA3Y1vdMD
kxDd0oarwKx5MVnx3n11cEQU32xfvMXXo897vTLyZVImaX8tWjM1h8u7WKvr9qsGXi81tfDuw+dh
zUZHSLWGo1WrpnhjSIzEgTW7+emSpexbDurzbypOs83sfxtleSL0cH5+LFNSAX9pKhBPHcqZAIeW
nK37oGJLH+KHdi/tkooefhd5Yq/9OGZ0TbWNGUmYpIUrqHoTfOa9mS32OXgfnwGvXrhpOXXU40nC
CnDBAvXT//drhPExmilCFzWaWlvtVehDXtpewTbb7/kCRI9RIma/S+aTk5lhqMzR1tRY3kY6tl6Q
+pDugWvPwQDJaHX4VzBsBLaQVw0cP8X4AeXQ4/ISLT1ixLhY2Ts2IzoTvKHaVTGgf1Pt2MCGd4en
Sc7d27wcvwi8mDEOMfUq3qFvwvaKGs2m7h5WYBbqhRNRtdSY8ok59llyXG/icwvkwLS9j5VsziP1
NkoopTbfHQi+eIGMTJIRqiZRC2cNBLxoB3T7QeR+DLsFm+S5pQis1zYurFaOWP8Q01KhSALTIGCm
zpyda+R2k+/MGR/dHwM5gQ1Wh5ZMr2bMQxn9M18zJ9hQzalmpGYbmrGCoLQV2vDr9x7hkoMOs/9x
RORe/jcSgXGvUInySUCskcZuTvgYqLYk1eBVrZ7BemInrOVj5fD5cwtqm/EZXHpkGBquiS8gmfiN
rZZjGWzKABHzdH9TOAh2xkbvRzC+DPuiQepH/AEjxs9Ap/3KfAtFmmQxNLzspcGQ81VgFh9oNZjn
piRcwe990rhK7b9AgJt7nve5/33F+ECPhdtcwARBspriOwhuk5HKf414AtooJaSS/gmlJW9Lbyty
o230gMNJAed6A6dcbNZuT1jgl74TPl4sJ0BukYhI6tGtN6Kqm+wID8MxEysa8lBRzd684S/kxYda
MBENH3OZ5R6og74Q3PHbCSStHGBKBAvkpgSXWQHXTg7XMzq8qbofV+sjfNdS2WP3I9jFSlyXROlZ
MbGMwvZwhUqp1AFLj+mU0iVlzFTbnXXUvNtLp5xEArkccevxTWoREg7l3a2HbtKK6eZVhZ+FCmHM
v1mKRcDXnWX8n4eVp2nYYWPJCMWt5vPO/VlWPsnYEzQCLEuIpJntc3Ml8jRUyw6+z5TIR/DqYEfb
Ktq6bu7eX5i+HDKEIjwp9YmfeSAQmSTe8t22i7PGAyW+QxnKKDp2OedQNqS07yGB8C1iy7GkTowR
VVwtePY2YUXYbM1JAXadpu5DU/EZ9caXqsE6seYw0TZ/ZfQhhl9l3fD7X30d6J9SBM1b9yE+Xd3o
baoca2ZJiE2lxthPduDLk1Z7bFVxKBxKGgus+7/wOP3cWGsM5o3Ma0dl6Yy6hH1RURH2jCvryL7o
H0EGINX/urKthw0cTw23ZqZTVAo2Gj74ePAGa3UP/iPSgE+W08m3ii9EkxAMSUCin5y+Mvvp1Vcr
ucg/hRfdg8AawXP8nsT0lF+eGbXiLhUSfqEi5Dw1tjMuyU+F4bdOF3G3fyi4u7zLkRzPqAFN7ymn
58hY/wWOnm26BZdVDZKa41p/cGZa1MZZAPK1oIuO0s9O8ot1LNqjtm7Tj9Uu2AjZqhpUZJ1DwqZC
H5VEAIm9pKjGKj+VH0738TXIIlBIxD27aOXg3H+ILnQkvlNM1BkjfBfCNdG6vQY9An7f2Rp1Ac8b
j695r0Md6li96v3UmqYVlCyrzubuTgRU5P3KR3AFVyb/+xcnNqG5P7ZX7K0zNKWj1So24l2Od5qh
bR5fjKV60jPONUtppNDZoB1IJ9YuH5mVB8wRv04FC5tAPZtMxIqri/30WkwwJrBIsvhx0DA+Zsfj
OaV3JXmSB2pyx6bU6EcwKEtRFyMFTH9TGPIo6IPhKpo6vkkJDVKJdJrdwvwClli8zHxG7aRlztAW
A2mk3lUU5zQKwZaKhgE9yLQXoPJdZXcCaUDRHMgpz9/kWSSrJTIB2PDfKRrwSXO976bpVActJ4g8
hahmFHw8ZwGtfotPWshwiLODaUH0kiETfdgHq0qynA1WJiTWz3ZtnW7KsMngdcMQDf7H7nYYJuNG
ccw60sgHU/hwBxgdOwH2scEEb3/cAPbqQboVDcQv3FBFcnRvZFwCRBWrMRPFAYj8dGeEsOmEGxzT
nz7jV/MvCAHjJm0HuwxXHD0IcV46EKtK4FQZn3wY4z7/UyH3IB9DxtP7xSnYrXT/dsi3qE1ZHCu3
IgNUGeFgA1Gomp0HixOkT4HzM++wLc7N2uoZuU725vF8sglJWy04fvcyEq6UR9Cn+s6mS/4agJXx
Yy5x3y9LCskE3CKTNTpMmnWo5u+421I7IKlpfSw216LGNOC9ByEvIj0T9BdrS+e43C2CSIGAySFh
CQm1PZnCT6S2uvUaSRA8La5XBqBJHFq80SjNp9KGSZkBT1jeXSOAn6F1TF+rCdXLymB7ET/8BwRM
TmDgChlEf1UF4t7hI4VUTx2gma+/ptZlkKmfstXYxybPoJG6hmck7NWV2JzJz1IjUBM8plwa5Vt7
UXnHMNRloBY/RIgpeta//4IT2PTj4pr41X7f3VE1qNoA/4iRvtRHh05j27j/n0LqjdA1GctUps74
7AchoqMpk85GkgEPRLXn2d4Zzi6w/mhwslGG5uC654BwHDo1PoYGxowfKLQdl93R9+X4ics1snNn
tgy3PJvJy3OA1/mgpF6lG2raRMEq+v071Y5XCARoBx2ixvP+/tpGv2HDA9l+eC6UlObsELeLBauY
qs9b9Ct3j52ctNsGLpgnTuXxbIhNELDLlAQ2u8+Onsm4fHCkE21S5hNCeXeocDLkQaEUlgurbwoB
BhSdbn22ryz745MDCltUm3Kbiu0cVH44oH6Y9liaFmoLSNqxld9YiQumiOnDZQo5pU5/rnpg7Tnj
Q0fWLRNXJnqphaWnnUsgLqPVb6dzw1OLZCXOeVFW6BNELw45GemLrW2lX5PVjleysG3IqrnfbbeB
uKBUylxQUA3uLeOFcNsNN65VfBgxEfefOmczuJXx3i5MKfb57eOLp8OcG3gXfUiTcMT8dUceSZHs
j5P2rT+S7eF+wlfFLdujzL+GgUe9bF0aM6myaKwqYGqeR054KcvNzVTjJMBsklTTpCZGUiPVGnIg
tnKehr4fs9CFXSCzAPG35UF5PQk6scbIwg/y8dfLg5Pquf3cs3wbkI+lk0jJG5Htt2djXuR29DuR
mY7RSsRqOYW3hrDh4rZW5j6iAytJors0X8vgUqkJaBb1rfpBNPU7YmxF3TZckCs4mjomnZReA3Ca
AiBPCD1idP+n8xemV1XRM0lKd3jz+RM6g/h/ytTpjRmJ12TM/j9jsv3yBNsyEXCAyFZK1DqaVw0M
K0vOvhjP450py8K21TICoVOpgFouUOYKbeSjXyikg4o50XN8UHCofGR51p2He5/FoI6SvOy/xHEh
Cq8JcRmgfoBjhktEtKhJiRuCcgPxwy8hV9kXYzn7r/xrNFADCuqvjAC25FJKnOhFIzW3HARcJb0r
/5pkzxP6lnj1qTg6IhNAIHQsnZ+mx/H0TmUUW13RP5Rz3xxQwmwXR/hWKOjWNptlTwOJL+/g+4H8
O7SG131e73GDhg76heCGnbo1W43vXyfwyDEf6a0zB80zwESATkXBY00IeQC19QF4Jjj4feLJvpE1
RJ9jPX4NWnvmSRdqduescw7kJjCc+elPiNtbgymVk06e15sKL3N+fuGYGrp/g/sAunrnGFb+Y39T
5TQqdiBb73ceulhu3heedS+KYdbJHUsm//rPFCPOJJiT/4oMBO/jGZCQ4x1mnKKhRpDB8yKrNYwa
2NuWGKUdWubBQ5YsarYyrjqbjKuVOwAY2h3W4ox5S4hfXyGpSQaGcEQCvxD6HmlYS8uvEJGZaU0X
PQD2lLfDY3P9NudiToCa8qQFAAXxoSsE3nOHPARO7intQ+JeSNXs/8e2egMSak1aHxX22SjmAkrt
Txe7nPw+/J5HWVmrYTCtuZIeTUJlBCy+guoE1ta2b2BhxyTXBDVAz6oHcOE7Twb4GoP0LZeeFUZI
LIIygLMfKYOKLh/z81o0igarjEtzqMNVRDYaFMwiHIOooiZhUPXuuAzT6EJjW8RYCCsZrRfd0b1r
27lS7DXPs0Ur0ZhPLKGti3zuZ2+xgDyUe82gYZVJ7g4xVc8+4SwCL4gCT52a6wlbnIUdEecu6VPT
8ShSxV2YeqQKpYe/kwLfVPbN4xnYCOc87PstPFT9g10MtH3jxj7zzEd2iosxQg856iSJToTsjUwI
O8zssKT9KDq/JUNGYFpP7mGVlUkr0Oenx8YLK/Nff/wGyau23NBN9R0ujahJ6cjZjcTOEYPgguYJ
1aoEJiBnZboxGvocJcscbVnNYceSl2GfOzrD5HDCcOB/cXDVuPzP9WoYSHjbdmd7c24F04LiBCgi
YDtViIT1jlw/Q5t9ji7OPdqxQlL0e4L9s1owqoebzChdzxngh3e7pC+GCuY/luBjGjZRsqgywEw0
QgtwppqQ3ET7UocxlVDkuoSZwpTi6G/OvwuHgYYowA7PkpAdisHXifEKC8GtLmWyQhEP6NZ+gfo6
sz3twhNs7SicSlncVuPSRdSJW/JSMR0IsyvmEy6Dd8gCxdQOZgAidpiv8hsUeVgf8L4sGhzYG34z
pl8VQEgAAKcOsort3lGAeeLs/VFqVCpU2y89kbL1G9IDqwBfctfM85VO5xG7IBRjM5Zo/KSfXn+K
SU2UBeCdlArWDCd1JgoLN6LRg0Zb8mFlwclJ8L2r2oIRF/qfYhGIvBJZ/kDfZoOwvivMnqzBXhch
bVSfm0Q+ZnIAew91hWWS010CmR/p77mDtj8rzg1ZrtTCCykiaoExUQGlPd3TzAAnVPn+Mtr7scu7
H6U32sLyx+GiBTp8K4hbSJxqoiPsi5i5lIvNDZ3E/mvJUjQMm/tqKJBeaircOEO9GLCa9htjgOg7
ipWLaqhczBFcTHAhqyUjzJB9uzXSu0Se+Kj1cFkO7CtVZSwfCRjdO74R9yr9Pv7POECSDyRTXfVa
tPF7C2SYFs1kDFbrLshEWXHcQ+px9KPfQgTg2OSaJrsuF+BX9zmzGB2mwkeHmNrTKTFeW/KT0fTH
rTR/zFxoH9sR4NswdIYvexrzL2bwVI9VMM24WnR3kqsEaQw8q5ZQDZQ1rbPrretnuGjY1iz8/G04
n7im6wDshljeA9ZRRRRMxMb0uBasHukfAyPJM5Kiz8zW18/GnsTnUES6p4433jaVqGFIoQVESGRO
S5PKjR/8kMytGWR9DTw321iJ4oQ5+Wg2YYxtUGfnTxIYptLWAkt510LhNrOOO+2JPjllhUomxzvg
gk5l4WydG9flMz3x2flkVBGGiHV/wbjvci/uQcIqiRFLDeQ4Z18Lynu/ZmYBrCVIOAcxvpVWbxOG
rVhZw2DR50vgVI8maOpdDyGRxEAc8D3mpH2UvUO8OMZ22IO5eZA/dKSXhHitVS9GcUSQO934l7MG
Q+rPNS8axfqKf5zsG8kzE062LlW/qn+wlG9NemPY2JD0KMT/twtQ+61bCxz6Z0a4yMKyp+vxSdCm
qEzrxDwAy7+TmMIfLpvdmA7hnZsPkLvQcs4MNOhupU6WWoZ5mD2bwD+wqdRl5UB405biyAFiSLrk
vmmnCbRw3BfacJkL4UzGEU/REHCCJ9PyC6YpbOcFxCodmL2xJjqJ9LQm2begdOZVndApNEq/KgjI
SYX57AWlmYiUQrUshUkzPc2WF1EDpMNtd2iCw5H5DSTBHW3FyM2M4+roJFPmg/YY+w4OhtDw9gXb
dORsF5BaGBLBw5M4l/NX5aTKLiTq2GTP36z6B80ggz6xy/AfFKAgbuiH4fLUsSXocpBfofk/f59M
hCcWIh/afqBEQ1DAXXZ4NB/kPSpQBhCg91pWSv2laQUuus6bE0XK1aU48djSiaIGDZHKjVjF20s2
rHD8juhEIlvlPX9KcEJ0qvo5+9iSZY1re0Qm8dwgiCJECMC5G07iyXtMujzpYLsg7rYeCWgyaKpF
VVmA++OWtKwDJu+7fmeakezVirvjKE7hGRsQJ8TKsLNchoQ7TE5Btjj7qTzpEzOGownAjOeFchzb
4wHCZIB9FnLNJH+NKHW24EjgPu3o+bSKFyvkkUUS5zxXkA8RVMHKZCmwC3eeOUc9h2ATiTnkkcct
WFjg1hcNFOQoWJkXBdEqV/1Er0//qtxCUDABc57TC+25qrf3WO9wBkphWmI++n1oNCnEihUQkchU
I/Oho2q8snrvcTkrhEyoCaq5zWHQdKG6Pb57Ejd7I7cQImbu31X7GLTraSn8wsYfC7H7Y/tFMpNb
17A7gN0It6S5X2F9FxOcpyw4xqe6n+vTQHsz/vxFULj/s8Ie1Kc8iqL6K3FPUDW6VNUWXngwPyBT
eYc4eHLDtk/mUdyzibJqYRyYnvFTHrxoh7VvhhdN1Vo7SoaLhlSkrj/IbiBAfAPdy36xC/lvQZoO
n9W+bBW5KzrKAaKfCNJDni74M2wOJxrRp35O39ze9GKJ3bw5oQkCjGwtjiWH9UfgpHwM/jzzfhQg
DVroBo/9+uom8vRKri7ZPAm2bq24BM52hkf5BmRUGjhkYRNPa8uWm6A3bVhzuQwcaofpuyJNMZ6F
P6ebxr2lpieEudopGhDqUq+fgYyp4PPHq0RA+tmG5Du9Mu7YRtw3IjbNaXbyfFGNGNQDP0rDqOFg
Ri/p6lx/rfH57foKqaNRuAkVY1fhQuCuZkFCzGxYDf69WSrwSCwzhUdvrljoCaEnXxhMMCo4yWXI
WFBmXQum4rBkCQvs6fTi3MZ31+pORBIUMkBlbbeHzBFnaxopBt034lEPn6BYPLKbsY0qqGqKSi8F
9b3o5G7J4KGoWWLQdQI4KsZfKBABNygGBpwfWvlqBC+KWas56hSXb8fo3XkIubmu7j0ck5aGDtZk
Ol7PWL3PLwSQbKSgR4HYQDgAEz0OpDI5t9Sv2eNYkrCiDMWNA8BfQh9KsFQUiT1q1fNseaI5v4dF
gY05ZLCWI3NQEKcU4bdO7696AUOSVIcCJdN8xcNscPL84w+Doc5cJizcyrfYp37BxrUn794wI5ZZ
z/0S92vv/acJcY2FVjc9PBwfDM10cMSRPWtdLJLegnqHN5s95fbq+zoiUvdjNQco/hSSXsDTqhnu
ngdwpZdWttbh9S9FNE+2D7/hIxbhPphGV18ZYtZ8kzdjbxET/bbS9vUGqfA5agnSB1RPtQc4EuRF
2u92bcKPhsOoHRA1T9HWh68jcbZfh9LKRozPhMSoBNyQkavTDtKrLRz04D/QH9BCvsZHyUFaxtGG
6SsF2/NzY2/KzRsA666LrFauWPj3hb5jtnRS9qf8ldMMIrixZQdRfTO4k95RAyN3qOS6n8NPWLBf
+0kFgFBqA+TpdF7QIGXYp0QmLbG707FRMghdSSi1pArIiJmSmmKXGGgH3KzcjYVRYimVqgkYYAk0
rIe1YSJDMHCwsdHRNjSwU+Dr5ZZHJ+8Bi7qUvH1CjTyNP8gEugKzgUUUun64XPupZXbpcfCzpr0O
51AKcs69uwBGmEAJIeK6ghtqYb53kb7WkJqgO1TbmzdXcVFlV1RtLSiymoWZh/i++0u5Fo7OHt/u
dRmxNVSjfKVNEfUJJpBQXmR4lEostNBxpX0jIkZJ3DVc2QZIdmRDRIs/4bGS/3uQUPHQjmxsvade
bk7ntdv5HvG01k7BqRnEsrTUay+sRdzTjALavfBDwNS7urxLlIshHO9vdep7ERKIZLuIhCrNnkUm
gH+aE1/vPCBXc9Nezj7r/+zRgtmEhPb/z2808+feCPFOy0w9/i0sd3sup7VAh5MIKhl0h+MPhByk
W09EQlAgCOSp7hnHgaRncYnPWLrzPocxUztDQLcLKjafgLj/85OSu4pbBgzFnZUWkUDLO1W5+LxJ
1m22UCNoj/bFOMXCoN0rSzvmVXz3y7PSvKTE3CWNFKmEfSiMJWEMtaqpibMowUuIVKr8FkaYbVAL
JrkXnOqejFv8ifaL7sDcrqdZGdW8vckvi+Se34kx7DKbXlaPLE34Nm8aym6xgDYdyoNWy1uGQafr
5nufJ1q7a0UCocCR82dOW77ZS2nfeZVCPPNpvCpAaqq359bUFwErKmGpx05CGn1Er1rEEcvhtI0b
4FN5mISeJ3dx20PRrkflQbj+dl1kbQIgsQishMZa55X3TjclrJg70K2IhWxiA3M1FjhBps6x93Xm
4CJd5g6Nfc0bDqSWEsMhbYP4Zj6OzImXaD4IGtCFpzRE4PZwNWRg2TYE072Rn4z28v/f8z7Q2s/R
o5tbuSILgAWzidNJG+wQRvOQPbYnzaC/AQgAJ9GaXY/3258pzpwaqOCRSDSODipF/lum7xzNt8iS
yQz4Mgx0OINhqTtLO7rqOzwkA0BbcL2FI0ZfLhSxyp8GU/7TGkxKumrlA4fjCJ01MXSCWY7tDTW9
LtIccyhU+Kw9waTMLKyhMGxaPjIMF/zBz5T/XyUo7oo7v8qFyhG8ehuisuzNwLFnNBTmaoMyR8zq
bPagy6U8OEpdm1rBgqhomPeaU2RLkFLunLkW2GcNsU+Lkop2MKnvdFMik80JX2/b+ehiA8ELgS9n
wJOjunXR6dypqRH7Z2w/ZM7Q4PMzUCdNov1AyDuJRMZf/HuV4u3Ua1+3ak9MtLTDZ2L8qnSLH1/O
p1V4NILm+EOiAshhCEv7a+LiWmcUA7uboyRRV9TP3pi9Q4WQqz2b0Yz1K+oTIulcIg0hovP8/Zxc
5vmpfK9WjKMWqXv+jlqUg1r2FRKBlP93guF5Qiv9FpZ9WzCryKCLoDQmaCIfGEpAqAPOLiWD2sO7
jUdmZvR9bp9MUkZqpWyP5GDHbxyCb8i7lCoJcfKvwCQMZ1JajFfwkh22pa5Udoxbcnzl6Rr0IjO9
d07VayYPjPn6pg3vdpXX9BtNrO2aqZfyT+StDvDktxx6eqknBS6+IqefMyNQ/ui8RlepETEiSnzB
tZZqIYWlhoUwyWKZfNBIZ/vdLpJNq7zLC9dFRJyRGhTCnANFHsc+ZDiU9TjX2HnBp8peljwNLP8/
cI4EBwKUV+MGtmkTzIau3OQec5bLTeYAsEb1fSGHmzl8TgBe07/VD7TBoH2I0d+Ehj35aIX/yyeX
+S5Xa5a1AfY+o43YqoWWCoC5ikv5P+ofooaLumDBwVFZvdeYM9d/qOksO+QiffpItVO1bSQeDyus
dGwmRm+MRuzjgLtPephRpDUyZDImwzpQuW0H45NNnlhQFyb7buyqR37zpPKr+2PNWShzPF5pWG+g
40/PAHJLVaAYZUoWwSPBllzZQZ+wjdQvFrJhY/rGJDiUPqL6ykjhohL3Zmn7GBzqRlII/4xHj375
eCN/c0kq4O71GNzQ47dvrABPbrK2MA9Ho5PO801j3cWbWZaPL3sjzMo94kzZ/j817pitNwiRGLzl
DaXbEMzupXtgdBmpE7nJBOh1i8ZIt++z4MpWVoxZ9efjlan2cyAxHo/djdNJzNV7MPT6BKafDkPz
YPme2xqhm2iUzCanKkAhoWJcubP3bGG7OQkyQMd56qMm39mRG+hOS7lSM3pkalNFi7sE78entU3X
LGObnaoGf+ztiI1ZZ+l0Am4lb5eM6mG6GgAsfSQox38hQ9xeQFJUYlEYmzGmwoerTipXFLgqV460
I1797h13mJlMCggM2y3+9WNIq+I8FhqHqHcZnZcjnW8twtbIV3SEacLYgaGcIMakk7TSSZi1coCk
WLNPPnoqgB/zNdfnQAaW31HO5J01dGYh3GfoDQCTMTzFkR4xariUceS0cQVl1AToiEEFVGd+ywGj
d07aCDIvjHntLh2zC9pAcROfllKsF/lZHITzLaCNF0cIrOVmTZ8WJxvoGI3189S4GCsORWTTr7k1
bCD1OYIPrHxgaAKRa6UGY1zP55z+8uFWF6ERxYrG3ACsC4EAAz1TnVirr6IuLy8LknaapWEDZC66
fBCVyfxLKo+bC5UhTmEcKrYl0H16X4pVZGgsJLBe72qnE4qiYrCpkQXNbicoXuGwZeSqNruYaXES
Xq5kslWdl43GxRivzbcHiRmkyZI3xx9BJAvi92QIE2a6mMImgSXkFqnVtkpD+gpGDzIEpsWoif9B
hDscQ+jcjq5c+KPx8G4E5QzZn2Z0nuyQgE7dWBzJIVNLlQKjSuXJsQty7R3/YUz4gHh+Jgvpo0si
Q1gkIbWFwYpRsIlNxWmeMcmm5q93UAnnwmrwpT9b8XjacdABtAbsnjLxpxKSKj3XDLiApHXQDrfR
ZxN2Az0QSwqYUfsA7SAsLz/A791ZQSamlJFvI4FcQtzSvzfqp1el9Hs8dh4sV4BwH6Abc7eh/Ecm
edqxoyF/0tJfIKUT+bVV4mWqjY4ZD6AnS1vXqmwlBWsVDe3NSD1+zmGxjrrM71eVHWTtcQP3WzxI
d3Nhd+//Wz35eLnb7FP6IBVPzOgd/1lSgNdyHqHVtf7eS79t3k/UO499kLacOgdGbZZnrDV7h9BL
uifMtrQvLjy5HYO7gqBFsuME7RwQqm7MJIJUI12gU4ozy8JARKwI+Xvcrv9gPbxhZVq4bKrXL069
brBmv8qikDI1zDRo+Ucf30sBzKxU1Og3uzmgU32VlH2e7+KojLBlvJb2iZPL3EDvjl8ocYDb2qQL
+/6j1KPQZ/hCV3C+u7PNORlUFfhr4jfx7s4dsP2CJtw61Az0HvAdmNSFxTfS87eJGXq6kwOp44Bi
QmlukX9BE+41UjA2WZQc1ssWqLacd0ZEAMaG1C3734mN7JeVVfQCuU4zm51OBuvz3jrQCem0vTR2
r2f6G0yAaU3fqFpJ22p7DMf+QuyMDPhedAdeIbtVtaI+6Wt59TWwp5S+M1b5t6ANae7dVkhnitb1
JFXR8o8eYjAJJlnx+O32ACmdBVYhYkPW65oUlVbVI85cy4nw/NpXvG4EVPcia8T/EmUL/9Njscjd
+XeLgFzuB90qpJBauBnLkfMdsJR7xIb+yZci1z1D7+qdkfrsC40W5gMMQ3Yg6gq4aPJktIkxjhK5
METbHwLQ8AojmLIzR+GixOtObwK9vugs0xb6wrdWViEM1p5egTEREV0bHlOxdc9Iv0DGfeNbdy9L
1b98bYL5W9Pa7FyXQ505T6myehNxDYMemcIfu8y+5wNWhfwD0InYisjG4KFZxYzybms+dzKr92/j
lmYCLppwUsU29Nbz2PQTBhAJT5s5oW8wwlyWCOrD0JMVI+iYd37RJurc2PdVnCe0lGZ0VytxyxdZ
nCoQQbgEIqwhGQl/gnrqd9ID9uCMjEPEUNJ0m9SWB6TA/ssnUot9/nYfGKDJc/DOvrBCzmJ3DCFh
qxnPGHZSiE+Tlapqouw8ekk4lzhSBSZJ2j4rtLygoUxhJIbaO7X49vRU2pamBvw0bDroVJjqbo0l
lwMaZRuvia/JW28mW90V/12zKmR0QzEFIsm/X/ncfGExiOyAR+sUv4Fyd/WpYkoFRr68Ysa3c+wa
3fhhkQjaZuy0X/jWPyGPzRevn8SKsZRSyUUtTb2MCUCrD2eH1Mk8tzk30CEOd6ZeTT3YkdEAMU68
DQgd1FZYlPxZJt8zOFXSUWIfWB+3HKiWkSE3tUeJm9BC2z/MNFcvxS5txt5VQbtmO6uScHlQZIEj
RBiOvHCdDa46nBOsz5Jg4SgGBzsy28BodyQn5y6H2vsZXDOgevgvKhK6t6lIBgbjxhac0nznd3W+
1k0EgJ+jPerjwiAu7ViG6pWRmzYEU/8NZoTM3fT8oxXmYwOk/EwXGUn0hyR+TlTMCftNv7gjNtre
JqB6i+0bhwtsaidXh+wuOuNCpjpHSmXCKucbr/lQ0jYvv+l0aC1NE12ZWA6gF+qNLdkT7WKFoA90
8QkIzUYyUssztM8kqdgVO9cZZT7eHg++qjtDAY9Ie7zc0gGYD2i/e94zGfkK6MCRU6MnzdFt25zm
T7l1tru8NIJqNp7/L7CXvWAeqVxRIDzcleOoDvxCbC0MS6h2NsBaXTUHXmiSjVeGsBsYQAM9F1Zj
n4UF/PkMvG2qxMJaw38TEQiRsFV89o3FXSIKvu/w9IBJErws1kXiT1ayKXYRIukrSYC7N0V/4Ek/
0OYZWgGkMJkqAdRrTPkq0OHQkH9QtwwWYujGNQZCIOTPeKG6SyAHEBd29qDsGtnBN3fduGcOEqcc
PDjD/o3xVXYhSvpY4zS5g0Fc5SJwq+cMm1M7P8IRBJDDxfGRxLa4/xEkMyDek8pBpNI39rVrMqiP
PMZrb3hGMgn0s0eCp8cAey0NFoxVMBhcth1Q4zGKCLF1c7feA28JtoNrco6oPJ31VRU3dehCzkJI
8uEld3BGNO30Dv/FxDfNQ1FdT4fSfrvgFlMu2/kgPtERBwXlFXFQpgXNeHusTPkZ2jTOb10Gz2dR
wUfENXXnL1J9mku9iBUzTDnH+ZZhHCKBc4PhbmIGSFLo5WDIMhdJjd3T3I7VibIUuH6gqCidnrE7
A+/ZkeuGFQSjypkCxYn43l5qjcru5X0zWDm55LD6C0qaCl1BCze721enR6JCtsMo/5HVj0KIb4eQ
+WLyfzJDHut6gWF/f+I53tM1C+5XroqkgAlux0CxQ167hPH1cqA5chWE9zaRg5LZn30u96TNIBLd
adgaOzR7utyMwMSqDCKD3pxYjfYo8UexPUi4iFoVoeEhc1nH4yTtl0ysBjCnflXnN2cnJQtk+Ruq
sh4nMBUIohwALmUpjcmqM5saxbjciwkfADj8JH8vkU/bB2Y0ylwTGcFSSjz/Vz3z3z8L354NoJ8N
P2BorT5bmSwy6xmypAQ3n+ZD4H2sVDdQKlDWKoWcv1no/zKSOI/cZez/dvA02oiYgASHLoqOr8MW
eakkW5K1YtCqw7MSp9x5Vu8p6LENrZS/98IXKBkA5cFmg/BF7GXcUpzD+cUdnOd5PiYRmxujw8I6
JG3hL0tcSgRsGZytc0U7nNoTzHYJIbKhklFxvIvP3xhJNIAPzraCzY7EQC1UfYeMEZH9iv8GyUBE
yrmV4V7lAAepqGR/gxSIG2O/eMMxFqcTNDfry7tJXFrN7oCeSwu3rDoeV2vNOjFE3qV9bJOr+lAC
IAMdXzu/ZZ3r9SbealnNYb/HhGn10ptRPt5zrVf45/OFIu/y+lChQc99zs7QP4L3mztmGEbtfI/A
ELzDBcRr4EdO3PiJ3cXp/+Jrp9eB4JMCUdQyRGUQC+VncAm3zTVzRTAe0GNWgPHlLZVQtsHgrzSK
3HhVpvUhpFlL3FIP9I3bQJySxtkfOf4WLAiiXZFcGsTgrZjF3lcNa6BS8NDASVjP4MNcj3TouOZC
Nb7ttUV23Z3S/uAbfMW+VIawcHiKEjRBDhv4HVjOdzDIEmrggXqsZzsI2hAyo3N4qme+EBMgmczu
PTZu8crZ8HB6IjC7yzZ5H6+1OpukqAKs4HGq91vPtl+vKH9tBm4nPUpxwgqtvCIySIip+3lhO4jU
lzKUx1oVn3U64CjD92QH0edCHbfS19E1opft2x6Xcx689etuL1zsTgZ5SAx0KnmUK7Wq5cRT/DZj
xhAsF3xIPD6FsKvKy9VCHeSTeOxd6dgscX1OPlEWLBwlK/wWv/jISllYEeqVJ81hfGnZDVm7pZh9
YFzshkF2EvDFXWdj40tjbvYUNDEc8TGefGOlTkUKomzGmTZVH3zJSHoW1xrSz0OAXQHfOw6gw6vq
Aqt1uGYQC6bf/3K5ITNZdNGD3c0vs6ZKaEau+t8h4z0Hx+NgNSiBdpP7YbEtHNgJESCWTU3EZUXE
KA/Jeok4/HnEfc4kNXqaq/NwrwKrFUzpiuEFQ0v//N6LX+Y7JYnbVM59/8RHUqfz6r+77n6F88BC
dh4NCSpgIsuKFRO7r6U/JgP1iKhBTZFGw/DWKhrX9UTDx1LsMjOOSnS8/Hi+sfQEVwD1Bp5/RFE8
NmNLTQB03v5HpucqKinbzIZuqkTDvf3UjgDDMzXrVMcfeeXEFyfn2RL7Lc97Vlq1gZfNrW6AvUhs
klRmcsZB26o6ULmGl77IARzu/3FfeIHU60Ba15YGFSWuK14rI2LR9EeLny3BWub/LNlm2kH6gkj/
5UlPUTHGY6K037wTwgJU5/z6Q5I3Gm1lpg68q0uQOB9UtuWTYdJW2IRz6aUWe6IJwjqlDBPZSwPk
+zsoZYlZP+UucZwsRVxWSEDmwB8Ve5RodkuMTaYT40XKIz10QgZFzfRVK60VTR4gJ5PDCpICf+Jk
DtIPubbZp5CckTx/RdeOhRli6au2zSZVYwUwnKEREL3dMboE0+6L5m7RQXAxzLQT1o8rjrm4GApR
ZhFEcbFYb9huB/JiC7CTL3eW2CuAEL06FoOB4hA1rO0x2Fi4NjdrM1kGMIDMQW5n0mwwDRHUI1b+
62fVrGnXRShApjxzyzpUeyCp1hP6z4OEaJLVj8zAH63PwvlkqIYld2yW7mXuMeSD74oXEKBn3NBb
4fYEbxLfphh9mYijP5oKLyNlVWJIsqIU20A7baVNPNQX/yYJkwN9XVsX6w1Ie/R8ROwowdZfJgSZ
Dv2mIYpNc3j/L7opztyhHHIM0putZ0qKoVJeJZxler2+ewh1SHPYgb93v0kq2oyU6Tj0HPrWxuVg
BZLVF1sA4iB+i4dS/Cuqvz0XRzolwH2AlNyaW26l28Nhw30xZGumKBVTT86GpYyGYfugVgmKWHlz
4ZN0GXQS43n9bi/fuBnRMPgffNOpPyPi2CRxcqba0fpJ2JK44NxbrrjzsVTh+yFCahNxNOB4miMI
hQJ/eE2W9nR7z4NoSIuQVf4az7DEq4uCX2r0nn878w/K/hb/Bb1q2uZ5TAlYyFPtXqN9H4AWOKiu
CKVuBadLvJb36NDpiVIim6lsAgyEt+RP7M+YVa5Xw9cRahp9KP2KD3LwPUiKcfJoyD8nWK7tg5ZO
LyqQA5k7Q5kphDyabTbRAjZjGtrTPpDdV0SdbAQdJMana3bahYZ8VsTD+Q/0oHkeEOGPJqzC1iPq
nKmhPSBCzDm9DgIsqPFaJRYMGhBdYRCIWSFTHlmZP9e/SIyLgnnFbV4fqe03nfzykdHWQm/j7Ywc
egneE3k70C1rz8v7hYWL8OmUDmlPJwq2qrjykvAQvjZ6WPgIgP7/LFRObaGLb3F+mHRc2PqnUzze
bIDzEHXJ0gwkn5dFhZUl+K+bgwIjXOFKGCIfPORTQ+1ZQoUrZz/l5ZkjJz4tDJ1nggK8NGctkeBC
iDkAIPtyQkxvZ4/M5DjoVnQaA1K9YLUNB73uyKnWTojaRESToyZ9ijHPunhu/v2+tJyOKBtMOsU6
4a6acPPy7ndxfMYkzVFbRlghRMI8LrZf7FWYHIoO7QvxALECo3hVPB5DQ5D7XgAsdnZCIOzJqew1
Lr+Ddhsb9CRXGW8MiyKpVUefVz0sQDS4vDTNOwARVz1BdVcxumHKrJFVcCV1v8uB8AGYQ2FvZI5O
ncEhq517JZIFR1+WDP4IMXVBzte4hgcYAQonZBolJtHVIQO/eadtDryD4A6XH6XoW5Nze9etjFzn
N8X5U4mHmNczHNSRbGR9LGs1/3JKkvABx9GNyQbqRlYvBTQA7YNJMu3PVKlovt6K/kw5rUFv0KeQ
4+7YYB1uwq/k0z8DBw3qStZ80PMD3fa5Z+dn7t35Zbt7y54hplAzEKZaxSjg8xeJUPgE1o/hIMs4
xi5xmVrHnKV8EbBVyGN2q6bUegWmAFOKLHIik12bFI8usmfadrbxcYsaO4fy90ww/7b+H2y6ry4v
7BkU+VFS9q8BsF1mn12wgyCsrVF9+EXBgeAumWaiztS7RL9Lbp6epmUHh25dLhY2kQ5nMfnq8ms3
DSb3mve/7yPYJPchnZfXtFNdQQoCDAikYZ3+Fl/q9XqUlbkbJxLfu8UHn1dqARQU6YXYJP6j4/HC
PqIVAPBo9bHI3R3tBjSfAoWAHSc+IQMsptmtqimfWWg7oK+23lP1wW6JZzl9D2xuLzr6HO3/3727
YYo1r0UIJ+I8YpnT467R17ktrnXTuZOJDFNvn2KRFwdTg7XfhUpvc2wUIAf4/ZZVdC1pPfGQRSAB
4Sxs41TyDrBLjpmG/BqNnOA0WuJSQJq6maq8Z2MlIfuJBXBZ5K5ltgrqla31eP7ptkpPaxJg69B7
idOoZC6F3QkNcRxpAb0L78n/M0hqOXi/7Ca00Tf4GHB8DcXlbMmItX/4SX5cMbu2ianOIfkeH0sm
QpmdUJdnk9NsOVH66DtRV7N+4bP6lr6x/XC6bF96vXQVmMiXonoLuQPOrdxYSpuuMAn2vypeoRfK
z5zgXPdJNaivIJHm5395XZTmdznohfLZMux8ysIItsKQfh1NTGgNmPejXAa3Ppbmnz6Wi0hKCaSR
U9TT7XbS3rdxfh3P15QXV2GFysXJECsQykYMQ3XIcXOCI7vi1hfTUOgZY3uAP3mMM0qhYVglThT/
0UXtyMMFN7p6N8SYOPCf4ktPRiBMJxUZvOWvM4E62MRPUAX07pdlgX1TOuDLI+8MFUE+XHsd9Y5d
WsiGtNEf0ejd3e1HPP4hzSCyXYTT7iv3NZ4KE7LuDnOzALAkqPUEwQuUUTHOTJyrJCFREXEC/9CS
94iVTCtJYljNxVLeoQaqKohAMq+hMxbA+DwQP+4RUZBV1sHq41SKnFz+S90h7ppa/CWFFAUYs1iS
FZKeSPd5kYjBa9c9N2S/FYm9kLFlKd5u2af2aP9rCO2LbkFenQfZGco1MX5tPmXLzc9IvNaBf0Vb
4i+dT05P/o2Zwodmgxgc90UIBXjf9D3nyGAPHIVXe6t2FMbLu6P4gl0imNlpiJNVshQvOqHTpXTY
80jQijrPRWH3t/uCUK7B4PAM2aU+WrmiVk0MW1vc20Lmba3YLvqCc9Ebov7wfLwZVE0IoejOw0T4
hEUBBdO+LVSbMnXpeaKYnIHOK7w/2oQaEg4QWFHahHZ3cI6V7+UqIa6Sq2PYt5cWxFOJukJoD29O
PNXw8R7gTxVq2CCRXh/vapTtRdAOXOE9bC474K79AAeitLIA0ffEggsoLLg9bB5U0/4C1RedX/uj
imnD4gOO+1hwXc9J9+DL0esSuHL5tB0FKGUQsjtU9iHVWjzrjNiCnIszlg4NCc64nuXqfd+rtMa/
JO9HSy+az780AtVMQbVz4M2u4igkZXZTWhTQZuO3kPIb196vD7F4OzNaVgsJ1S/arP1Vwt0U8FNd
dhIkMfS4TbRcOTJyGH0JKFCHMUR0xpBgAvBGtldMFu01ZFjnAI1L0b2LMWQvBM8azOYrC072eNdD
EMU72bP/f87Eo5utJEOGQaZkR9jrx5kftF4qQWbq5iQt0QlVJ6EDC6QMjhIyY2X3Sd1GdbIfo6GG
9pUdslNSlCQrrh7Z4U4KESfkID5lmF3M60r2IX0vhUJBZso8MiuCFUp8AZL0ut9jfypE8UTmmOqr
xYaJIeXbWS8HFBdAOvfVJugndCx9RKAGMBkKIwZea7//KT1RFsTpupf3r+tWr5yBQrB87v6KPad2
rbfi12PihkIMnNkeSjZaAqjpZhOJ5IKTMt8s+LJLXqnRbLsYZnRgttmT7RbAq9s6NNlZVe7yX5hc
V8BEC45DpX3u8haM7Pdi/eo/Z9PsHewu5p8AaMSoSFfcI9WDxQdkVIhJn/07s5jbMApMOgFwF884
OtWM8QeuzCsjXHJk5VtadTPFtJ7bgGSKf+iFtC/+0dJBMe203fxxEslp0JjyyFQjSRt430Y24vIj
yk2GtHQYy6436bBTGVy1eX8A5A3CCBN1YH6hXvWTNpy4OQS3VBqsxHDzAimcx1l+Oi9dI5ILPBII
jnlIxRjpZhGunxeOwXmf0K106/Yy0plBuH50iUUvzVcCdJRSN+HEnnlNhwEvj6TARsi5vdlcR+79
rSyIFtkLBS2WV80FQbwAlzcYRY8KHB9hqPUf36AX+iByi8kd0waakAaTi4PEVx6PMG0q/ykraTQn
S6GA3PYbnu1/9Xr9W+DXFYRKaU+yB0VYN8aYkNKomJjYgZFptGasQ7dN3wK0s9p7IWZepAR6DgQy
3F6PPEH+/ttVc4uSGrKyCQhVE20aXibn7+0Fvc/hapDtkWnYA/p96+te2yivvmoy+FjVlKtVezb6
NbUZEwhb/QWH9IZ3HzujnHGCbKgkUJVuwkjew3LCZ51xcySrNjD4RuYyFKSepQshjljBqk8aToDM
OrV6AmQpttZkqqba6sYPXjlba4uWJKlqzMrziI+GhH5tV4TmjPow5am+b3djmljWlyPqajG1bq/c
rYRf16lFIHTc97n7NL5IZyETBIpRvJ/7miSGmB7L95DarwiQ3WI0vVL3gRhdbo31t3NKe+K62VGM
fkepKoqhrb25MUcc+TICCRdGyRP124tYDWVKKqPM1mCxHKGjO+hXe2zvuKI2ihnnYxzfN0TYQiJX
cz69I2ncIL7JneDFOC50evceCcBNfgViwQrxWRJY/iuQaRgQ6LiQxFNmzASU3/9vAYN6OVa9ZW5B
8TjHpbuH3p8+zwDLn6/sorZJdndAa/08xidOV/pT8+ksAwo5G4uu07A5kcyCZ41zn6wkzbIwXJ1g
Nad2xjvnHogXwVLSP82QEyjvHdRTH645hG03/8lyhktwqF3+CVMA3iU8MMeu2bhk6iHj5+pQ2aug
69TkNjNM1M3SRsPquvcq3moj6YjUn/B7pU2WjSFB5Ytus/9XrppQxkHCOq22dJY8iWLU6ZSDe5yN
hIx+7tbpb5587x3RyLh4V3PB6Eclta/mF2k648SRVSQXMYKaHpc6Z6b/Jm7tw/H1hERMHfA4I54p
N1435ebwOYvP8puMxM3m9HFCBJPNJx17kGML6yGcWB3O4TvlZP3gQZfboKrtVWK5rhfW2a3xVkdJ
0Vqz/hnHGEcCHd0OtxgeW26iISrSgo2PafMfu8sOmxq52Ni1mXj1nwJYr9LjSpU1DAc9wL9MwI7E
AbBLSjhRyNB5WojYjesvx+etF2XXtxJPjywgt/E9iSx6QTNjdwutZXBXe97tobqxa1FurZrmzMDs
z3RBzLFOQewgomMHuniGMZEiq4gmVSNKF36lxc4SFRW4bFtGd19jtOHoNKmgAdqB+erbDEXc2AA4
QBSwCDD6x/46KQP5FQNChe1w4ReuL6YVqi/i0PgegJY2JB6W4SXF5bHQk7pJwFsMEZiwTR11kXPI
ovr9mb2afhGxbzhxua7cap4z3YeKttlrF/tmBZBr5SeL/aaNy154dRo9UMz+cxR7177Xdbj/Qq7D
fh+UDKlWLpUvSTIC0ZXAJDVDXdGwLM4641CmEjD6xWVyrmMhXuHwcxJqMd50MNFU1cjpu0rk/KIb
fGJaWdExkRmtGDBZLrltSANXdpQKsuuOER+SrQdkGgsIDrBXNa6qUeIdmCi0xJXBgiTIuR+muiXM
4YuFbm4vpPG+RDd0eEzYMJfYtjlj3BmhudCXzhJEGjlv0kOCkkJ6ITUCoV5vxqR3Kj292UvtaEkx
Im/FR6VhtN4JSyU9iLIL0sN0E2vxLSbuKpq+DAAyafcs5YXfOi2CbOWKy/W8uoqazGYS90YQyaJR
LPSq+vFlUbuIkcQnemytofOq9kxK4cvcmsS0Y/vTNGLopOSEDzZ3miEd1tB8vLYDIpVhofdqBA4l
QGFcoTOPvS51MTIB1mQN1eDw1gZSN3WfjVpsmHI29PYb26cOSObByt8h5Af9On59sgzNiSP7xIVF
eqIBva44POOANz1rLL0fvq+KZlUDMQ3D/kRSUIw4aQF3gcaQMj1/innBi3q8AvtTibR/hLYlRpio
pSpZaCW5oGq0Ezx2/9bDufLwfBN3I7iMBp6r1wNC4EexQIKKLaR5HzgqU+zLMDFh9XZbfxlmca6O
ILHPUsoTTWTq8ly4d5NO7TLhXzr/zDCoDmcWhJ9GPlg9oC3qPAHrVjTySwEdldYnjaWkGJtA/SLV
uLVxXXWZ0+2Vh2goH/5OGqsvjYcczSxyF7MhHQIgh8q+pzuGQUZf4q06fWMWKMdkYuZba9YnN0T4
36SacGPwDI32LLzl6kQKhRKtdNfoze1NGP7j6bSCgnROBlJa/PB8Tdwz3YoR/kpayYeeWiQIddBY
5sdrBTi9IWyrAuYcHw8r6SuwsQSiWg08WdFM15aH9cLehwC0yBcwMew1rH/VMY68uQHtswQoMaOo
tKD4Gv3QoEaA+676i7C2jVDc1R9efGPTUeTveYXuM6LQ7ykkce6/LSzUavHx61zff5FdJVjvBBjz
cGK/QO55qUoWapivbByHYnm5L/khym3I4kQ1AfE1nS3pHn5eayDJX2AuW7Ab9kKiYTw27zzXEku8
E65QbaCwdnCk6Pzj3+DovoCbnEwCG8aY8C8DfiLjJeVvWTb5+HuU+NLLvk3fZnqaLjqYPi6FvkvL
CZMKWi2JQLcmti5rxqHKtDHJ7fpHNzBF+7ZEdmZhVAwOJYV00dkRQnOydoPMjmDsnEXz21z9ns+1
pvp1K80ybigIjIgnSvwsc0djMXXFYQKX54NsdAQ8qHg3nMhYQL1OsLBOVS2otcKyeG+HqlgBtQM5
hdwSpJFNCOAChq8oe22ivzUTJ5g6TJNfb3FMmxeNPSDZi82xzZZM8uhUB4YWl2ihWRMRtsOJYxDQ
+VpF/DewOXOI8JCAZQJ5phbxq/Y72zfJmIlhmvLhNbQiRezlyOBYMFVYLfaiDoywtBET19bACOjD
mzPrvSGKGXlobl1uZWBsP/y8UUvzWH3lUm7xlzo1je/ouvCVu+G8TS7EKCcMiM8Dy9lh30BjaVpI
S26LxKLOkgddQ/l2KKVZOXj5Os+yC0fXg3bUAc7kT6OOznnN+hHz//FBQO95SfptS8aJCMLKS8gW
Z+Om9DcipNbNTMcfXl5g/mVl9c67IsO4eko1XoRqIPajjcmGY8KE6vnfMOL4VtyTQC3+rX69ybI8
Mtw7EGLS1rVQtZhhpSpSt9uZQBlfEvu+hJMfx7+l5JmqdDqENpy6Nhak0pKjcLFtoTT92yjxvKRM
JNMPrDYc/rGX9P3+F74RqqLmvZSkXaGLaNjKVeOLLfbxOgQkz5aqkScMdAZGTN9TFplrN6w9nA/V
7bg+/b56ufBoqTGTCTcXYxTlEQfqytoBBvWEcWtodDu4NySnzYLK15OSX06+4xOgUToAI/yhbAm1
zMb8e2XS12gXpOa0eCcM83Chio/ze0Cu0SNnANagMWn1bV44c5Ky7ydtfU2oWuday1U0OCcSoYB8
CmcbbFrooWTy5FTE3bdXN71wfI/YQ1bLb7j3YiFNTcfXKt3sQJpbdC3D4tEuXcnQxBxE7ZguBzJe
7c3Y2tdBmbVcGoOaW87GWNdVbMh640WJA8cnwPzktZ0WXniJ/du61Thaez5yO7BhQWNjN/qaxWg6
x8BkWG1dHdlERThrI8ssKYPVTow9kjFFU0aOafuVWxErQhEk2ew5QSG0jhV2zYvj4VEhdevY9GEh
kEaddAKUSU38n30Gm4jLUUtcsugvidozlqG08HiuIHl/VBQLO54IakUFpXfPKhUzUnbGVdY36gVj
Y2iP/oHGdNmorPJwG2nQ0FGIEGwPlr58tF88z6yllvFq3qGGcgADiTnZGsaOFP14Ms6kiEPx4PvL
QsQ4la3agNWv1KoZskQRKr3Zx+oIRFw1pGq4ZrV5Wdl5zLY8JuHJ5h5BJ0QoGWbgSXUBjib75zW3
fnMvP2RwdM6Jx3Jik3IveSdfMg13xpDFwikdC2uzlPEv55Yci752TQLfdDhJDxN1YuMYBJ4DRJfa
oWCaClgbbukNbWEhqkXW8wF0MHqrAeSMxCetCSv549dtmMGHxzWyq7VI9rLUkDXzS8Xdf9AJLyO8
XToFnUbstJStnhkgzoy0ggHTq8HbXSMQMo7Wi0/ajDfshp/xNHouFD+N3Xukfdy4whPYXm7WVuMB
FBtWl0tsuQD4YzOVvbGS1sU6MFEZsNZHNF/Jp5FL+9+WKuEJIeD+cJf1sBzf7S6IWa6tuL/WxGDT
/KkvAxklWjdhV0RjlWYk6+jsrrFX+RqWCNQYhl3gsw1Yjvp+hj8YAoZUS1mbheF5P88zgud+hrBf
kuLyuTfxHcBWcE1i/lqTGTSjMckWtAX5RCbDRg+eyACCUsNCdk9PdiVZb6G59PMB4XWDZoPZAsf1
DMZuVpaIe0wCdCh0QOH2wzRiw6Jwtt/NAIwILvoCOub4VAiIC4uXcDdmPY8P1lKVf9P5zO0cMWoL
+Hn6LP/1dz72f4Lj8DOXT2eZhmHTcvdivDwyKGeCgM9nvG/6MNluvICiWzrBaKVuVrSBUyDCcGqD
9jl4u7Hr+kPKrrFNeDi+373AYd3Imik7oxh8a0rEk69nHB9aKpZPHQg/DSSwd65dPU9N4SVRmZm+
uo3xdgY7yZ2lIb2RXJPvbGZEm72BucNvHbjdWvTCnq+iQ7Tkb0mkQx4pWbP3Ojfp1+bm//VTMnAX
kA1q5WAtNYNThveyvr9z5vnhAIaX1g94LHZv4eDRBWkS31bHTt1e66ub0La/xrc/IuUdYMQd3zvk
CGAPWTwvLTZvyLliizid2pohO9Dy1egWYPwl2EbdzJhUheLXGaDrSddf7zLg6/Nxptn4/n5x3qlc
GYoKw0eT6k6dIHy8Nb/j7j0rVLwmVmmx5TOqULT9PfYYIy5BbpBE5GsmTa07w2B6DOGal9c2Fpqg
9HN0Ig8XsE/jEsoNVpls8uskHf8EEocWvOWrv4IoS4NLOpLe0MCN6EX9rNoHjd83XCFX07Wlso+T
NqbFSfHFJHLkrcCaTr4fCzCxKK7N4p1sF9Mws9ueyyfQAUEOu1No3xEgnjcJDv6iHT1V9HVVXyfj
IoULUBOS/tXHT4ou5XFg0WRofMR4BkvrM5l+1WkRkIWijRLNELmK7i9CzT9xQSuok0YovDbjqgQC
BmP6xHymEjXCgFORl4vXRhH9p8xNnGRMSCtCrorgQsjkB5ePf6KSeQcby0TEaN+lHtGVww1g+QxL
o7O/WeqYywnEdKmSYpi2alyXo6zrSESuAg7OBE0ZhVPH/qOS4HI62I7zGQV8/FUNcpHJuoYDGITN
+H9onjltKMf6tv7/7gTV3KDecUtUEtEJ9FctCc/RqhO/P3NVwLLee3er1kz80afnrWrgjFEFkShk
Ww0rBAh0nOzPtYJM59AsorhkVOEIhcimddgWc4EA3lxnjYDkIroR3S9/1nqKe0UfugGmmmLxuojk
tnNJUmckHMT9HnftZOr2+OIN02UsQU5q3xqD+WYY/2t0XTeNCpwDljlmlUrTditnikGIaeki8wbi
A/hBDtxiql9xMXoRvpVvJnkEEmFpeMwDkscTdtTTm+d6hNWkB/tzcavfn68aTRxbPiBwsJGlnSn1
ieHwAnChJUGhB4PL7hBM2RhuNPR3X9Vm+ywWCvp533MKlJqv2EZJQ0C0Uoum5onmU+JYem/jDDKa
ZoVER2WxBd226Yrk9A0lNX5aAo0BMzXve0c9zpofQGnX6flKgfDb17YRRBpDTCnWKp2wMfHBGi4Q
QWEGhW0KP4FYJaodQYlv0zFUU06VXvAMjo8dBSunkiNIktDfksk+e2456cCN/hbOuilhZkRLjG1N
mxllLSUL++ZAiVFZxDF6AUfx/jrdI/qfnBbdP2cWT1+xKOrJbIVVVL8o9ZqIrs3laVrvFoc7mBvH
seURtnZtd9qTF339Tfu4ObiFPpFMfhZJwbY3XYM46RV9AnO5gLvrgjyppDAPrNeDxTxM4gwoTVGx
J6olZ6BcbsgU44nvX1YeuCyRUTKQIVsX3tBq984Y7gxhso6jOSFYBnWDK1gIG5dLq6O85Fs/QMRu
3jfN2qDZH3pbWCU1a19Z0u29ywzPETYZiBsNL7wE60IQf5JwzyvbQvFmLiXo2C/LLLy1Gyc08mKo
Lp5IpVMCVQ4mPfWPewFS/iyodJQcfz5OUQ0ZQOAFmmiFIgUBAt4mdUk1rC4TEIEw3uMPHHEBkLB0
9rV462V4U1Pr31hmAIpGWY4Y597PMwAWSonno7I6BhIo9LK5h4BFOn0UOcLvt1d1WaGhMeOmJT3P
0JUZnoiZ0MldWexVl+TMlvHK4uKhea+RrngX8KPwQOXq0HYyKRiUY59R5uyGRJ/FgaB1mQxIbBjb
Sk6XVyvlZRyFn3QX8k3RbHyspSJfKR/z7YlM5akPnYMgbsK4a0+0xM539jpU1XkkdcTijXqADcBL
DTHapydYYpkc5ce2keHM6iEjn2jf8Tk2Y+/JlXVnviYYr0P53GtKoz08DDCNnmezOUH779Mut6d4
azkADBlbQiPeln7BkZgZl6kTMkOjBxzgcM3Jfd+HEHzdvGhqjlBQ/RgnjK00raJz4GA0ddJC3voG
mwmMp7WSKYWaLa9Kd4YiqwdteAWZGMHwXRfKZfRkQjv5LnaZdymguYMvT/hOivhxXCRNZH5w3EfS
PhnAVH3kLHanvCBq+EeXTWTOGVl1eypJDYgPfu4dDcONoDCF9ISYs1M5aN9rc3AZKzcYZYeAC+q8
zWck38ZRWiWbpXXQmqumgWWZ/0U+GXpsvoEdu1j4G/az5JnPeOT1rCb/DGD5ST+iBx6gvV5cTTdN
pIeajND5/0VDz2rjgomDx3dxoZJuvX281dg7spqiOtXV9v7iYmH+1E3NUqgQGzUzpYYlsUyGKG2U
pHC9/CTPYn3iqROAFpQoexu3xA2sUZ+Etu9YhnuaPSbroHaVnyQ44wwwqERaBIQzvqo8gnsldpFB
4Q6CkptKYiLrS5Y0OnhU15spbMaU6tBYdVaOvDhMZVX90WbkIOQ0mj9y+BcMIvuqdo9+E81c1iG1
Yj7ui888mAUAJ6vn/LJdHj0kZSiNOd325fSYCqE0RMw5DhN93RUBI0DBdJBoQNgMoPjNZSVFb5hR
nicXpWV/qdEeqU5WqXxTiY/ogDr9fsbuXzYa74USNHI7ub7VzEVU8M4saG+9WSNCepIagNO39HNb
+CEiJ+hzSfLPGgXVEj+9zB46ZGsLJgFDpzDnLQ95zMWwMNQUsCa1vqYbemiVvZjHHhZsGNqEfVuZ
Jp1U6eMbeZEgfUu0XocYwquW0qFH9rWC7Qe4LLEeKUSwLxzan7sj0/QVWlihPPi/wTEwupxCXxGh
S1gwo0v/YYMW9nC5O9EreEBesFGcnHkkS9VqFFA81AkAbpr2+svy9QNDaDAuMclV8ZRaJ40exC+0
SGDHcGuay3YM6lcsUnAozFlprV7ZHGdbvEoaqi4Oa/S/7Gf2/izkDSwJSt/bECJCp1cS4r2ZOj3V
aAHUvFhFkjygPV3+KFxt7Xop7ZyKHjoa/tOuFPvwVJGNCTosJnbOiq9xj+D4UPvXfMLkmHMlT6l5
HJGSqA+0E4wanetcl0fnMZZzaczAoyw+PYzJwATJ++kMcnAPaDOaNp2TPBJGFpRD7gzEaJpyBfj9
rGjO6vGLxqqMSCjMWe1jNl6ScaaBFsqY79z31rxQwQaiO9IFsQvuSd0wx6ijePpsAbwhYr+L2dac
r1ZLrtW38ZtBn1r3LNtvIupySHOCu5a5V8eA7vSvNgGIRLr1lHBGVaPPSVZvt1yKJY8d6TFldIv6
U1+uJ+kWyRqFoINH5x9Lakonx1tJb8128+ht2Z4zQpj1NDfIjqO6WMf179mvhrr9x1YIwIl2uA8M
3hDh0160llb3igHLj89nDcSdZKPSG6Vb2XF5fe4SUidAD5jTTOcMtk7OmHLhC+LzkUPbYY+Or2ey
USJsu6HorsZXGagpjMIK/qKq+nwx+RaDBJBXfMypP54rZkAtgerVHou94ZpDpreUA2eZK2zhwry9
I3DiM8UvlzQVThqNmbqATYoXQoJLYLm2X3iLWaB7lzArc3sSMgQ6gmhFeOC+3YRkniUuQ+wUJveX
2e3JWN4xXvWFONBovZHCJxtl75PSiaXCSMWPLA3LkBstZJIhDuF/XuHghPEakPEB4GsFyRERF7Oc
kOMLg/yRM+pxN5LkB2bqciJaH+YfZdqZsGG5xAe4LXjp3EpHKHVX47Pp3i9NIjar4t9rtWMEezYJ
5sfW/UbMGHT9DZGjeKh1cImxXNBEk2D9QeV8zV2OhkPm4XywgClwddFqHeyTLQqPNOKs4Nd6tUIN
7KhqCfHBCqSX/OsMbGS05eLOdy2c0hPL8XyINCB7BF7fmmq2eANEnDJxozK2A4In/1liXyYiCPxd
4fWdD8zi/7IfMaRw/6ZKwDayTbczkOXDs40RbKFsMm5UBtp+roh/OpafURzGpCrLKeQFpatjqslw
NqfcanchFd3/KQym3GranyOadsICPiEirLqtdwT/RSDo9sywAmvU6obsCUDN3ci+2KFXulfOvgvK
eD/plHHpyBSTzN0emVa6ayVcciErvftSJK4rcreUnlKKgQ2SBo/MuAI5+PYi1f+Ask3En+7hn8e9
+VBHKJDsjB4BNPH0IGUy4HcwoUAvRvQxIHSAJ8mkeuB0Po2bdhtRTMaqzOeYRrMxRoRMOmpqyuXT
Wc77mlwISG6eWpdfDbSkEBznVgv8ambraBKQ3veqZMeBQ3HbTMZxWoxWH9BsWct42MoOt2Il0fpF
TVayegM9+73lw9JBlvBsVzeycosyGx5uOi2FOmcOQN7FYj8290KYQ1EX4gPVbY1GaqrA3Rt9xchi
VubkQ5hjeS92pCOQxLLCL+qfZMojthjObMF0vozyRhfAKXpG8//m5EsYM/3NLhU1GuLfC8JNy8kj
iWG48GKvXsFZ6GKfqztpF5lEd55UXe4jYJJFxOsCpOWKKuQN3gkoapPalO/pZajde8nJYCvqZUlL
KFNo+R6zsAAUz4lpOXB4pFqWPyLxNhlnuYv5LvYCh0ThBbdbxbGsACnQTOoymg3DPbxdk5H9krVj
kmUjGKmCglFInDgTGMR2mpYYiKQXqX2EUbb6iuFANXUgBnODTLPiSeT49lnRg300bsVlu6G7snDo
f5posEXL9C3W8v/yCquYi4RbZ0Ye/TQB4aD+eRcVfOviO+04TXmVBFW7U/cDA3tgkq7mKMxwJFBK
WGaC7PIzuGEPYbwJzla5MqcxJa0vKjzKgdWTR64PTqaI5T5dKqo5BTwO4jsUrEUpXPLXbSjoCMq/
i9QcujPJlHCnYoCxnSLiHG+W+NEWTq8gCtFOxC0VHGrb9xTFhTnUh2+S2Gt2lWsuXxcRm9PfZMEf
68eNdqZ94TiXyPmrQWzu7yVPz6V4bMbK7EKSpHrQuPiH09f3AvDXCR26qABeyPupnAWqErykS5iK
LPQP4cAVTuXFNqP2AkJcM81HX6G/bwNYhK0x9fI3dfE0sU+KidYogzIM7TcsFiJ+2hFG2lfWj8oC
iz5F0jzyIQf0B/1ZICTXAPlzU160L5KwTLE98EUfCjdO/XQ3TIeLt/UuFYxZ/X2MFNKAMMpBeGzI
TCJUaoBzqTHsjqrQ+t8d5zbDdTzuKR98ngV2mwaZZhJuShqtN+XHt20WIr1UAqc9hgcFbf5dgppT
dCi9C5BqjWwHjSyjSofkCt8Ypkf4OXJmkhlcAMXK2vjIC3RFCq+czahx5eTn+GHXTeThVcKULheN
M5XCMofGzzVhkw0muwk6AwmiK/PeZMN8m5XL6Nvq8LypXW7Ti/yspXGpS0qabPOSy8Z6t6Ms89lP
7uH/ZvhGNhm4y9deCTL6Ma0egzf0W48bgYe32zsW6MFharpIc/Fb8mX7+z9V73uJFVC+JfX31AZ7
BrqSDh72NXBa3HoRkTlL6EyVeyOHHPN/7vPT6SdZtzgODNVdkfP8wub2guQxPPmxSnNu+P2JcYFT
w46epExm8LYSKUXzyUMqZBaOxTPAhiACM9Y8TxR0XA1z5LUqFlx4HQHDWVRvs4P/aL+R4g8J5MHM
6fxrO7jnh3sBy9B+N0bzWftNKyHEowpkH9oOanRmxmJKPvcHGvUrMI+LhqiFNUk6oyZIEET8Tb5b
VdG9D3zTxwSpBID5qbcQJTuPwEhlP2NsKsV7tHN5pW1psE/rVkAwt5NuSDpwdswjWZJshcGtDksV
rlo1DtESY7mpSF8cTPBuxW6RVKNjbk6ONkJ6FAe3U8xfnFIag2qPwsJGgd8QOMmCGUt56zvP/16Z
WdrxhA9a97dNUUm33nUqWsWlhfRZtVJSp+fMr+owtarrDFXB53rP6Jj7dC0e03z+EC0o2onOKbjh
5buiSG7alRLKnxwWexsrxCysv01MY7PYKiI9Pcubdc+ZyMKYW759fTlBkv2gmdc+svATtSti0Qf6
mi+7Bz8Isyf3m6wixFh7lDkIpQRcITOOHAXXYEpgK/yRTlQMs1wv5BJymqCZZcCRp41k+ECbogxD
PNcd21Gu0OIiH268K3yVC9Pn59dFilOx4LRQ+BwRFlOB7gTWihOsl7Nq5Pi+QmUu5qVJAEAAkSuZ
SxFex7sseptCDiKlt6maeREcXTLEihc+Qpa6GJvucpZQ2VMjIk9l6uJkP7oQMi236xpH9OyYwDO8
SRyXbyHDC/3fW39qq73qFRY18IFoRY1L5NXMG68n99oBgPjOFaUMJqJhQ77tRDP28LoaqxX02Jdo
aEFZt5GH2MrIrUzf+oUo3dB5By/kHO92h+5VviM+gd3F/aD0cUBdT4y3UW2TpJwGytHy3mOX5qd2
Ih2iwS1ppzHq4fIVvRycARdQYxUDeJxN2/b5lfDFH8Mni3hwdl/26TyEH/kHUrnsdBAi6buRV2vG
fqA3mff2/DCqNTU+c+dX7Ep0f8d74aOXsgXyjyzKCsZ65MeovGjPp7PuRY8Ey3ZgoDdfNkIVN0Ym
4FqUQ3yYH34tP6DNZ1knrjkjLvn2qnw7iGoB6uaG2OCAtpNqCwD0f+PSBB4C+L3lNCbzaHkjyLyZ
zZZmfxHQSuco0eGAcmIYWK3/LPTRPkWw4uDX4M7o4LOq9NZFlOQUwfgjcXVSReiMWPS6RckVN2Bz
McZHnBjj4/PMyG9yWCPyybcWaJBcqLb01/3EdA2byS8dWO2ZD/nLjTnKYlUMXkaLBrroaswtRCfW
8kuKskTI98yLnoEquDeQfGDI1js2/0nd3fyKU8ipN07fYlYP5gumX31YCdRpkNbQlPx3lSG8fwIN
5UaY56U0m9UqT7p6RMlwJ6FTcWZLz6UPvgQVnnx7R97TfuBRL86PmOr5eFNst/38Sq0IL/CR2jQE
vTDLk8m3HkP8R2LqNjOxMXlv3la5F/IkfcOTRXDR1WqJBBxOUGYgavCXY+gvPPq2+Ynjdiw260tj
ObGvxUP2lNHckc62GiIWXnZjscbxRYiMJxMQ73L/pm2sDjNwg7j+h653BnkIv/y/kM3lWcJjIFza
OfY9YodGQj8+3M+yw6+T2IK7lLc7nrfZxpKK1Jc0FExyPpjqVdfII+WUZ+BmUPzSMXScUwVQI5YP
/wFy8hso/TuatUgLIlv1YVbaO0H5yZhlUuEFsRKl2yEAT5T6TUqi3CvJWAu6jf85+m5UfdYEORrJ
8ud0rmPfVciZGHbkA0CmmeIaQgki4yrTmJh4fjlqIwOdqAv78v8ozG2bHgnw6L23pH4s3xa26vdW
DAbk2Vm9TewtU/qx5OqP5EZW6z+/OA+N/I6J+qyAEC7qejgS4t1R6N5DGHqpLKmXKNoSQkRs/QQy
xF3t2jmjicEbGXYnX+hQpdV/ubm0FkRl9UTx5uS+j43sEZhYxOMjjwiUtp/HcPOp+27JkTVks0N8
kfQXDi7EtUgM274YFJeov7fKd6MU/Hh7NAQDPJruCQ77S86ps2yD+IoZQsZCGJE5gh2jvhb29L+2
QfxKgmBZKU1yAPYlgqlKzEPh62x54z5ydhRkVw/aXe70QVIrRwGKxRgE1PXq9uTiPflzclHy4vTE
w9S4PrRjsHIuHhQlfX24h/GlKtNB2X1tTsVOk7GW5iDtGP52taNa5BdfKqMXDhL9Ybar+xVFsH5L
cHaQjWwP3rPasen/AnTGA7W6vkR87kfRt5dJW8nNiepMqsQ1lI+Ktp9f2KUBxSZxTbJds0GfdiN8
3YNtgkeYYzgOdMh7XPw2O0ykMDHiHibJAJvyAqUgjkMfo5nypZthPjn3C/obw1/qfmsCbVTEqoPm
CG45Ik7LySk2o9GUMwj1TWU6LxxNoLQTdGGKuSwUnok/cUIkonlD/Qw7RTWsRLuLKyptkz2uzUEJ
upFmeBq6Qmqg6yMVR0SscQiVQdhQMtzB8aPd9v9CGAzeR2goKb1R1vWIM2oL5MEwNJ5BXTR8Y93T
2TXAFg8eCoiukpYzsXqTfV/sS6i3g+Q6/uqbjJvbyFxaeOStk7oxzKhOItKQ3tCWsbLyiBPQgsaF
kd9jr6ByqCFP82flntw4+RotCSCg5DI5i0+/68p1/DzFj3E6Oz8+wjDtdcCV6a5eafgDLhai2QBe
GTGzE0gtaUMMsrrJMszno+oV2GCFDP+faXcyWQe0SHJsB/fXEt49DzNTlSXE2b5NbL7Nqzq0c+qh
W92DFDyIDokT55Lb/1MzMPvCHobpzRKbS+AZa2Qp2BSCZ7LAf0p11lr9j03frV3Hicv2z7ElnnEt
lvZWo6B6yzrrHsjY8a55MzyD88CAD8SSIv+5sdYqiGaa6x8LiSdqu+unpzInCozYtEsmVLRtnziu
ZVQiLqGbfYeMhSTVFHMgAnQiAFMrHnorjVQ1azGN+fFDoIJBI86nFpk+ASEeENIaWyWDqi6wRHac
0zAI7yIq9CQqxA9Fz95d/AHeQT1tj3qDflKYBsQqoKLKn4qgvz5xd+76IR4/yB9TWPT4fj0CxFVc
RQ89l3krCK1qhHV82NHhqgrHlBfgGfmlSJZ4TWm1B/i2oBIm+ySEAIZSU4q8eXGifNFh33to/Eec
DOYu4aNkJAnG3pI0k0+cGzFnYJ86y21WnKu2xlkv5HHr3Q7FtFQ38yCqxsXh8xLDY7b0yvGrZMdB
uX2Dn0NB6CzRsZLReWw2L284KMKK0/r1eVbUbGBUnVc1AyMTO//62ZDO3vKHRqka8Kvr1bT9dIk8
C3WNEdhWxC4GfuzctgZ8ajzCxnDP3zlgTVNWPGFZzz/78zp1FUKqLy8IZwYpeaZXqZ8I9DTakqKu
LGVvpTLKLm8uolQj0Bsc9pF2bMXy8eVWrxV2nioIPOB0cg9R1WGFwufclic/gZjWUKpVCWaxL6fx
3S9hH9RfIt4aYFw1tC4jbmTv+HDDTG2KCnfIrnMkVKyl8/GjLLUt5ubFnRWHlwtTjA4y+R2Vukm+
kw5DyXOr0798gK1RU/u5PnoNItFtTFBzn3qd18gzkvm2N2XRrLvcp9KgxKNfxf7rrMb8vzleAcIx
lvqNyzeQbCS3UPDqlhS1TUooUmg28I4oy3qXUXX9ejPnV5DLz1SPHUTNuH/fN46w9ppgSS36GDGh
mXa0A7hdQlXYQJP9FGhzv/itm/y5m43uPCtnmI0/Djwf1jtJf06sTDVIfuS0QlXpnB86NYbswBLq
aTiFgLc5acQqHA4L/Qqa7nJl0XGl+7Z8n281LaIUSGYXH2EHV94+4sF3UOoomp1pJVXUB3kLKR4y
/rBwXGZJko5Fbgo1rYtzAmIyERa99WYcUykFJmSUldWIhiLc/w38kSF56TcU6tbjQcIBlARBr/OY
yoFwgeDsiTKcf9OgX/dZJKNf5wtQ1vtS3PIjzrbGmjFJ6NzTicxPuRUNZrare9Wv1cdLBo//91Tt
DU7fLpYvtd9rNJ5Qc9xOucgWVl4zpb2rrjLtZgpkAcp4g627wAVYuWNvV1FQ3u1MOw1u7aAlOo4f
NTlLM8M62emuQ1+3+bx4wc+5lblH7+JdaToaLMuzEa4h2lAF9FJTw31KrdCnXHGRzPHeWAuXH4It
7WB/ljkuSDa3b30lQAodmC+ogBdcgzporIok26gSB5OO45SkmTtIRTq3wa1XmZ0LLsFtzIw2u2y5
CM0Dl2gpiJJN6AJinrL4nzGHe8m8vVKeNxiXdxdyS4U405YKC8nl0I//POMfxKpGu72KZuintV55
rPdNXOn3rL+qdHBnoQ0cL5RiS6y0+irQjr3dZAjyNctcF1642pldE2db1YJ9RrnNPOa/GwSxw9H0
M5JCWQvLt2K7Lxkuq6L9JTZJVpjp+4BnbQCrwRas1cJSJFI+0r4KAwhirneXtGbvpBdPEyXEFAzd
nksJxm2dC2TyZYtlo7TniPwIbq0xu3DgVZOxq3pPEJz9vr8PDadQNIddjTUUtu1CWrO5hluCZ40K
wAaxwddPKGiXR8lX7p3p8oCpBnao7gBxpJHr7j03px/6t+mIIxOWsRBFg2GICoVwjGs+pIlhVMu9
bWxzdBhP8+h8CfmaY86/zPyznDrsgsiFnenaIyQYj5WyqP0QLYirmwme9JPr8aeg1aw0AruxyID5
oL7AUG8Rf8azNbQyF4LcYnDqEVDFwNPj1ObY6K5Q1L5HrzQbP+I0YnafxMzrUB3q197vgRzy+uep
V+V95t6t505+agTtboDGpPhJTDKVWuWiI8YiMO6NxBKXSSVUs+UWL9KjGRdC+Fiw4EfC/PpVaJd6
UvuHEo7ItqsoZRmzeXTUzlNzcA0eCx0lepNSEXxGGmdTCelKcHBdqlouyux5Y80Ev5JwX6MFDYIK
AdOlbckqJO7PG/KaHI8Sc86uQYJgYE5zWkH7CELK9X2S1SxRKI0YsBmVN2LFaAvkGPgjWe6eqG9S
3/LKIpkRWlEJ+9Mphc7WNnT9YCziUuu96GTYVxNDlHt4M7rapTl27QF9Tg219HtCtqhH+rBNpk+2
kb8EqIYwviHMDAQ3yDZgcdiN/EMl5cxXiAvARb3iURWRMA9XqUlueDVz95z2r2odLd87SrIMXywX
kmMRzGlOuQ6KZSuaJEvCxoRgvA8lC+MKa/YWANeAICu0VP7C47IVPqJEE+M/ksoSg6KliFmBsF1R
T2H7EGJsoIBX0ob69JsRgjhNK57xBqqZ6uJEgm1ltWNgiIK7pOaVXA+LDj3BGcCPKRE0q4GFBL8t
Iz4dwst1MN/tYgZt+2Yn2RFlxBg86Kz72z+JhfhlObvnUYD+ZJ49Vp60hFSjwXSRY+whGLWjItie
E+O6MNMKsrybZG/HI7YHVFNpXdOe9V05OUWRJ+ZeZQJYq7XHGzBaLwSfHVKh8Du2vDSVXGTZR86o
7eeIENdbnlFYUFEQg5gMN+LWAPBwbX65lo8X0G4hk1vr6RLoVCxsq7JCLQClgsIVweBKoOHkzqRR
ua+acYO50TjN4AXw310Ux2RtJwOkI0n8S8/xPF5dcWE1MB+TMg0t5X2xQXSW7OB9VSxtfZAkTAYS
G3DzL2/wKPuuWBCl0mZe+odLptGmTzer2n2QZzq0Vu41wiCGBMODredjF4phq3ax8pFwrHeRKUIo
mtliAHlRWC49pjn2VZTy1SUVfvO7GOY5cZwqZ+XeFsZpnnjbNch0xLcWjbXekMErokgAbPTB9HjH
S9aOeaD+uhNwM1nP0/0iauf6SxbeNDaMljaAOptmRwse1nryvfSXPMpgcsieSGScbXfkttllw6Q/
eGr3FMLufKxgf2LyNXtAK0/Zkx1hFLEvsaIfYuEGV7NRR6w2V64usb7kz9nwmFwceE1D8jCvwN23
NZK0oqSzD/HzaZB+D8dZsD4wehZmF78ijosdAftM5FJvfU8urASmPsJP9FF4pI213jSoDEvcGew6
9DoS2nxfs3Rqfr7wQQf+aYGmGSyATVpwRUzCcnImMABJG7fBOZ2xqwYSz1daaPkTUPkZu0XKV9mR
QV/zA9jn/blN7EqMCEq77f33gEMBbpd1nQlICZXBqbAVQ+SBVK6rFFJ0ZX5npioh5YIIqL0EftQ7
1KCPvpBhW2LsLwke4tMPuR+hGCPtWx4lMv5jFype1qheLSU81z2+2v0Gz5TC8PQMBMFRRp9tUodP
LQDBjzjI15ZW10gerSDEu1R7rkF4rLMrrM1bD5yKqtmlL9jvEBlYhcM5Pu1AQr8e+/5QuZqyCDeC
OsVxbMVjmyMAzjprNeSio09Tt/kWJK6GeyFgzlVGgF4oQWdu3ybgwqLId0Gddmj3r0lMCejCtrer
aX+LkO93BXBlYqV1SAjnpJFIZgIgOo78rMl8ww2hUMTALzplAqjKdYYbqK/qhP45KeZh6iXEKE+B
cbPhd0Y30xJM+nhIo4TcQnCk/6LEK3VPVOSOwZOQ5Kak+2EVmiCW+AO1R8M08iPXi3cn2RyBL/xw
2taHOkzA4sAlke3QHW3EtVeO5spxSZRSEpQxtlZYjQFDTjqmorXBngzKW4Aw5qHOj9FsN3S3vxwj
XOTIfNuEzJcmTFi/CAGuEMO5GRLlFkxqlWIkis42VUhqVxw+jJwGh7UH2dmeVCORKf/N2i6Ig+EH
Q5Wsl2XdRy6b5ClKSegt/4z6Mcw6XJYs7BLyoU8Fg1KoTDeCfr2fLtTRCmQmSqBtGEcKjwIvZ579
RRwGSHa+wZZ49+pv0n45qegWcc2fArWxyymR2bL+7XG6i9jp7CnxWwFCxh3LHoSlp+4pCP2Pfjaw
u9QHB4T8xyuUC627RIphc8n/lMVYuBv7054SMUNRfh27W4/OLkC4wPIGnMu3/cDuM2c9Eyg/cjtd
GcTwMhEXCSH78bCOW2BWRxtPCouOPUDiC2T0qRTOwoUKCp7d50SueADa6q7K2WO9DyT2L9CSU3PM
XXkMyiQd8p1jDA4XDlweeYk7eC4/OmcRg52Ei5s1Q2GmqnBHJN1m9v5Urp1x8i815JUoc7YnwvJ8
9QPsIM4Z5bxjaXa/9w1eLpJuyS4WT9RFErrmGA7vMwF67kVuzLoA4lngI1tftemxaYbMOT8IRy1A
v1RUK9NZevHb91HOXNu09nnJFXUjyXhN+12mqxA3nHiVtrdOMmq4YiaWziSz96X4Haa1/TTQMQip
5uNNeuu8CuiPN8Cz63+3JN/Ii0Vuc9rNAFpm7j78QRwE68klcM1fMXCpKZ+oYtkgEVZ14h2Vw1wp
GtUcyVX6Iu0GtRacOWKHr90xIme6NZ3S3XPObPNSVm3bBQXzLK4o8VPYKNOUv6jdmsuvwqXtMTku
GdbbDr4foJtQg8REVawf4YYMKSRXBthCiICjduibEFhWbqWWH7Fm0pJku/hkBunH19DqMjzj13vl
pJtw6iP+vqo/RWv48b39SgV/LWuc0xY1EjlFNKn9uJe8w8CrUJCn056EeRc8Jkth8r05qtO2o9Qr
PLGYuREnu7mdBG89OOcYSLN9zdLBk3WHhDuqAshSDjTc3RhDOdmjzP+3BDafofQeuXTCZthBVNm1
DfeqU/HAus3RpHqnHmTOTKKpl0CVyxK/NIh1u7NhueguLJSNTgXn5qPrTEbkSKek2ekAPL0HpDsR
XZc3EpjPVaLU4I1AAXbUnF2UXiHrmIBYr+Y6tQLF++PueoGIzNSNJYPkAA33TAHIuvA7CrFdsCEo
lGAHKBD+gNxgaH99PbT3f1cDLcfOUdOPoh047CkdEe5feg70DxXZAY/zLRXtJUy4TS3PcoxGyuIN
8yU4dUtae/HH73thzOMsVNi5y++Tewyq12e5Vr4HH4/MqeSqmpezEA3JXsvc2i884wWsnrkc1nEq
1VR9Zqn3geeYiBJcLb2oGSdXd+DLsIMaNqaBwOHcCFphMGGAjDafiM/ZhZ040JlXEBjHfWm5WJ3l
dfb3ekVftpJZoINWJ86kUsSsnM5tXGOj6b/pXox9RwIX3znrBEvm1fGVXgRLezEM9zS3BSn6y1EA
r8qCg8gwT+0Kwh2yi4f54ueErBbrpfKXkOg7O47XvRpTEweU8T0mkmAeEDLzQO5+scJ25K2/fwa9
/Ki5HgeJ1jbCuR9lV6gxFEnF+8b4NtPQpw4N8EF8LUc1oCBHjfX52Yyqd0t4VnJKotHL1FOLAxOv
5CiB/es5dP4I1VZ58tGPnjb+RAs2lFj0Stknm0VHppbsYzoFtVuPSWUjfZWTwsx4WXlWOmnjtwlm
ZQDj3JoeFBGwiq+IEwA8a1Eyf9BknAJqcPLF8WeCbDU2x8+lsTl1WMhV4YQX3C+utsSX2GJ2v4Me
xhIkmKPD4CMlB0a88AKcpjjgCu1vts2oaRWOTs8/FYcSFP7Prqr+auunZWHVY/F9zwseRvxsKuJ5
lGl1gRzJfJnot2QUidJC6G3TJ/nKQrcSVMP9+ve0YLFsCJG/KWO7AMo5R9BXTtp7BrvJi4WsKDqY
auR5X7Mi4sWBcLDwauleBhrRtNsIPIucrxD797w0Bflys0ozgCgjLz2O6JEMUZjHTd9nYKe+qQ9Z
hLTRX+iVMbVnuLh/eMf6HxFBlkVgaWB662hpszjh0lwtIHrXdZ1FfiBbe1dGGNKbEN7+C9Ctl6s+
m5EBEN4YKYxrOYAlQIpyYhWKBxSrldgM/sWnbdbUOTU0XXRpIUEEOL/vV3o4aE1WczyO6FwnH0fJ
EOnO5deLlc2kJQylYuJm8ScoVCrmjuYR9B7fZ7UozuKmQimX73PJPZ6qnuN9uPYFMgvrM4cYJyaJ
IRG9piCHuXum22WZBeF+T8dcit2p7GW4fatuoZw2STETNP7GhpsPpQV8aTJ7bnF1qOR/nndibxpf
BiBzj8NNM5OOlVmRRgsvDm+5fopY7gwRO1aelxkXfuuGnJZxvnVTbTdlnVYbBUSnMlMmI+fxtHqh
w9BrJGkNxJW/NGUHFgt00uJ+oYNoiwe2HAqgDYqWiyxNPk6DA7AKsLjhZfb6s+bfD/zHXGeybAFi
/ytqiQbTjUwSMqas10Kaxd9n9w5e/IjG94vsu2isEwxp4jFe5ci6Cys43a2mAZiK7g3lryPdcg7F
zg1hlEUAnorY6J+0QEWuzCS/aNJaFkdSdou36VexDi6/naLD4gQnMxXTl4rUhd2tycdwVbkA6gY/
FwplCeB2aVmxbT6FlEjbGN981dXv7P5Ueczg//0wtFvSUV/Rz6ebQFrwN5RQWu2Fgnp71p+al/1X
PjNgFlwy/UOluOxUyddaKebV9K1Jd00DiYZ+rTAgEX2wdrKCAvEhbZBdLFFnBOP0QPbzlnNqgLQA
y8uSxNQgLNUH/Fc061GoU0FZ19g2O1l8uMVpXetbtz16Cfd4ayQGOOHZBaYU5Erf9pRx2mjR1byD
WtmbTtofhdjLLAbJZmQBY+08/627pKwYwMZ6Rlv8edSnbUb+ZhIYU1SnDpN7k3uxShNdivfp6oKT
4dhGJYyMMpjSc72sSQ25XS7M4JGMEvUWbWPiaFrEvI5QAqoyfDVH/WI8JdxpMZyTxekOqzQxXuBA
FCIKe+o60pP5CL68DOYJfC8sdD/UgB2I06nl6n/m2QVuP/Te+/06clYMzKzkWcw53nC0WoqN9UX8
oUC+FyJ00DtU9npQDiSRhVbwDIBzDv8LUVNt72FBjxEBatQvH9+E5buWcNBMkncgbELNG+xY3Yr0
WQvFTI+Dk8rcfF+zCqlp4YkjFjidBCtcUesSgsaCwt4cQCeQEpO8CJb/u5AyIMEWbBnExN7+w3gb
xPttQ+pspQww8UQhGtpEY3uVraCnGMTNYopoaGGfxOw/LX6ycYMpvpit9jeUTQf0hZCALuahTHbK
7BbJxsBTMI9RvFFz9YIHzKwilkULIuXKHnl0bigd+TGN9kbDCnjCoOS4lk3T8CumD+OC4/WO3P4I
OgNZbkofpSZx+88xIx/D1c/pBJy8EKdXD5oliBTjJiimPLj/O7DLOVAjfJDm4/MuaeqeQXH3azEV
rE6R72/dTQga7/Vy5+c6velnQ91XEqgstXHxMxJ7vxEQW5EfM5svOtGQ1kgKYhXqj5PUR70w33Jj
hhhneEsNk8cJOZrSUCN4NmWTKvWHID7IV8WJYz0fjT2S2YACL4ZvN1tv4xh4fhGrTHuOGfCQWffP
SrG1FCCfpu7vCHtNuxAT2t00o715P4md8Y79yDke7hACDqsoFKZx1G8BI6Og1aSj4tQfJhvqwx2K
0t/LSkvQFT0xG7mnhzpHPpB8Gb7nR4LFJG2j7Op+D19ou8m/6JG3rN0a2rq5iwgZnCStAhdL5MDu
MwwF/FotKyk/cJXbnBdeSU3BuCEWol1hkpvhZCcgavHom7fnigYlA+s114ibwOQT5NJpXZeO9t89
BeLmabARhyiRbxxmmlf+PyWJ1QGW9r0HdOeuJ72LuCD3C3yTXycSWGvhcFZplmWBzKhccrvqDFmJ
+lJk/hZpxe6Op+MU+39bTR+E2gfg85G4MFDn/LgDBxft6bABa1GUrKCoY2jBqAmKOmL4bHRPj4yP
8NCBZYjE5Ugu9rgIyWHVuUZL9PUNpxLN570WxmePtQC/vuqs7zpSUtSTpUWoL/noC1KpTPMEbaXU
xCWAS6vfjCjlMoutt7XaJ86MHBkud4+lba0bmqeuuxplVtKvreqknoszAOtxZ5LBz0F2sjYoWJTP
yUTqcF383OmA7v9zWGzNl1Bt2X+qns5H69UECxqo9kTWVGr3ZpcqoLVQmZBtxPeAxjRDgzStn3Vp
4p6tIn/g2dUX7lEBIGZDz+kLaAJtIBFX6bK+WTgvx5M9476rj4+BKxlnUZmt5EeiIWQFx5n66Y11
kTV6EPKKETceSfLmSBS4G9tnWQCvNCGbDW1sXBevG4e9KlXAC0fB9VvY3NnBBumk3V6X5HKc04tJ
ZeMkA4LxwSFAti0ZurSDcuql0b88saWE3kug0ZlmfBdtOkSYOlgvMewWeImVkRl7PhT4igCs7DIR
OGlGKYquvBVqTxox39Kage+Pddc/JXLreb6P3vBre+H7NBDYQ+wVSG7ks1XoK/Q9Ctkl8lWWrUSy
4AzeL3HwChloDDFbyAj55U+Zxz0vKUbXI35xJ4u0BXrnfxxqpKQAEE4tcWHyFReAPjMW6PHk4Id+
fbvCfim5D4zz7iwLG85xFhfGUMLddagvmx4/XvOiqRaKq5QuVz58OLRYU7okAfaQM1AcKAc2vPQp
QgM/em4eRNjaMGNq8Xito8cQ0mIrs3xmgmiBA6nP7gE0kWbPgGgSfCiGbeuc7PfFysQn303K2bq+
2F1k4bE3ja7vTDYkFCC169efz0gfGj5ZpqUF1MqG64f3RDVNS0+jur8TtxTQhUEKG6iQojWeTgJZ
aLGDt+8SgdZP8mCf1DqyrCNCC4hUwwjhu9o71SgFd6qtyEcoIDnRTODVZEXyGgHXzURyGIs92Lcu
oc9DpT4P4+2SG6XeElN3g3JsGn/dnSpyBbRqvPreMP4k95BrpqT7gtYS9cIR7EFD/F+P/H9231mJ
RTL7xnpM1sEeIBgC+vHZ2n5xWfQBsL6TcRARPbPpzwGMEwJR8aREvAo/thYPEKoik/zGQr37dFoA
SUY1ePH+9eshQbgIaQZHEP7AKjE0tPGd9Q0kz3YlWYSa0NRsMif6t2LlDqjP3lmrW89Wg6U5rJiB
vGt0drvhYDRCHQ8U8KuQcmeGOtGQDyX2i7/zAb6g/nZAj36y/8wbZmFFiK7im++jrPnIijl74bZ7
6UeL75UtU3P3Ca9OpjaKClzoB4Hp6D4o4YLpH437OZz57XxjPizc3LhDT6COQU/8qnq/D335BcC+
qUFJ8Mpju9z/FumjtriwrEVZgsIjvZxBo9Hw7zmbDw+JDpBnYnBp8ciOLMP3q47bcNR0MR/NV/td
DelNJv5o8mqsJPoubFb/QXehmYQMjgf3y1cno1MjrS8m+0f765CZbBMZltqQld7pt2zFWfDfxi67
RPqM93OgU7R3FUVQWTADQwdfEdiqKht5Qa6vXL+arbfM2KgCOK1tZiMs7vQRZoKaqXxLvfNFSeRW
QenraNmrkLyK3XvxC50Ow27A+IWG63o5yBKr8nD5sLfp2nwnelEJdli9QIGPznnn1HTI735cQAgt
qpXCttFzey1YYLIhjptGJKsrsYhmCxyFD45+JARQWySmcuDX7xQVlh0oucAsyugnToh6Gmpclqrk
pUw1guGW6MkofPU7U0HNdU9uXO0Qi8wq8nb2iA2h6qwnN3C52SvZivnzhstZhQSeU8OGZ+XQED6E
KxhoNoB8uWbtqTEI7eYgwrEIhHg3/hniq8WRBMZe1yjqGnIEFji5aD4UOix3MPgZlyCxBnpayFPQ
2vZ7QC5BvOJoc2CDdiWMpm1EcDlx6XNv/GY8vCrI3BykKev9f9X8HjiyOUEGh0u1LoQkpdMN11oi
ggsBEzNgOGd/Eup/LfTD2e+zo/WWjcHWI7lNR8y9l/K0DuhpVxmTEVZJ2UYFynLlrGgWXhSwWnBb
4svpBkNNon0xIeymJjTcTDk9ic98G62k+NF0LfD8fUJ+NURhLyX31uW1RGf9w2JuLZ1XwsCjQxl2
Xkkk686rU61LU1Nn2BBxB04imKXwZ4mMTZE46SNtA7JzMtSv4HALPItlOoTQQX7wOKb9Ld+iRgCR
tS7EJmiwZrTUwQ2ySbZ2/BCLmSLHhQOKKRPdrgYhW8U8/+0Kdcbn7SpXB9uOuB6LakCR/dVi/CwR
z9pdOwQzNHvA5hOY+/wFppK3uED+gc/2JBe8JWZKPyULYJe8fLwGQCQeC1HVHvWcSnaWtYgZTF8I
sIGlcORIBrX+d1ebP1WAbosy0XGM8aqNzHqqioUR4Eb375nsS3sEmmZKmIITTl5c/b1xXlofeU+K
V2rVdgB/a1oBxwx6790F18I6b2lwW2bYOQJ9I8BMnrUa4KVaGNwyHb2v4oouIoSh1HxTW5mRprrA
jW0cMOYWBe4Md9u8ifRCVpbIfM4AoUUS5XwkKOrNS64jH0gNo9HRH2pkuIq44d/n6t3wRJYsFSkx
bvwXINNJpqsxYjmEZflzrOo9SzoZGgmTi6Yxcp4GXOzAYSACo0RGcQuN4g+64uGIP4Qc7Z+TBk3K
BhWfKmEzwWWKwS9kTPKADK65j1hsl8NNqix9CkIyJwkPEl0nTgmFpnRgyXHdFmfBMZb5abQW3uFt
SPX97NQZXGS+bA1c1n9wP2rUUQ4aA1j4HWZI1RuB6zJWjd1U6cQomqF6TWIQ8+uTCJGMZsWXerUU
RPs7dfCL4zzerafX1wFVI91OwEDWjersj4sS0fjphI7f6+wheOnFcWDBVxhVRBYmqxqFVo3f0XFt
fKw+UgK7MVdXOI/p+CBXbhYVA9PemMFj+EustdZS+G923bgOZZ7hYiKt3FTlhjTYKuZ8UBMA1VrU
sHh+LdB7VpZaQSz4zPqW5U8keD+8Kh3afTaE8Z+RfrAUvUQ54/6nPLNN0dbQp5lCm05iOZ9xK01h
CtAAOnFkB+8OUNoRHErvzB8sFWBCsbbMSjHUOurC5U4rlk4ts/tT5w5UaSZnI00ijMC2VkHcKaxM
uejyUHIVecdoHSV1yOvx3cYvz3//BdjYUJ8dxQf2ep0yx48YnMwd6nrkQT3n1tCSDYJ0JGAQkw1S
eeDFHWJPYDqBaDZ/nSOStSEGZIijuNEM808tk6j90Ke4CIDtlKMIaUy1gHE1VXybucFe6xYrcUCg
s2TTNRyyblmnsA4TnCaeOzx44sXdXhNSW9Zym9/54vSriCh3yZh5/paMJI0ghF2H3vi9eBA6rEoM
cySqyF/4W/vpBxh0fz/EonjXqc3G/k8qBtvIsVlTZHeTRuRdil72nulkQqOzm0s+pWnIUXU+3i5/
fSAqVhg4/7QyKPjRnOHNsUn0OmR4eMc0E9D6o+zW2hzKJzWmksWx6uFKckQQkZ4/jinZFUR1tRkh
ViqxZbdO+nPtXoE/w71cj0fi9d4otYaZ9q5WJfFqkmYZSg+J4JiWOFT4g8pVYXZU6q/2aFpbIsDs
ct8h8MCbhx9UZcuSrxdaCQw2gANLvUjTe4HB74FX6G3yMdqnvUfE702QmEZhlnD576x3AXinlWw5
fmVHjBeP3Gjq3XZFxziiotExvdx5JL5JabSNmExdrldNTtAPG/luOhUc8UpP/oqLZE9TdPKIOKeg
1G3lLJG4/P8vqhZNUmDmRR1DnQT3Xdo7ziCqN80dGTWox7PN0Y6ZV22VlpzpJFqto+K45TZdzUn5
wdqBgPJ694iBj2nL67o723KeDj8SX1aRMLBvI+qAv5mu+q+OCnp7+qDC5P/hZibJTtPTRLcblJme
pqj7ealDXDuNNdF6A77lbcFoItcx3oGs+SJJn9/QHdOBEMd8wHqNdhbvBU4hof4T3Lr0mWPt7Iod
2od0eMRUMCZE4caLlK3xTUhIUifCR/PKuVWhv9fV0OTbrUtbHU0jIYxI/W/j5Xb+QRdyRYgp28rF
JyEJWFnQa6H8Cc/g/eEgNB5TAi0NM+0HlYxPvQxqhdq4YhtZYZKEbG7nD+AzdL7XZcxDLkLyrbs+
8z5akloPWklVAm/MnkPv3PrdUn/vBArZxWim/upymh6h1pKUQiTcv6Ta4wwCqHE+mkrDOgVGHo/5
kEYRIn4cB3KaQmgAhRhTO34EwR1NuWuK10e8Uvrx5YdmYFzD3vWq4lXmwQdqyGZ7wk7GeRf47He0
yJxmwXlpWQ7ioo6/qkFIift02k2thz9J+8o2paQiY8/ODS5C9cWCmEds+bafvYDAWlpXs6EWbHNa
myrbfHu09g3ch7FNwd4Y3tbFgcMpUsRB29eUpGBv/wuhxM6rrn//0mqYbG4U1gf9v2d+TmKpvE/m
iWO3h7WyvDUwjOIL873pV0hiSC5yMDt2pCRa0PX4uPyWzUw8s87FF8AD9wQSYICeYStYs37FG/ol
DIO/mRkTUKBnSLF1IRZy3J4xPNiQRGDSEH+JXM/BDCMlq5bwDHSy1aPErgrgZRSm4MGkAYALRtw7
DbTOwBW/ZccFCg8/HxZny80AtQY1m8KkOtXKzSEGB+aTJMp5xZY31VsZQHbRXfh8t3vIbIB5B2Ty
zc33QZKILftkyO2hL4bDoaygYtNK2ldgtRbjbmLtPg991JtDipfnBZKz4SImTW3rV92g0iZl3360
d6UuKx+YhkMg19pZXeVYijoOr69N/Rd1zG89hyZQFX7m/Zof6/S2Y226wsifHTBUH9DTypiNS/uO
+cr9l8hgDK8hu6gWHbtlzs/RSA0R1dBZLDyF0607au4TrqIZfZ8K9qESt9CSUrYn+d+k0fKi9MEl
v6Y1ZK9CucNZ64LhNigTPM3iOmj2lfz5fqagojpDWIuzViyuQDzngrMlahHRAEWMqk/TIVseQvJp
L/O/evicerNcxTXZ0Hhgt+sw95arYwjze3GQd717GlQsrFuC8+XhnKCxj2DhgGDbEW/YGFQy4jZh
dWFFG7vpmag+JpE3YAC7UYarOdV2misAp9k9Yw9PdKbddZfpZ9jm37odu6BaWwMWZWZ1lxpi7onH
yh+YpNWriaNd8jwtM+agFH1j78V7sUKdR6GDvXI8fKjNO/RwjBGAwbLko1UeF5EH+KpFA2lHIiiI
djxl+v8NAvh2C5K75aa9Pke2R/aKjnSgVnti8gZeJ4uJF4o/f1T7Lwe/MekVoiyCtvCSZkaQy1sF
KBO+P3vfmrTU4kzHPUtsvMDEzyPkXw353zM46NZ31th9gHjUfwdLvEz8svyt4SEfHRxj2YxeVrhl
3KsRvR1GPqifHokQN1bglKA4cVjQbzH0stwgGkgJhTKBQUEzf6+wc2exS75zyZiM530jq/hYBJfk
Q93X7zWNq9zgvofnPlQ4rNPgSQo5XIRXQCI9rQFRtHjssh6GyCZOys6dQOBKJucRB80FFbYsBj2V
wZefWUhY9XeOYcuTa1tIpjIePaGdVdZOMyKgB8YCw7KeuA7Eo0EVcrogfnBIkjYtMbzbV1tSvnp8
IVH1wFYon2u5hSN4RRLeXmtdYxFR+9V4NucYNrPEZwTcjILheGA+CKTHl4grPHGRubCSzqIlgeck
bUVCrbhYcueUEVjiNmhVtXjS1GWfybr8xk8NBT6XyKH2e1tRdBqZM4z+J/vBSOBcD0xxoO4KG/W4
b0sXKmiIkG7KYuRdc/aVMz5QfHnxjEalFA7rppaISoE0E1T+2iLQEoWwaLGr73B/ZisbOP4cs5sX
ExUx2r09X7JBpdUAKF5xMkkpp0yvxjBE6EnE4/CSlu2zrwRzzWmGTvf7C94uy8oqaSFlcsUwdXob
Bjxg6Tlvbth9utSHSOHciQci107UTfpLW4UEJdSgzkItfOKEcGirCSs5NhKpI7a4o7Lg0MjRAEMA
Agud+VNhlX4n9+1lHvfGXGzeabm2XGFNr3jO2ZDHoRzNs9rzPYhuhXVdn0tcsUhZXy1e3FjoxmqE
CR8McOp0fEiTxNjZN9+ei5J5dqDlMREWG0VNvDD7psu1/0ldpOofQqgu6weGU+05m3EyAtr5h5PX
okA1sL/s1LHT65LAf3MNqzkEO9cZta6al6rby4BR9QKlYHouSCXId5+F38sf3zFNCRlov+09uk76
yhevdGa7iFudKYeqai72diiqD001tPZMMbAMuQxvJEK1iB5AJVBdHsnpSVmSqEYrEcPBubNWm8qE
itBwG0V1sZcgOmnzkcLFMNxdgDpY5z6FplbF+z1UvyFm+iNmvmrJzcwchSWD9pezPeRxn5XphBei
IzhYmb6Sw8haWeSJmNQvPSMP//5r1L3eb/mxK1FFKoYv7PHcgWni3SQvxXmrpIUsHO91syqofJvT
+zJhC0mj5ijAgsQyT07DS+e8PnwxfA7yRxWUQ7ZMqZLC7NZ86Cd0bEE2XxbufEAgQxIO/AB+qQdb
w2KoadbNOuJs9h5XR5ER6YwukSJsuj2e/cgxIugQTF/KTv1Y73GjvkeYJJekrwiPBzuR1TDGgr7y
AjGVBNFxzUPTRdGyjey+rx6G/zcWv5oI6j4tNs+QsB0VJEd56NCfIJ7xjC9FC3SISGWHyJ8gSOUY
lFEc54AKxdNfjliUqL2cT5/+ZWaOGY+YDCjHDMxdYLXxOyS3tUPFK8rk+MTJ47cT6OtdV5juNoSs
BNUEif5zKF5ee/jZ5VGQtw/uIy3Xk7qJfYS/7c6qZHmjz+RXkTlSz3iaAE6xQmdj/GYrIKtKZymE
/7Verl4YXZZybv6QXzl3FAZDgJDM3dFUU+15dJ7TFDLqRV4yKsCnzWZKIqGkQfzdtj/5dae4rKuZ
YDpgCGoc9fiFaOCAc0A3fUiV8lpIulovEHUiDsg236xFdIcdgJ1qqfNdnhJHmQXFRnaJN+K32lvl
SgGnmdfsfgYgi2clwlaROy3hjfYi2BW3hcg0HaYKJPFuOyiz8cSSa7ltA8o9EU3YIlpksC+RlIx5
lebG/afAAM4ZzkftpQoXl4b6zCHf08ATvexJ5qasU/gnSt2DeeME4c6fQnEMsB88gV2gv4EAlIge
F7Qqx3jD9hUWv5vn3DsdOpUzD8nsIdmfLQ4xoIG9s47ATvYnKjr4mcQp5U3sySb8nfy8oZ+eQuau
ofcogs69nrzWeD4gTX3m/PRQJmmmF+K0ZmrLH2o4QkY1iR5mbFYb4ja5PfSWSSLxSh0JRF+ANjEq
22E5qNd5XUGQcrSQXeCHtWV0Gd4AkUL0zVrzfLrBN/TbCOWp1HJ0B9PAeMKWUQwxy1sBCrP9DCCM
8BpYiPs5NIujzA+gRnmEgJ0q7lrx38Aq0T7eHe/SQOQIbh/7DZpiH4zCFo6HMax3YdR5vTc/tww4
9umSt+S4BceGqOP0YZW5c8TDWDsZahfSkEq210YQkhsIa+OsZwf0YFeKn1BJ19xEdIL9BoP5IGlC
NQaryBzLklEKaw1VA/6s4qu84mtL69Eqh2vGVk+u7u5xNJ7psgdhKcfx9/pIjyjzCY9kmdqSU0mg
AlPHPbtlCnrZ2/pjkfLtfiTNFptTqdMZb4yXPcM5Qgj/VSlBLMkJjr0AwwQtQfsPsJtAKyYt2M9t
PI9uqrIL2aSh/VJrfX3FK89h/299l4doPH5GaEA3wFmRfbIlKnRzQR1y5tp4RDrsvmJS+WL+cq62
9eWZhTu+v822UBWWr1uhBW5lS0LU2w42a+hBEcvATn8FLQpwdsiNfCxZ5dIm7czZihy2VpajIchG
fNcZRdXUVbluOSNjsiFjO0Br90KRFqlQAh39+Li7yaQCg/RZhZhuXO6w1kqn8/Cgv4M/S8zrTUbF
uNN3EQ/V/j7RIpRvEqjpQahRT6wMPC59v4p8i3Ka/PAI50BztSF5M+HS/ScnfDMNRedfVE24EDzb
Rvp9PPOnPx2cpCbzXjP8ZJj0CdOjaeIFdRA+PP7zaayCHrH3iUDL1sqHDDBXO9NKfveIBH5Sqhnj
fW1tDD6eFVHfk4IPQOeoQwANoZYgKzNOdg1orLYW/ZlCreh25wpZmR5wsbebHLGpgxF4iYTZRbBE
TUjhA2Uq1nEsSLvtavlzi9A01nT2WFzzxnxsgX5Wn5QTmU/lmGxPgHr0PUicXHC3Jr/gxJoqklcY
D4ktVw6/k0ZpCdD9C/9XLgaakpxKWqZj3mcwkMJ6XjkIk85Qrv/vQL7dt5QQXmPuXZ46+PV/K3En
B1uSb+TYmBIDEm28XMPozXviFn/L0DzXL9jz25rTgxiY03fGBpOG9HMD0Fcdu0qxUqsjp7og9vuN
3uA2HNUwKmeIaVh9Zp1GADky3bhzm0b9sfUnXhsUOsoXE9TuoIQHBlHgzUvpGHD/YG/1nAiDhC8n
PnN1MaGjhKkUw/G4+ZvKh0/Yq1JMG4SW77toltf4cMyJeJ71AKW0euf2BdGtoKAjM3zyng0kw8AD
EW9SXI9VY+DtB+PNvjj0wodSinn7mI7it5aGsG0JM4GFt/aAQ0/P+Ow5CHPgTqyFF1zysLG0Tnnj
tkbEW9/NG7nLLlylrjhvzIGPz2HNoiRlfcp4zmwYPqPEE5nqgQGAc3ap2IzlCVsfGnXgJonF17w9
CqzZufV1VWW2kKQHmmI8IjXKBU4Yf+1OcIDvLMsdRRHKlVQ1YA4jyfh9oRzXDF5oz0WeFHAu64LI
4UMuhv/Rz9Kev3sXLDHfOqJjxsIR1MjehWs2k3JFV79NHL0NYwLL2QwtRi6Kgu4icV+J2Xhi5rw0
3gzlXPT2mAjR9IYr2/CZroP17VSqC2+qy0kOQkxHpy4pwhNlTNdwf7BcFZ+ve8kDjc9iuQosZvA4
5thzbXI5LFU3NMvA0x0val42YUUVpIwyD/+wDSF18i4WqocxoVRSznNmAfB3iN0I3brLcjVW+Mhu
fDP2s9IVyYkybGWFhPmIqba+sK4X72YMAhwt6ehPQafk59fVesBhzaFaY6cw7yPBDnQ8i5hLUs7Y
DCrmUORryCfj6BVLVzPr+vdon311mfdJm1Qd2Mx9V46o9Tn9oSZTM7Pxy3xTzFzpodAGZPjqTanA
RLKJCwKVCSpjkHdSv9ZLA8K0cPg4LUxhovyONYx/tzzgPEitUJx2bz+uegp9+ThkPX5LYhWphVLJ
sEoXBe9m28hY5qHyt5wk9L7qMnh5PhET+pdT/2MDoqccTT+DKmD1jmkxGhNEXCpE1rSootsckqzh
YkErZC9DTA7+MZU/0b3QfjOyDPdVYUMswE0CHcOE2yIfyLvQirxULYtM7Cy9qHUHO0pTDE4fNvmJ
6oAgUtlKIGTgOe1R9j7yEKxhbZLY2X44ZfM4ur7l4h1qAiMzNSWCy0OF1iSlgVFwS36SFleOXgLm
6Mo67Ar/x3De2lYdKigDKWQCggEipcWjPHi8jNajEDGIxL0zP1SPF2A+etd+a4BFA+IG+DqhzGpl
aVKFyefNbrK3ilB7p+YIHX4Ob1ieRCM0T8nICdwl2NX4asuMrJWnkTnLPsojBj0GGF80kdA3fvFk
VDeEzpISkC8qCH7t0U9VO1tmD7GopvyFdNTEEip4atk/WJtpULj6vDmb00p7K5vENLOl4jDQAijP
CRGjQdCB5bUGz2CAFPAXgsSCRPXZ/gLOQ5h3SsU27ZrTTptOWtcDDIRcwoslfrturk61E830txdt
fu9mdu33sDykco7nPdbNLYyRgAV+9tovg1TqGjv4xHgL+p8PHpZSj7tT3mryCSZcf3RoQg+Cy9Ql
bFWb7uCScx5NqAvoavdQ3a7RAIbEMmAf/g/c2fbhdke0RN+q5yrNYC7vARJBQi66X3MC5OwMAEtJ
defvBSloeL614RzGL6jGvB6axDcxAw1rV8ltkSQDlQtm6XQSIpMhCpwJ/GMtB/1BdE6YiWaikh4w
VB71ArtAb2HmTr3Tr7U/7y6wnLy/Jn/S+o9a4k2xbaRVbCeFMHfwdDunZwomKnuPyvtyzVTLPeRc
ky2tyGRTCExr2lDLHHBfSf6pGr4vhHSKZsK/WsqO4wmycjbFWoGixXJFzLlxkpTvXcBIW86BMQZ2
Ue62vzZqrWWFciygu6xuL7w6arzGh2/6ex8UBt//yd4HYa4kzlnjYmDlAzpMec3OD4cRCAJiFX+X
Y6juuBXt7knRxQ49dZLCyjuaJsde5UwyD940lyeyy0T3s5UDk/IPWRfcKGYnD2uyqHkICDwDacxO
vait80vsuGyNzvw2nchMEZbljIVmzoow1leo45I3XzlQqJfStAI+0ZdQQeCxvwHbpFw1nxiJTrYC
KaiDBKqQadKP93Z8QjSHR3mvhFUjOFwP0casHZrw+azgSqdtKIzV74DLXbgp7MNLgO1LmaU+OFac
u3XOBZUhmY9MUzTA0s4mtxHZNECO3mY87ylKvMRP23weQq9MnSyNAIuEioBD0opIeJIeJGeoxZul
brEOXKMBt/GTYwsuNkDZEY1MQJGeF0wdo7UJ/+m7JKPDz0MypOV+66vKnSdWK6q2bElDnTEPM0/t
Plf4mm0yilV/LKvE/NNPTH+Pr5kcdqTX2NFXtJode4SFa9CD0++Y7866X9AkxUZPBM/20UkIHyYd
RMPgC5lB5NvUsxUZwzmQ26YUqu2/NVG+OG0QCsZPeVCUDpZhxgZnKMGNFGMzcae7+kqjduy42/JE
SSnAeLg5P8CL4LqgHIksijEfWatGUdJii+Sr8x+S31ZN0uLTq2NCbaAjnj4j9ULYAOdQ/FtQEXh+
oQI3neoNIs0rc7xGZ2m8npKJjF3Uuo3eRLaIeVamBt/5RK7RBCQEXGHyyjC32of4zR87bKbwk8+s
2Z/NV2ZLn4W3dMHmydD46eoZkjrKGGjYrESaqO8JZYqu9wsTZrVNBUqJ+hmWXjfRS2Uq3E87qBSQ
48EHzKX66VsjpSQDKIBSvNEIjP0vp6oyrDV5LUtJBj25mJ9yjqe2lKZ8rGQd4FN9cdrecZFbYAQS
7WWJg8UV5lNId3ZR+tBjxBMtepXr/Eh3HLqo4YxiKlTIPbW+HJ9x0hTXKK7szHRR+JTJHnoTDv8C
K+XJ0NUvAFmlLeyLlAuJkC4aZsIRt8MOcTfGOMTjsUKx0wnJPB2autzwFn0EXvvPTZP4bCKPMSWq
wJp785nt+4cs2apydS07+CkfZjohg3ZZ+vYV+hfxn4ABjjzxW/fr+zRcKGSDymcrHMQlsLST/Q/c
axKciqohmF88mahjwcZeX/SEFS/czdozSAwMPxs0jK7JN2qmTmQiQIYdfjZuUiN7SV/XtU8GyOEv
EeudJBnxdxGLhtbRGfcXRt+MOuk3I9yFBUQCX1l72E1S5cXnN9+ApV7udq0/rUOfnEvVguSSS3mi
UiRLgso+kBcNJCl96YQOQ+smshVycGiLm6XEDQjZy7Jw3AMNk94aKAoohCG0o5oPM1a/C7Zf7oaj
LWzze2jnLSCIcTuchGGtczJAihXziJ7AMCmmR1NlUTdozsBtGTmKTc09eKCWflNo7akbwSbUDihs
7sPR/ZXwo9xlKEDa7eS7W8tenJPgrwORnE8m+xN4WcGviZ8D4C6nt3VYDp7NAhycZEkk4feb2Y0g
gbrwMnSHmDBqhXezup7rQM37aV2U73mfbWSxBriE3qwVnAJnwD0fL5E9o9xxIjdpNTmMRXBLdGqK
dWuGy4EQx0Kt+s1HL+ZliM144wWw/vKrvjwMdgeuDO7M7sSgRlEwqiEbCfQtipDL5+/tiGZ/44uX
/+YUl48XEoWBeP+JwXkNPdtzUPPX3poJQnI4U4Mg1RqOnp4MGhg9XjOL7aH6QGcFdUKOl2hXjfiR
Fw20tFDQTPf0mzGoRcsWNjOeqx3gYrRoNjfjyyeRrh4RIly82h1ptZIQNlHqbLH3kSAH4QkB300s
mNh7BDy0TAiLqvLKbfaAo+nbvSg7Yt4csanS5or7IgZq3ENBFnyOAnYnaKO1gVPb+y023cRJh1Ka
ZMABkb4B9s1H+8Kcl+L5RGKpGQdUhQPssxSZxF//bUeZFwCkWg6U8l6EGA8udkJB8HRmb1646aZn
bFfqK/Esoj6/wyGYxD4KO92gg2HMzxZ29SN/anEnSIiyWCjx0dibcD9oWtn1aq8yRQaxdz6YIIAN
n5OU11cWGFvQs8DZbuRPV3Iv5WgeLubpocucwrN9zDjQ9n7T/IDXb4xmaCCATNNcae0uHip8OtVD
naIPY8gUu5ajh0HZySAsF5H4Y9y0vN5Zr07MRu9M3qi5lRRpxT6ZIihnwW1aQMnA5ZfyJQTSXMo9
cccW6SUBDeJP8lpgdmgoJ4EeLjYiF1ayOsrTVzf4mODDFIcgLFNKwr85Sn6Djxe2vEjy8n85WGQN
ycUoNzAn2ZEzp++eMTdMtE/6gdtqE19gTq+HQi6DZyatnjvSgPGkKV0kDOgMwya26Tyskvu3BWvo
byXXCgu6lQ8J8ovMZjpx02x4fmOVafSMOijudFoPICgBdPWG5w12LbDWD32qy+8dP6Da2g4EDdiD
0uzbQVvio/COErCSbfw+eJLz/U/wnlkLhR9YZQyKGSu3g7YY8uw6UBZlrJJhXRv97nBkjMaAWOFk
KkR8pZ7oJyPymKJYsakt5h2AwkNTw2AFqlgMs/lML8pdLO97FfpO5OhIt0zF8jGe9SNoXUXrFXOP
GaX5wNvnxnt22snEX+HVhOb61iDiPRMFXVvug9wsnYaqD2eJ3r6dHsfdmFfbifAN/sK4e2KeRycf
jvGyX49Kbvz2WcHtxG9yy587x1qp1GhhX6qUjHI0eS5Hwme3n4Y6OLF0dombf/EB/zhwrlR8dxwQ
sBbFmZWmgPkyt/H9Aop8KfopTrne5mhvGFOFqxJH5zfIjC8wuNFY9RJDVMVFEvy53hshUz7msuO2
Iju5G3zY7chyHVsKXyZN19sff/Llsd9iF6+g2pVpzu0SCSzDhvbxjljx2/1pwKtmpDNitObaPv7u
xnPXNDn+nMN93aiAcCy5EZLBRdTCfEkTt3KwMNTJJdgBU/e+IPExIg8nzIlrPOMLX51qgPwWvLLE
K2NsIShfJahDSH163yAS5xltsnQAb/YiZTEpsByEKfQZc5vovHw3OgZbzn3fAFFLWaR/rv1If2C6
3RFpFnS6yldnQcap4Rsb83ApL2jklaPCs4gl0qmdJGWWEmvToWvaGVzsYwCpts0c1/3Q2lYzWgq5
hyY8fFFsE+d0HfGSiTXUvJpxHFYZxZcFfAzRT23nI538YbjFeQYGbhibx8TUoplZzqOFn5/s66+y
jr4eqJ+Bj7GkrKN1ZjYfG9gqH9LfxCoFr1h+QQ68khfXC9ODdC62I4jUQ1cHTkCCCNuJL6ap0Nab
OhyX8Tu0k6mWm7kKn6t7CyY4NIkhadE2YERUWqYEsaWIh+xn308Cfo2+a3/YsnIVx16G7Zqt5Pcs
QTLwUH/m4JYjrTcKmhKnMxNpc5HmixO4A1zbG5o3qvv4rh2m1GgZVfZtvmucOjoc2oRSUo4Ysle7
4l/kAWVVj4aQecTiRgASAJGaFBgfmnf12fSzZhiOOsTBtnV646nST5UjN+XEDjJg4SbgGQltHoJn
iHrgAzfqGzj7TnikNpRRU8YmnpjcWCGWaYzffr2CslSe0zwCEBJspUy9dXZ0YfCU4eBkXi1lheDv
P1DUEJBKWqDQCUh+8AEtjRDE/9weR5VqRyjyjs5A6Foe1U3LE1Frkqkd26tRBBdCpJ9O0js8H+b5
YORBjM/7Cf10t7s+5atUTOH3AJ4KxzmMdbsiF5x6oduGSKPwONT+Z61nsW5BV3ao9ljD4pvPilsO
tffrXKIxsb0Mj620CVNSoMhDwUyOrR5AFFAuYhY6N0LR28f1kykpP6+Ti30V3GqEaswVEsTHVj52
hYJ9/uXzwGMFR/wkfI9ZR0eYw86GPJyK6o5y7mA5qIW9Yoi0LFi4nFBxi8cDvGd3Dj/GX8OOO5Gd
Ia3rlueAv/DV6CcLP39ApJZB3pvglXMziWZ8kNHhDrAzwGOnhfS0QB/fmJwsHDkAJZSMN6YrL3dG
2v37cOL+7pdW6J8L8Nw7isr/Bds3Y9n3s35kjM6nWSMAXEBDsMtyiaTBKRCWqs6HL78ShqAPZoJr
OZiidH3dovqZKAz7fFG7PM+J0nK2xvVXr3y3p4YyqLn9FV6KMpF8QNliBVHw3N751VMSfawEyuUt
8D+wkGx0hugxLVbLvvPZ8ESMg25NoJdre4O4FJwIEAjm8CjoL0+/otaCxErszx4XBo3NL1CiT0bv
pIAPxAp+W1JtAPPRtY9ssYPyCd1/SWacGHjOI+5e4qcUrDdIvsTAzLQXLND24604BOWcLx/fU+zw
fNjntF5cX2g5gBAfIAncutFFcF5bRG1eSplkAx7mSai2PoAEzS/4fpdyI4+aUvqYb+nKgRHhEQq1
0NYDiMisktf5o12LpchFXOuDkaJXaIzBZE/2epBlAGcZZYJsCnKs2140BNj6ot0MzzP74b342MGI
68KWqzMAlESTr1tj49ieIgdN3n/dcPcn14rJDjnZGhzOFbGuM0s2e4UaT8G5V/MfnHK3T0xPJFio
/QjTcgUkNabOWpXEC7mNL4EkH2UfL1tP6eg05Y/YxXf7YzmzQAGLQAYzlbMOeREJQdL1JWXQIn0k
0AQUnZh/h1HTKE8PJ5EuPkmK3jC6ITqc3Lp0KpQZCxfzuvNMh+pl3afIOssk/NnWJWyt9eadRt9K
Nf33Z0XLwzbNK9/a0mQVNo/f8G7Gg08czgieqLpDefyz08y0dN9TFdgfqH8doO9gXe2pj4lM/N/X
SW4CRC6Hb8utvJXNzmNUtzXD+sWLx56zykATyt8Hqkdkz56icw5yGU7nnQ6NbEFIesn5Gipx2TUY
ItA04ZCwVywp0H1/c4TwLsKg2WXEKZYIXMs7o5KMjBq+BMhs/gSaMuiacTKk0Augprj7rG9yZNFZ
3L7LnvZwm5ReUn6eM4Ci7IaQ8LysuI72iMsCsA7yZ311BFAsSZC2hnrjMeY6TqsE8MqV1JXrP8bC
gc7EF27g4ttProiuoa3PAa0I7ZF+IJ1Iykc7lNoOICSYCPmTU+pgUKeCQgILSQYd+4fdLpatY0ww
yJv77Od35oexijbyoda2lFSYu5LF/6KZDakhkSSP1kMXwRpMHYy+TseUNJU8puUj3PtJ3wA0Sk98
3QYJfbdG3Pll1Jv3j+7bK/TQVDbQUD6jDf3CfgoDe1jwfv1t8jNVNjCZRk4KtNSmZynuiSbWZihg
8ordFnVrwUR0XYmToSdJtL17cLPhSyk6X8OjWWdjXyfw1o1p1QzK1332ALO0Gxlt3o4WAFKgwvC8
BmnAh+yDTJlRN1Idf6HTk1pb5oApz15IMx9d+SwaPgl0AMcPp9PnO6uAC+cVWIGlBFXM+KZQK0Ty
JNTHJ7/M1Nh/YKrvz8+RXTuhUoEo401zssBwfPVREffegaM6MXb0on8NxOsO2j5bIrjawteoZrU4
UePUxetsKEHJwzqyJSAJ1L+fXceoLhhZ5BF5UEH8EZgXKV9yoVN0wPlEwVnY1MTX+rRyPHNlbVMk
mllgN1AUytqKdfi4nLJ+/FZUTORfjmVElmQt6IMtjHs6TXJMLUmIjF8KNtESCWr9lYrZtjPP40d2
A5WrFv6gyHm6RaqCkSf9amUnyRYaP22YWPm6LSmd4nK/2MCFPjspMs4KEphenDJJ8Cou2DdGLv4x
QxYh/vTOPXy21K88tSzqSgEuIgej8tlbUnQkYxAjnSPTY9nnJhwSfWzhzecgKxjjzTKXDX9szCOA
I3nLNi4iICHG+9i8jT40ubNkXCDne6nQY2ZdNA9K1mWM7RfwRO5OE9tcBWACN/hN0MkS1liaM/Kx
n6K94HIcni2JDqrYCsRBrZ+1DMjt4RzWS7JaCIevjDHMmDW1ATYd4Aj121dDPjTVQ2FNG326uGvb
kOMLaPjCZyBQCfqhLTzk5a0vuxE36y82VSWD0MuAy4HgLOAROKNSAjeJ/l59h+yKswLlAm2KSB2Q
82fk+SWcY3sqYuEd/rG17jKZft8SfyuDVFb5UmbAjPv1xvh7uMq5/2j1AnQZaQDyzYZKh4bLamPL
E58FILQAB1lJhJTAUVmivSZIfuuEgLINhPOhOyPfnVvQ9iwZaR+n3XGcZ75qDAqtWipBwPamlhDZ
SeQpoIcYWt3r3W178KEPGhXHSDZxV1wgfFEMMcd48Qg3jNpqHqMgsx0lrdTh2E59ytZtB2dyXWDl
9vj+tEHELx6+qLXXqDRuYquA7S1tK7B5MZA7qiwsFt0u3Ou96yalChr+gY8aNE/EMK2cqhZnyuY0
W/wKCdkv8mA959Q9hAjIHeBQXbn2wQaASPIc7pqAr+H0N8Hk6r08JA8gFcvA1UDewEP4oji3jYJR
7CR0o1irlpxmvOo2r91KPaVZvnBrKUgaI4NNuezZUIzZFXeMXpBMqbdi7vx/W5x1ohkpoJfBWnPZ
ewn6hspEbIhBu78Bf00ILhaujr99mYkNWlsSPb+WQT18e2BXyjne3l4mIXt1Bl9wVCbLjEGD07oo
JxFcM7DVAVQK/FZGh+oPFdEAK4/0X8UBE1rQPnYY19HndbSidvs6H/0cgvK+ahwvutkQydNo81K/
xTRX7mTTEq2JRTJwdGVNpbNETUY5GjAfspFTlT9qcTn75bPBGNMI8LZ9DD5ZuCP6BogvVP3NddNV
JTwfcpBjvCAT8dBpZYX/s53ynzzZOMlgFwvlVw095cfsq6jT47K9tadb/qKeweVdnofSbPAd4V2n
ApD6nrBtSwWiRwiROe61iu4nZ8T42/u7m2h+3fAxHtmmhTzoQShmcftcfUcXPdqDwTJ/xAbovras
D+MYsEvSI77vJIdpN3dYbakP7CDHKTkDVqG7SCrF4MxYbyAMAgEsIRh2HVfQ0Lj5uDJvFtoqTRVb
pVZdpiPsc1HOnuDHDCZw6qeMtcj3Fo/onO97DQnFnnQ3xfPsOiYcvONZMBNL1mk4o4vb8xRz27LG
kVe35QBZQ9wJt++/c/dE2SkyvXcat69juVSuvHJH8veRah1pzfVjCvoMhu3x3gZo/O1wXU+0pEH9
dPzccZVVbwOIgqZwobQJ5w5Zgi7CNkQ/QY2pXKeaaguLspQp8UgSMOUdjvY52NjoMjsZ+WlQ017u
eKHYhYf9upFHpByvjVOdq+zULgLtGkFI4nFStBFzWzsyWkdukzipPTsyPvVERI9m2A5HD1RVRHFW
M4HMhh/YY4S8r1ZzhEg65WEZ0DOEqIFRTEPo6cEQ4L5jGlEqKD5NPWnnLcIFRpItrM8kL3zUdI+P
S+GF3UD6ol1KQoZXvr7/X4xClIjz+OkPr6h3jCP4ZDWPe5ZVzMQ+q7xy09RBA8lVNIThLhzHRcAj
6ZE4RShEmc2dArxRBlU9sK9w6WzeSj1aVGNo5epMhz45tezODPRQZ6kywaRVyIbLmmikMCPe0ZrE
z6dppzUfuUfW4E9XaRuPmKvHnwCIxOFujnOMbifml+WH17sAmlY8tf/QKv0SjEaBqETngLAITKIP
44XMpYXXxQ5SHX4/LaSexfL11w6Zy1T0cN2w2giUvKgyj3sZrNeS/X4VkW/bANPBjAtQCRECaBkG
gFo0/FeEhcOLMUv+OIaUSKZvAVCRj4epXoEUS1bZvhZrAsaBvb3KZ1HzSPsh2rNNntU4YKhjDe94
+kWr5mMtmAJ5LKXevUsGbq6ZWQyE4Cpa1hOsAEEJ7p/URh0IaiaLB/BG/CJCvMVdxw1ljj4KRYSe
FrlgIoPyEq3bwYv5Dz+RQLjuaGY39/WlFFazqX7XEp9g6MtV5WLrh1DNRxjn6GiZZXc3eip8Vn25
J1KcPh9uzWIHm+XD170T/QEThrmMxpznYmk7I305XWJpyegpz4miW/zlYmhFPM9JhMWqQfNjVqEH
epZpXCt8cecbMYmQKYuMgw/inYuHM9sMkrJrtCzi1V8fXBA5vALcdmDk8CGz9SOBkV2dxTIeCuJI
eObzbGlW8ISkiLdJMTzce7Z5X7EdmNg2p1TntquWb3Y9qirE6xjjlyPSxzvCozCzbY9ov9HpC0ku
0HG6pIv/Gwpol2CrCzW0cY4PBvX+Aw5UCGUhtk9MAhPURhhpkBXHa7XFXWpk55Xrsc3lV+w1iva2
WpIWCL0ESh256hO50IbafIfyE246P9OSrqqBzOzpMpIY5CsegYVVS6qt6vsG0FJcgKDBqrpwkNm5
lm//9r8LI4JU2dfhG1l7rjvcFS7fRByVkzJhOJVcnLvu+5DXXEjf5WtJg1ODAWYKK3oFcVia7W3Z
6S6fk6Z8YjqwBYyT/nti2c5zoj5EmfVf5VPVHOJJZK7b5vom7YVPJLAOcLwKFm8Tl/ZP59ub6dBj
cG1gO9hodRsx63I2DfNj/tF2dS01vF8jItQ5Sm492vaIrEzcPt1OHhww8KWLDuw1ovwk8V2YUl4C
/F48sxibB8NfRRQ01zIi8sb7ekh1dOp0YGClzXoR+H0IsaJUMuYa0O5c0Hc4Dmy+uWgvsUjwFTOd
W8+qxt8R4KvclCvoujaHg4bP4HdKNAe7NQfG/7lzNK45LOR21FkNmntsJIliN1pAJm0Zb8G2vzxX
YLY/qKUtj9lOrTP/a4S9Sc880nTNZxCpCtT6TPOzzdkywuGvjz+JLWxBlQq0VufjJR3ueDk0YYMz
r7mPCskNxVHUqOYy+oYyzE82twLDM4BvXnEC5lA2MX9gTp0TEJ7oUG1l7htMsxvn1ly0UJCbITpv
8s/hxcUCQLLOisnNBUdohbxi6yOy6np8EtJcBQnhn0S3qw9COaVGepNaxF7h3Vd12n1+orcx/hnI
l0LJjy6s3KShK/CHK3XiRCfz8ZvGoZ9VA8d2k93FXhTZBxtI3/W6Pqqcq9dr+S+upxFFeih/oCyJ
/zsw+OayW77AxGv2O5uaGR/zoAk0qqqn0/ZdA4lqsbmcwNwXJsfKmykVOsohrAu0f5YMCBQxbwt+
Bv1TnxKXRnI+cxWPTYoy6eNqYCHwvIvOaIPa4caLVDM6HPGnxqxgddW3cU1iani8RVXV8jXk2Tmj
2OB8kMhVNp8GPR2J97rra3y+ctL9WmqGQfmGbdi/0jxEXJRFmBqO+8X/ZonuYbOIPe+h8/u5Sr/B
R/7AvnhmpavEN/T3QEMu+DVwlsdtu4B+jVNJEhTDaDI3TNK9YT4ajOE3jaOEO4TBgTq2MlUrer6h
fH0bP4v1f/EOgfgg+sIC+PkNr5F3zHRi+ZbrY3KQkJ0cLrzO3EoShLSv76yZ8hr21suLjGLLF4tn
ZnzWAi5geMNGWLFiKy3ZPPTmfDZz0UKUjMOxC7BFXRXD1ADs2tiwLOPZ0QjbQZiruTf8GfeQnAuX
6+OY6RC7GQDWiwXXC4gOSCGZF4yrAVnCOXj8+huCHlGIHUx4T+78H8OtGO2VrA5Pl+sTSZqgs1ke
7O8doN0X3/GePWy9Y265LPKV2Q7Rd9wYX937hHAOrlLIHAlWphtoshQso5kT4IzO177RovQCV+nl
fgUU+IxkxLbTCiqh7ovir8zHv+XMNXR39dR9avW/szPhaggNNm8mnebGAovPt3BRsLaGkuIKNsjD
iMHF2PKWuHqM5JLoRNOiyXh3fRUmIBz6tF5cB9STq6cj2d0/Tu9pnycInhhxAId2kpmywe7KAUEr
nsDVaKSR3ppR5FvA64sLz/0l1hXI/+ypUNstSqd5tK7ejuidgMHAmezmDHJCpiw6NTCbN8cKCwvr
OIcjUXszhoRxD3OYp4nccm/YMMHj1Gbc5jRkTgQFVOucDczz7Bu1zCf7KTYC5avIznW4z6LpE6Jn
bmsU+45aP2I+0u1qps7zhK8CDQyNDH/H2l34kTTMfypM7Z/JDmPJFRJ7/yRFWtaVXrwBbW3AwAD0
5Dq3ugE8UJaLOb9hF9bG+ObAXJPE9dmeMUh1VNMLISO8eVCTGe+WkPcbgcAyaMdH6564VYuCjsUx
Q3MGBJsW8NPUibleLpY0f3U/g1t2aoi5SJPiujUTsGDzzpy3CofVO+b4RkalDoc+ajgRP5AU/LV+
tOhBAdvohVb32A/wTHQjtJ3auh/M1hLw75HbE4pfhwGO2KoE3BEWCsR2XvB9Ky+cjpXALmLIcdaa
cwuYHbPddrRxUJeHSU1k7LqMv1QjUZFpUWUF1Gj5vvzGlH257nnNFGpjWuvfIii2heZ3PjVhEKCY
mGse+6F+yPY3cgV9y5Y85VFOfrqcEkvDvvIfvsqDA1SmwVkwWo90qOeI7o4rICkIDgeFwV6Ul72S
0mjlAVvLANP7+i1Yj79MzAakm8xKpPfaGeUdAWjTrdPJuSRyyhNx302dvgoXy3SJ+TPH8UCDLb2I
eFhN5OYRJ8/Dv+6auTMqdM5sC6kjj0qhcngZfsQ8pmVftmfIyASQfQxm5dHmKmnZLkJOLFOp/7Ci
cNxRFBWZnNm3VBgFk7TOJB7HNKj8UESWT4LOHXPyeGELfFyPWbbpHcXYg9dAra77/EpRkq5wl1t9
pB7ilZNXwOt3I+2PX3XmFQbt/LnKIbWdNT6l52oyAlR/xnk3XSrxwjjoEaNmL9m7LAsL846Tk6NM
Dsx2NyLUww59bsXIxthWwRYwDLAby1pg+q9QrswamUiraTUwapyO80SWwcXGaRMBVXFWin1mHxV8
7u5krdz5N6sHAMvPJ7mYw5aqoS6y8U8hyO/CjukpWhipIePnlyiqyanrzBbpZCLUMm5WqVqOvBYH
pAUpyKmZI7kryBhGUdC8axquioHg5SIA8O+FjUWif5CEUfqnnqr318Ls+v4RHwpfegqM7G0WNK6g
6ZOH6p+iRvEyHSd2uvFVSasE4HR61+kukr4rC/iOdvkts8iwJqofEzEmouanRzFkMytmsPTxICRw
hkSy8uihoeYbESIXa01etKSp5FfmA1QHwmtqGcTGqIgp7DJo92f6M2EJfnJHA4id0Fg7WQ8H7GVU
fzPpTAcDf64FladiYd6WrObmxzUX2YuvhgsSgqn3QOjLl+kQ27RZ6KChO4kjTbmsuX4cV2DC95jC
qk8dc4T1lmLns2XMZiiU0ocS0wDjCPq1I/LBla8vCKVw3NFr+KFWKVbqpkryDswM8UWKki/VlA/p
kW3i1x+j/5Mjd2hRC1T0zKSF3oLkM6CG2DsQK5HjgcgNkhVD3lHHXyssCn50g2vsBzqQXKfRP/fc
lN0EzT3GxpuyhY0isU5z2GbMCsOaVjdVLpIzezctKUcH1AyPnnDPLFAWXE/cpbNJ+YoE3YD7oBty
YFvPbYS9zJbVqzh5MMvAels3n8PGEiZhCbGb4TMi4hVU5n5erd2v28gReaCb0/PcOPCaC4s0jcYY
IzxPHVZ4glwTXf2kytCfz/nI4JmxA5o8qThEHmiwcytJyJ53grZyyykL5mb7NFI9Yc6MCAUt+Dmb
ve6vDEtX2nt86tp9Uey5Jz7J8Kg0cYYncg8GDlVoth/ee14/OS9g42kixryufYN08Zmuuma45ssn
b6ZwObml45YI4rxTiDVhj1oly3lk0s9GY6ixNYOnfnxYmwRacaEn/Z0XwoTUfqCe9ugdJ4bVf+s+
hINpHjkeAeyR2zOMdq/AMuKb8KvDT53v0zxaRVoEMyXZKghihrTHxDMx1L00y4LC493gFq7bqqNC
TFiMcWQMgtVXtKSSqNtZQ+fNPWiNQ+iJ7IVxLjnUFnOL1mq2EoSN+CS+kgX5C3QxT1YTJrhkkDZi
ddvFn0VBkBBKG2JlmGp9+dAbDa+zzMPvZi4YSIIFTLOfdtLjw2EqRTFFyo7aI1h+4MMQLUMgUzYg
FKLzHHaF42nTHsqEOKSqUMhef6vFlt4It2S44nxEE8mr7QiCExOaaYIQQZ0y7pBnJEC9kHC+6ze9
o5QEP8mopMJUKGI0Y7URhyRmFgNegHzlW387hcoVeOcI4/p/SvK2q0Lc+CRHhUWNgPdDtc2JaZ/H
1rSZgWo23v4NavJZ5oTSu7Bk+oCRuMg64gj2gG9L/BHI1HbExd+R6fZWnhfuOkMl9PXXXYoJFJd9
0boDvjL1bCTKOFxer6t9/nqAxyh9UrP1eUQIxeTRzD3NpX2kq4XmhJgFZK1NZPgCfi9YoYd8dEEh
PsJBhzqcjFwaw57N/3ClpV0UtDQRSpc3eSoi3pCQRUqhfLry0wu7Q3akE+W4sv2xErm4ZwdctvSw
/9JAXaUBAXrASDsjWOBKWqpLdI7XTnzbHXe5f19MUc5/0AwYkcfbLbNQvdz4TNlyuGDgBeUUm+i2
Y5+2fZZQzb/MVrhGs9mMlFYfKCILhrX4kdc7RAW4Ts1l8IIdvqwxgwzwxp2Aalu8WHPoEPeLZFV/
6QXVqoDwWpt/3OYRrQIsjDzBMNnLO9FS9pAGCRpnIlxqmHcm77FpVg24xWqFGwBpgN5dxG0mmFoN
7vbDlDoE5wTkQLxsCFIiMM0CZMhcZzzShZLt6L5INW6v4ktr82Vc/Pz/XCwRjM2qy6HSgo9s2JVd
zxXVAITdzbvt1o6ZvD39V4zZ2VqYvBTBYEpttA4r+c5XfbOJv9BgaOAcHgdgW2OjY6Oy3EcSASrF
ZNOLjeVBCRzp1qozMVnnLlzZPj2JLiYuCnsE8eiuIYiwcQcjyYMLzNGjtGieHlRvh6j0FQXleHo+
izKIHUDSvs5C+DHQRlHzPKDskG4e/9G5q9pGlA+c12EeaS6zTYMqxIHlJcaovu7RLh9gxSwLNj3x
3LPwDsE6fUaVTLpoz2lgKc1NV4F65qoyON03VdYLuc/ziEztRFj4G8W9EW0ybGxQ+KE2v9h9XSd9
Y6nUSZjC/77n/QdjQ3VplBpy1wxye1Rn3yImW1ovrDki/KD/HIXo8PDQHOQr4xzAidqItx2thafI
GhLlrArXKOlxVr0FYVy9xUPZDAoeNnme9fdCRzCggEMwDvZR1gHuUlMgvAkfWQl7nKsUliSLPLzR
JlNY2eTZwgaVIbFQO8mpaUorB/SJQtFkvcz0He2RWEWoOfhnuGeywjr7Px87Pu8whj9P6EulVsGA
vx0eyls/D8dgmoiZfPXNQaTWovwXIZCoZAFNv8DGMJqp4nx1sy7tR/wnxzdg5wj47Z/b3SjjAeGy
4KzthplU/imyHlqWog/9pCEuiG2a8XrUJcXP8UNg0Vs/GrlAw55/B2hGIcjyOhkIooOh9ry6kTAZ
FZFAtWivW7EBDWSL0oyifTsB+KnPRGCNdocJtDOtFXyWuBfgi4SE8uBO96pw7yVyhcf41u3pgXyK
ZVb1m/h+EZ8qK8eD/6aEabPzQF+tjTm/EdT/as0pobDSPQ8QU0DUE2HeRiYpBEJB2LhOurdcsWTM
kWrT2HUj9N/ZqcvyOrHivVqK8IP4NJE4Ke8JZ+W/LBN2GpcgcCU4Vo+4m4UlGgFSMV4l1pTCQDBP
WXNjC71+swFXUu/YdSAV7CTwL2nICgkNXZN2qoij5CrX6gIZ5SN/FVFql0DDpMuFrFB7v0HIZfEu
atB3FngKhIy1rLE9TESxgIibpd+NiQw8wS32b0lxyIfp1CW1GnzlO+X/JpkwTi3w/66Lg5ICTNhd
+bpgoVaES3vLLD5TJzPv1tj7bUGrjweSoOZ1NnkJ3HPnSEMo3PurTMky69jh5wRJu5/PRlqbrcqM
oy8zo9k1X3RhfRs1HT6jQ0vDPNcv3WNhTnIYjwOsVuru6TK+BJnHuLUuCAqlbcObfOPmOdGKd/ck
uh/iYH2eYN+v2JSNZ9svMRkVCBi1eRKW2ZUOlgKW1n49Si7qvOQZXgGa8qx3oUrbkkIegWQ4RU0x
vuSOfSeJL6OupyacfbXm8+fLvP+zWSrGru2bYEqvmOnOklWcvjQ2EIbVnjONeT2vDE9QNvFMUOi1
lpVftUB6VcliBEFcTS3i1rx2o9F/4k9+fOAlJRDuA+e/qfjZnlIJBjjoILxiIvvv0NI0KtIfhC8f
2fl/f7PuAO2hfNCfeAp53s0AtlMZdase/qGvBYlcBFkaW6QQRKessLpLCCuCQeHApyd4/IPzhQCc
PmF6UoZL/rrZT+PGWrGv9rcq/oN8T3wOcX/7MWR7qRYdn0uxhzarL9ltCpsTL26hvYQt+ZQCJ2ES
tgAQAH8W+6bId+Rn4CFX1sggzgUTwckfwaM7iiICzv/FP4ZMRUbY2kx7kVoZ1y5UHVNQ7XMsqIFW
NY+Z0vN3fsfy49tTIaMA9JHUx/f+8sKM86zlcg+3EQuZbLz0T4vUgt0z8e5E2D400q9i0qGMIqeL
slFfxz5cZFNPCUCWS4dX6x7rLD8oeRud1TauDsnAOQfdlUyaiDnb1ccWXqo1Rgf0S3Y9J6FgdEOk
iTyNj3iGrPLiTv09STK5W6nd4KpJA5m35X/3f/idOGVnEyjBKqLM9VwQIOofu8lPmMWFtO/l+h4T
v/o/uoiK442R8pQyY/D1LIPLd0STEFEzrTb/Ra3kdNEGEcykVyCKlhAApKVOeXyiugT9DI7Iekxw
cYavntkIYVGaHfehJgx2Kle/FKv+5kNRMESPUXkUZuVpfMxTyaBSqnC4leo0y0QjXMTUEYfY3adA
cbfX0Mk3X3Bvt33yGYx/yZNmWUh1qmhJeRKpP936v2/nY/BIdgmynQET8DVKZ6STTq5Ala/TfWS3
IsRuw1NwoVa4moZcB97AsxHEEifqZxuTdrfzbZ2Lz3bSmGisP9dYutuNAowyIrYFhNWaajTehZDZ
i5moIcrycBFioiFeaMdjRmEvrmqWAf8gKBXZkSCRZr+TybinHDjvSLTLCzYsjlLsdOR7l6ADzDsV
jR0RI9+TFlNpHJnPPl4Ttq65SMMyq7N4F0P9JsvpYyK+mAmVE+NTfNvL4Lk6Ik1ER6cjA3jbW1b1
/5LgTnCSg9za36yp6vSkTIbuc6JAc7LQQLM2AlbB6yv81D6Sf/BABTYzkRdgZ2NXq5o8ZOaWWHG6
eHHZy7xrMy8lZrLoxaYeoboJVplI4VW1PoP5AW5kZX4l2Tc6zPiPED1U80kmlMegNNF+O1VXgaAn
PQcL1smJm+Q4kt84OytJ480PvfG2WgoxbbTTAig/O3EZ3Rt47eIe5Nv0kULurffH/T6s41lvWwOU
xoFyes4o64pbN/jf40yvTBiz//7cIZbYmtq6M1jlKpgERW0FPaBE0vntAX/k2AZsxQGfizd9GnCk
a/cOQ2BdXlFjODMdpIiXwKXzBNTiRJeW7F0PpXDMe562SCny/hDSi8lRBIv7ZccRlvFPX77/dmLM
bz/xbhXulYtVHsZLn/XC+OD9Doeau6IxnRboxH3Vrbbz+7QIaPdoGTxXZXcyIuNd/0ODqGwUILbf
P/Ybwsp4x7QkfUGhJ29gQo/93uPkoi+y7vQZDTrm2C1JSFr2bFav+f0FPDr9efgp4E7Ua7RpqzwN
MrlfwtA/lOHVlPCnL/AGRXnu7aSV+T8tPRntWOtK/ukKHDR6nCrtfoFWY98k4kiBjP1yCUvptU3x
6qqEr/2oaqLei/O1/xgIr6p7Dqs4fSRAduHkXp1cWI7Rio5toCVQ47gXoHAKBu6bfW0fK3pl+mMS
2FZAppxJQfmNrcbZXPLHi54eq4bQ+jwcVBXytHVrg6mcxi/F/UjtcY+2ngfUKvNZwwCu1f7sZOtS
RbWBy+iRkKx7nR9mk1ArebOA99QT+J+yJcegyS0+F3MHP3+gfi0Q2+1jVbiwsvVTWJTN4uUOMNTE
7AEJeKcx7H9YawRjK1Vam/V8rJdqO8h9ijyOefHJ3BuVlyg4TtqNALMpqwcRzV6O516mEiuz6mUJ
nar0UPuLrFhJWaMy62HJ95UdZPgGhxh0ilwJilPB2KZ/lWiKztJ01zbyOFl4KSjLTCO9OtQ97W4Y
fCdv+CoTX6LqJKCF9fxIqSJWr0zcSuL0K9pEHrOsrUVpuqAICRCQ1Xl70oOkXqEs+0rW88hHBM5v
/5UhdAm5qcWIu/2Qz91zbKyG5kYC3CzGwaSBKVb5Y0C+ARPvPnGPglTdJDN8u6743iaeO+UjcSki
9ZAMq0+W3lpWbj2ldb4hF2O7pjgoJwHc1o/BYAnqBd2ispK0cm/z6hBqCNbrHf4ET6EkKIdgdJqz
zuY55lTRD2n6XDnZUDwXAabM46Rhlxu2T668MCZC13O19XZyLVhzJjytszJKMQnhlxdobSES2X0q
WjrQLx+c3Vbqr0VrjtitYmrBkOjg5B77ge/MIelnjnozN6jeWLwu6B1VmC53JYytiITw031Bksur
T4ZRo/QJRejr9UYsmAnnbY4GjwsjHMmaCp2bURrDpPTsjhCcI97wXQoGXsRaDH/AKzRNPbavsY4c
z2HZzGEGjupSujAImmRD0g4VyfNhOXQhr11tI2l67/7pzY7+7/QM3WK9xQEgqmiLR04P3nFhr0E5
RkfBWgadCgor+kMGPua2t91rpPWSTRD8UVYtmO8olM1UQtih8e050JBwhuebqPs4ZDhASXUkRBoV
8sPyQO0HW7tJvM2MY+yz/cyzu0vdXsyxjUkDw0NkKm1Wn/CtZwSc8mCVDr9XYXUYCB0tOWxzamz3
lPVA1zhjKKYufKSh53ngbtApuF4O31yn/sgY4MaF+QQsWL/nOFDiTn6JuqMH7vgfl0Opv3pfkrZ7
LChD9omYl4M9041SoOtSstRb5KW04+e/SqTJyVbZ0dV7HTUURJnRRQQwVk2cIewpfIu77YEaVNHN
vSHkZ+UqINlZlb0phzxbtQdqUU9TjW6qQZQ6Do/fKs4bL2GJ57mC/fwacqTgN9grEXwVTlRVsAGm
eddTEWsvX/4WvgzKS3eOY7Aq26fBDn6GFyL05WMnTti0bOot2ybvInTmpddlZnaJOsRqF3Pupxd+
5vOyiTc/+/ByKzun3tXm/db6A/f7NuKj/5v6XMmafqyyeYn0IO7n5kYyJOt+6ejHqwpzMIGwg/K5
7R+n+VkOLBSlqjnlB0JhR+s6j/4lmQPWYnbjGajScRv8kMxKyoL7q38LOUqsjf18TO0uq800PiZ0
kv0KGbHOLKZguCnJNXbJVBMhO40sE50slExuXLs8ePq/UEnrpNqlU3Ye3fbYHG3NIpbYhe1Op91g
QG/WIYwcMKN9ovEG3fUzTg1asWFkYx15SxcSsfw9bX9B8oa34FoHqPk31w4yLmKj4C5gvQ6MiqqY
s60twwFsJYzcQSLYyb/tqAop90S5MO0CczbtjFh8BjcWnitrHNmFPugiXmOVrGVcBPdCKE8rd2t0
g6GSQdmgh7yJOCtnUhqpbIFcubxME82YYcmx7KckcdBp3/hKa1NgvjcacL1jTWXJFGUK74ySNlU1
eK4672iev+kzZyCpWfV3Y1ycVSQUmv85JBOvxGpZWeY0zKxcSmufC1WA7Excax0+divPKoOq3qyQ
KX8s5cJQTx1tVQLdJCOn0lIimJprIGHL2pb6phlnY3AkCp6wllQUe1t/Cnh/lRILtJ1vDzGXSdXQ
TbbjAoAkoCZR6R3R2LnNtwHFSG5IO3PvOuY9A+UxSLGV2zyh+QQ8FQte3b/yejEhlze5KW7MADlE
gW14q4ZTgcUfT0RLAZjnyY4vHcmwVgvcF8P0jpPnE3H7y5zCEZLkzMdfkBwoKq//DPw8qAqMUYHE
zJzDUAn0cTBOJKQxlRo3z+NzgmTydSk4xleZWhutRThme7xQRxEXDgUKqDcmyGt2f6lf9aNkEPI1
cD/nk8/YVngeT+TFOkC7nUbnxBk3XGxM5xGSFoKN9yxYdMLucrzF5PSigtQWOFhDnI4Piv0tXGsx
qiredpvfysYTLIV04f+6nqSDiEZr5ZofaXQW9BuZLG8C6q4vOX5eMmlxu7sWsOMHKkjsJFoU6h0C
3MSc3YRDFHf8h3z8uMU/HnuM6JcW4Rtp4JLaG+EcqHu0+5qLUFypJFMzbYvnl6Wjn78XUk70LIAP
JiK8CARsGUPRED07Uvb1934J7zXnrvljMvzA3vWfXAJTkJeocZ+UHPmlnXigMy6ki1IhOn5bz1tj
hSE0rKK3xHrf3n+sVz+hYDX9cbtCEDcW40Dw2DaJ+xIzlfE7xMVjAmu3iANghftKvu+1jR8p8d6g
QdlVbHLstg94DseU6nhFgyK09DW6oFmixmRQ4UDHt5jF6e3nARP9ITA/ZxLfWGMmVOaoOSdjz+on
pYe5O+g329cT7hT+ovfn8G1wqsDZRUDnp7H3FruH345XPArU/WtiGQpeVMbRanXqN+l7H4Gy5Xji
PsdOeBVT9AoKk+zkv6i9MKw+iZuBxvVtcq+BnouccxlHU3RJCGxTnqGPPMU9AoHkC1DhDZQKXbeW
fBxLIhQxDEsCuglxXG7/dQ9x3sR/jERE8EejFKaT4hqKS/DMWDdwdArHBcZAEX//kbaXqY4qQWkR
cqX0uOyKFImT/o7KsXJo9vnp6qp//KXajt6U5owD1nk50Fp2xX1Wk+wvZhsskr2XVclZ2X9gjqXs
olJzKFbefN9RV3wMD6rJTKmK7MLqtPvWvmw6zllA9p8dbwyqtljQyig6rzGGjK5MRNaYBtX46zPS
RS2gWcFJ5gzHwuQsMTDYhOT/Zvm8RvhLRoDBb4gLp5MvO8DdqxAVdL4FvWGpkFXPbtiYXW0aEOOx
4lF3g2jvuktsXtuS1wgI/DDC8r9jDYEOdOPtD7EokC7qG93snDu/Wy/6WKeknP8Xd73KHPTsZ+71
haZZusKI4nDh8daGIk0X5p6ZThBQrwivVuU1mJywUl0H2hB/KzrRe6Ulp3d9A3/EGO13RisAaEg8
IGMGGIs3gDEbE0IUHHCpvFWsOFdOrHXdUj0djXdbud4yv3S1j+86nJAyrioIJlBNrH0pcN8Lu6H/
q8lbv3P9sH4iMkjSEBcFb1hOLJDClbtwGY+Yia3g1p7liL4JJrR+zNt5agsFLJjZ2CIL2NJLp3MQ
jTvExuFvTO0eLyK4PxxipHV7CSmuhTzlvpd9tCoY8QR15jCTYtj0iAdXcM0HaqgXJ9CvXqKwBvW9
tX1YpV/hjJED3K+oDYQiLiykPf4AyBmuFywmVMragAlka2y0QHt6qpmaQUTNfFAKp4TKhOimbM04
VYALNawJtIASaVMXmuWmA4pZa1qgejNlA+NN7MjEpjhYKL8IkSMALmmK4eQ5Wg1ObZOVCEG3agis
dy3ORc9xFUZVw+NknS6ojhrcMPb9B7pALwCqu/n67c7UlBEh4BAATyurMtHzmZ5QkUeGPcH3hBlg
j10qwHORQBBY5goGDEx7GWSbLsiBCOIv9VyHCS7RifYpxNIb9UFvsftNxN40updItaKhFuqhXlh9
DFG5kxI12gLkbUKYztfH8nwdB8UzQ1t93y36BagkoiRyH3mg5LI+dpcqteV6frzWmdZm44rD+/Xl
NbJScVeXY1964s4kQEBSpcXB21QOwVqeLrYNrxHPVCTOcLNLZ5hq0aNiW0zW+DEnR+wPcbWNnyxp
VkxEAZyXlmjT9uBmjcCGaEc483uqI8ImYe/r09Z2hDSLfG068ooMp4ug6Rb27eACNtF6q3UCXCNP
9/uryyAW0qA/hBeb0ELrz3goJhbPjB+1CUCgWcdJJWXlAv0VknsgikfO1IgizNyhWc3FqiDbih7a
6lGbl9omIYQrdjUzexkWPYgb0/DW5fLJU004J8o/Fr0FEZZ9uGp10cphiRHOliRvd8LyTzq+v21N
Ns/ChZwYYSj7bvIO5bJXimIQGPlzHhkmJFxI7xucF4k28idF6uVjMRfPtOYroTieW7F+Sox12CO8
WbOeaZEaJ7gVJtfHCGOtbu4EAJcOvtwGGXsfUwMqrQ2FNpQ8mRmD5G+hz5pKz7kIUTibxaBjyTXE
9pzhYx2XXEmoaHXFe2Wba1gs7MtCTbjYN5jdZ+D+UjcpSpZg5q0h1gz6IIWjZwZ+3FVpvfSvNru+
f6nFN7cNRNoWim00kT+EGCToZNNTlVC3Y1AhtjfFvyHqdKmhrZL5hGvtGXf9RCCcxTfe+B7+qhCa
YXdqtxOsyJP2SFPQk6jbpGtWzCXb48coI/r8SYAzbVDr98qeRihx6utO+8LuDGCf7E8cY2eiD+AK
gUd5i9YtmIZRgqcLt+7FxdGOo+PJlrkJZQ5Lc8gOMxH3a98CIhrdSY06I1E3jxICqyTMkhHSFCYC
3fWVyH1sD0dUnJyArtWkN5Zi75WWNASVCn4kp4ERyRX8pbA0QcwWi8Td0BZ6fhJG9vpg8naZ5fp0
iXtIiwLCGDFaeXfaXRvD/W4HQro0jNa8uj0ic6hX9S8fdcLFy0hZ+re2pl64SktUutX2KJxnyW0V
s19B5TTC8dy6ipT+qRt1GZe+uBksiLCMh9TT8LbUDczoBhTXr/i8EwINHtMQY9yUqm2upEvTSUJz
NqHmjiRX2mTDYFcGdiBRO4SKQkHkXdmK6acXYQBwlDUpvZQdPxfhcKkCoB3wGalPtUS1SkCfbYu2
r7Y0QqVhq0kTwqx3BTrs8PfsneNB108rHJPd2+ozlvaeGWcTtSRBBaoQkGaIJQlJFmY0m0EYQndJ
vj+AfD8cG3qbETJbnwdTu45EXXBA5abhZNRBtZhuMfd901tyJkWe6YH9UN9bsfh52B+dd7Rhhtbw
gtyBvPGwYzmZjoJjvrP9dXSNZe7ICotLajVSolmegqBTlmhN/ApfukAvZWeCHo01FLQI0cWqbG5Y
9Z4uPmgApbcu83/zaF2vug0RX63EeOWFxfbWBUplZsxwe8uIbWiST9gA0Pi676nECoGuOOo0UdB8
qsQkgw2D8if7b28GJ4xx1C1mtwdA72DvI8kIklAlJGRbQ6mgbsqtsiCfh70ZEA34fI4Uf++8Uo/c
EQo9lYVm/1nfsR14+SqnR4xa+OntZBuDyO/K61d+r5L7z5KePh+xxTacYkkb6N9wseYhJ4QT0/yQ
P7kmQMrPuHALyCpJYkMWMyyO3mMAsqRaBfta3Z3ATqSmt64rGd7lWIxJuvBwUvbOZrdMn3q22UvQ
bXbqfGdyHTFEcNZXHQdAMuwVyrwpPS1Y+CHIQfiX8Dc0jsV0OKYFlozNab8tN2Wn1q/8tKubaGbH
DABU+B9m6WyKxhmtkgFRuboez/PmTl8PTRTkaeL00+xVMa7M6QeD2GJnxwLMVKJo8s2RYNVLAvu3
OYL5WwPANUTK8j033WOLCgTAvjjbCrATyfkCHDV9ajWcbk6wr7UMhfE3GTah4txBuQmxr5oPkLk6
YstL5167VNNPlKIt1X4vc8FQIHrpnGrHTjpcQYmsyBgo/IOTto2LgwfNEoGNwhaG3W+mzkPvSiOH
/dNNwMvQvQjXiBCWr/aLAFxg5M6iV1Qudph4ZRskrtr5wXaHYbnl1Anz/N6u8/q6YOsML9EBbmNQ
rzZG7w4l5EDgm6MLByWcrJ3cjCo/ogfH8I3axPYtPwuYVH3zLY5TTsGf1LsnD2ibmj14aMLyvYjN
xQltK5HOF0g91+Y+fP069lC5+68rq4nnnQNlO1obR3tXngWngb6uB9D6ugUxgaLjjPO3qQMF8wiV
0rTRkHHm6jWqyXESt10QvP6WzGUOK5NZEUdZTbEVyvSxNKtDqwMCXrz3nr1Yqje/wS9xx0q1+BiX
ZQsKXzR/TKFB+p9Z+8AQ03FEAEs57GJD4n2eSL1Cy0z3OZF2FL7uh6F0mLlzHvJUQuMFW8C3V7nI
RK61t1j2dU2+bmbCK7jSY/Ok7LItGOTPDsZMYGlmWcSgxhud5fjuDQY+Fi+3FE7vwdnlI4SP3HQx
mA5rerFT5m9TPg4Sx4le+Xc48cQJ4ixv6o8W0ZHy0TxgOn//rtJTMosQCWX8tXs3lGJiRVmj5/Qz
oew7/CWfw2DwGGOLW/BT3lX6/6tFXOLJ7BEjMeri/iq8SpN+UfCDVOJq2frK0Q8d4s/yZh3AzmXs
8TQgn0WY43ZA9szePxuBOrIgzq9PGPTk25Ei1cj3dDYd31Rrexpcb7z7NaqHdYL3610YB5aHeYCY
Q8jxudWCgZnSs8Z6EKFzR0Q17parkIbTZsG703GB08Yx3U0JCYDplfAAXeRjC4mg+7uJnLWkMnhA
WMx58EreXSrPcD4aHXAJoux9fcGgaUGxdB1TEB1JwpCHsooFV05nXsG2ls58tMUhwqHivzIfvTMB
RU5t0xlrdVqdyPrNzr59ydRZ1+dwlfDZJexMxkpe3yzjaUWhKXs7hIqqtxmnGO1dhWDNm2dyUtnz
+OfoRQjrYbai/PEBAPrvRQnJt9YiRWxYsw1/5d6/fmhYll6Q33i4Mf6Zm9hWCCZZeT8XDZUMLldB
+u5DRXCGRIfo7ZgN2UZj7FljM27Wd2i4UZ1njELXtouggK8jp8/fIfK9+BM2KnehkjhCUpy4qLzo
O9GwAJlJIaqfv7hkQyYIidlBOM/BB4nxaECuu9r23gfSROhBV4vyOZ4nOBOc7T0Phiy0gC2XaA1n
Lbf8Twc+PNKc3a/OP3xBSZomkOKsJq32pVWJTksmUoXBVRyuPUQrBKbdRRXG+hOixBDf4ZcP1XJS
XDIC/9xWCz4boLBwj2Fp3/0hgjVOqAoneNlS2pmhPHPjfYcc4UC7B+O2T2Jqh5z4NVIH0qUv704M
tAxkdN3+wxZfZAwichtOcCypli44/Im30HJwHudplknwKLzse7z/fVtKI/D17Sz+gPOzUKo1Xn8l
mE2L/14hHSDRNAwOG1o37scKhm7JcRneQOe2IEAxEUdDpkQeKs1e88TILtDCZXk463xVjoRZRbpn
mrxk2Qjf65rmDGK0aJFCJxLYMDWuVdVxw3crRPo0wzqIHl5g9L3jGHIATEr/gCLaXs6LyvfYPmbN
prTzWq1QQfk7AR1vABu5Iki/pCT1LVRTcJEK23/hUBEejofLQF4mY3CsyRspEQpoc1Nt1BgGMzUG
5beOFxF8JwRziR5oqtUELTHDGH0n/TE0jUdLyYVnyjgbHS5KlGbooqd66erzgrg5bwK39PWun9+q
AJErJVXJ9atE7FJPzKwiVzMClNAC+il0Nl3pz63G6uz4GoF/8+wGtODJgeapIRrUuWytBLT2CCqT
lPcf7XxlAnVb2mmzNw7YXwn/IsJhU8a5Vyv7YBOEdDLmeND96LGZ83oZ7ItQpbr8MXIBjqiebT06
4FdivES7Hq/lfPZHSPUn1iGNNSrSkMdrOWUDrHhefHyq38AAQJJNWAkWN+lvNz+YlY22V0+Qmq0r
YjMwLKrZT3GjNbWyE2iZaAY1el/96E2CqkX/Aserfc2JfkQ16DlcU6xMvsZfJwy5YRjaBggbtXek
fNB6j4OYTCyS/kztC7LMOqvC2R6s/iiK6y0cEp3YELZwuvi4XRXeL7YDxrkWuXOojK3wIgOJX4BM
2CQbHDk9PVxHhUOsatwxdPmj+nQqCDHWFwBOt5x4xR2SVH3ctYSQNoc9Wyp9K+L345YMimC/4Onn
c+107fV174pWKvICc2Xr019pd+nZVkZ6iguaTPBemcn61xW+ruQ14A1YD76+kVXrEGVJqQUAHudG
ne8XocQoO3j+x0cMPcjqvo5v/39W4qEoBUO53iLyuWnvB+Mm7nGGmBTLJboCnGJrTZ5S6Y7X0wcT
UohbSdlFDm3hD6BIeR9F9D/EI1ydaLNdhU/6JGdrOjrrBZD369LsiBHMg/ebmK9KFRbJVtLDNRyF
5vIe6m74gKUQEl/KYoIzlkJKD6kQHliQQxtRCiuTYTzZMw9X4vgYwJElRMPRE6MLooupB5C2wpFP
CiYoyM4ezxX4Rrj3PkHDlhgg8lFgJcZ1ZYY0+aVpMqpE/dZzMiqjqKVgk3Tf7xTt4io55LQZUGt8
6FDNNbg+PljbStC4f6T0XhOHroBkzgFXcK6wo5fqsLN29fTFDB56CyULdfR+nwjfep9cAoA/937l
S2MEbwD5/eBO+UmWf3wAqxq1voDqyHHkrhZqheud9T4OG6guyi9SD+i2x8+guBv8VSWVeYkLNIr9
fEca8NbRoQHuQmonZ0l47B5BvASX+bnVTtRuHYB2Ot0PhvNO/XABYNtcO7S43lcfahBnEYrs/BPD
SIyPwFwBwgEIQdFxXb3oI81597VeQt+poUMBSYJZavgxE6lmTPG1X3qyE7ptTvccDtl2QGgdn4xv
x315wd0TIpiSkwBxjzLGMgdmorwW3VO+hhG5HNj99VSjoJJxaEkHDKJte5/2jDB11fXsom1FbxyA
79PfqZ7lMGOcKbe7QoCtxRRLFngpr7dbhafxvdEwqY35sGiYtXtCJnuAbyAtTkomF5NLELYA4h37
0BW220B+f/eGsujCyp9MpXAh+P+eon5iWX4GShM65Ac4MmGUuov5fNFsvsZUcP+CPxp9NYKvsEQ8
jdgnln5zIyPB6reGzQL0B0SfpelUZ+2pIUbHyE2VQzcaQggR3qtpri2oTsAp1W8q3LO561ik+VxN
qqRijDa+1UIuwROapKVW1jFNaam+qk5NxPmT8jcfq2foicuz5vxkpjQYx0M5P/dPjfDrP6oAHn72
iBznZ9zgmQkUx188WY4S7QcLOn8VSz9mQkrlD8hMrgcsL+tjz43C7ofs+xeLEOSYzC7RxIbSI0lV
+6VdZu6pf5JZ81GMTl9fnmoY3HluiUMeLuWbt50gbW5XADZYFBWn12WSnPTuODDGBAtIkZvtJBk/
j8GRX6sTIR+JvJx9EHwBFaepONrwzloCC0LmWGjz+BmCy3aEuvITAKEJkMc6nfwpYbQrfkxXp6Fl
22Iv56C9i2mcnEGJBKZ3FdRkjoy4Jr787/hHDcSL8zmNNhurdF6y5W4+1oakjVn2KUQKPio1CSI2
doQqIQhVd2My3JoCtUsxFwXjm9wVkxID/UKyVwItD8CQMynVhcEQwAd6Q4hvdT0qmXc3ncFGT1kK
JcnVIL3wO+Ssrl8agM8rdhKScANwmHsfow14l7foNs0MFzBb0yjvNqf8XOT0PNwklJemEDgSBgya
dZoYXEep67rQUyUuKdqWIFzDY3TZ4YReTWJHgQbJFzPvtS91Ev8JcxLYV5bFJ7ymW0/0nT5IPwP+
mjPnLyjGxGsV1tBgzh8sHF46fuavZo3ZEcXzMDTPtx/5LeNoQfyr9x8U5RhBqUPi+n1mpZf1Fj2Z
Iz4HMfigGfa7oobq5Oxlxxf+siprT6zCMYPWDVEDhvoDO1a2GEC96auMB6e7eqq8x7SZ/TjEXcPz
nBTVIlRmrKuxHtP3FKhROJJp5xDbtPG+Rp92oYf8hhXtZuLiScjgh8yq/wFq39ckpDv1KroQ1OY/
AIHaoFZ/xGsycQtIA1NQZaTfcMaAyfFhXFg4JnJdFp8MRalPzyzsk53q7jPGXK6qcmQdgEfBcT6k
VT3UYwMsHTqEHTlqS5J9WXv2eajG7S5kijOUX5yidYV4kSKDoiLlDvuVRQDmfXOJ0JWGtNLTC0nX
ugyOj34Q4a0ay/X0pKYFiljlapKIeVqGTPvn4KRpVn43lwrOFoDimPGgO/ujJ3x64tvv03GGmd7j
WuUlh+KjwSdcuDdaZq2FVMY9KflPw53RtiDX5KrW18BG7E93frhI4gByls8kBRYINrRuSoa9NK2K
FIF4smYseAlW5H7cBWPyTXPKseSv4McQloi4N/qbQ325NDr/KOGKhu8IotWLXC0aimv0oIP/iNc1
JJ8+BNEVXrw8c1eRGrmhW666G44mDXsEc/Q+GP+IQADKld13oB3UmYGleakpb3vFZ5xKZBGO82aT
RsaS9ld96x5QOGsKUSUdhv5u0x4pdBt9QYJ9t7f1KOo83teGKwUWLfeqlkOs8XXsgu6xs71eAjYW
9swFL33WuR8XmH4Oy4aoLtplaph5llWKHk1dRAeMxsRXRv/ER6a/Xgie3iCCHSIOgjWk0X/foIhz
9Qa7UrtuA+tPFLcHYWgSrR6FOUu6IJuFwrw2bG/tA11xRpPwEGZ05mw94uFF+OhqpF/4+qkI19ci
TZziUIVbQ7URlmGStO70zJtBA8Kg05BZbqIfPyyg0ccicPAs/S1//mf4JFAnv5Eg95hkiZRxDGdq
pUGDKy0jHDhpj2t0mWHwO+oFtKl3uS6TKacIxF1rWorSfYftpcKI1kG5SKB7Uww90aqWVhua9eob
mB3WgY6HWKIJfUtrGJee+9FpX7J3usNOpXg4Hzr5IGa+elwtbyhV5K+WeoY7iojEarOJAyuNHO+/
4/nWafQeR0OAMS40oAIGjqwIRU0jDlfpNBOAmGXW+NH8mYcRYw8VSRJNa18+ztzElIMFNHD+pFN2
TzXgPPlCwK6e3aoZ/iaOmSNMguX9PXD0UkYH9CT4ZwiFe8p4ZHsGpxhrqUCWONdp2cRCHzKjqp2z
+ZIt9y1zLx2vDkhM/UT+HKp30tNPx3pWZhJnTrAZT6no/SfEQ0/FHNJfsxaxV2yPioqjDZzqFhhQ
J+JkafQNC+GDopxbXwBoDKvyhH5X5kZAAocNQInDamSdaSBxoixKRFdLDP6sNOkuywHeR2CU0d04
ifWnaiCo4tgIworkXGDrb9R6BvU+B5Ke07NDKVIolV+Ov3zkF91mIE5XXwE596JPYJkHgN/mgIpH
8VBUh6N4LVO7x8NgGdmSPTAgmu0FjByfNTExatZsYa+LQNGym77vEyotsBoKw3qxkq+89u+rYgTd
mkE8D/+p5VhGcuME9AIwhasISUfRXe06dEonx0RPSAnflF9E6azZgWmeCgZ7saLuGlzuItRrx+po
P69xK8cv0qm/vf7WepeduYJyJbT4UzEeCEKPqDx2bW9LPk92XDEQujI+rm/ldcWb7aJYSCzAgUED
WqmvhfVrfDrWbIwFl7g4cO4acMeGOJIda51lXQAtQaolqepxIMp3y+cMrvdKr4N4Q0gcXkj/q8Nu
TCZ/EWyULyvx3DQcRqFYkknpKEfZY+wENT3pzOPy8wjo3gZYZgp/7m1UXqNmfJoPhy0s8KQzQWL8
NPxSd+mM0/BQyfiaGb7vqKVTfIjlYGUZU8n4mtMg2QXsN0O0xLK5fOkBmZnZKF6fEoFuHASFTzlr
PbgCHx5cRbXeW3NNilsSo/OepeyID8nxlaB/GvhOAx29C7XMX32l1XsxxF1+fg6Nyip8+9/0U6d1
3BuajVDQR0W3Fr+InwoO0OOt5ikadmi85ndSECN8fXatjDa/Q0am0r6uHaYLQt8gcP0GX98RTfJ8
tPdhyFlljmyaZjLyOAaY7SWA86SVjMDl27Cl2eIJWxb1IgB9gPyDK5xFCwWBa6vPVAhJCqkPKeYd
xsbg2gpVQPJrM7VUiOBZBkC7zUBmRmKM88bm8luk0LEZDOlPx7hHSdX5d9E8SX2hmmy5SJbVkcKX
F29or4CMbFTcPDapG6zIpzeEZdlaiTVPKWLCPmirN7/YHXyBdm6+wWLnCKmUKM198rALj7bMAVcD
ru++eI7J65UY0+yVRcrU+DIENGj6yhPPix4LPdVImoE5yM3e1/BZnHod/2QsqR+JnRtOBnRlOEhj
6rwZ9bo9C62t1rZ7bbj88I7UYKXIdv6c3vtXaHdNEsp+erY/yIIKg6OmoHTkwInjNmcR3JrbMJ8+
q/03UaqZjRyGTAGHUZuJnbSp/xseVXiq2GBgYOtDViibAtPcQwXJmdSuEQ4k1W7VMlNAkSuceKRK
QfJGPr/gNa5hv77KGaqm1POhTF7CLqHJTSItcdptKYxkgS28pMRz3H899DvmeFWUgBiVGYPDkVQH
2MGh+Rua39DRK4dn6uXjYnBnlmu9yeobFqlMWq3r1Bo9SIpJZqYemIuW06jgwX9dxZ32nwQ3Nbtk
o3z04NAGlYO8KPXwiBOrTaKwBNFmkkrZhWptooYoEL2LC6HM+55Hqf9gIDC3ggy+Pg2v+NeTtGmy
RFdeanRdp5GDngTDmM9Q0NZmQAVQJCl3G5gX3QcnCMnWQf0CredSQAZsIK5S6uA+VC5ndZ0aV4dP
UAlUqDQYJJVxohnoan1IyHPshiTW0utDeiAzkj3bqdgNqmcX/3t4FK/jcivDpwHcyPGcK3Tjmpuh
EgxpFE9aYRseXJah6MQhuEI9xrBExS+r4haUvkI6BMxLVALIDfMUKSj4m6iU6sLnR14qp4umvClk
+F1sV79pOBDU3I2fhw/LzrBcxR6OGfAxyULEU5pqsemZqhlvaBoySgrnUz9HM2lM7tfVSvCo5Dcx
msQtnzSG5w+vjY4INnbLeq9AXhT1MB9pnMXUENo19uTZIl+SXJ/FI/LLv+XtReT+DRY8FukEkB8t
r1f6WiwmsV3KYSnel00aDHqNUuek93uFtXEdjpXHyFEgR/VatMkooEzKf4Lw4qJqNg4+PtKM6iPR
oeLRztQkJtvx6BW9ufAPPrQXDa4cj5rIQMyigELlVop1WA1pCCud7L7E3gpufsZZUzhjxj7ykwvS
0RqAqXRYaNAqOlphAbT+ZJ/M2abFxjhU0XhHlrlx5DgK5O6rMaNvmmcPDBZdUo+wMqlbUya6Y9Cd
RmZYg+wn/NtFU9xzDLyeXEMceNXP6RnLLdbZ50rFeUfoQ6W8mjRkHjYaL21ySMDPG5DhoQIr4FyY
v/2KjND2ikELWzcsfjRiygvBvZzmhkMfnYdPPydjGrt8OJTa/2Dtgqqyof1p/8XMTb7u9HEg2vab
TnqQ2Z9/AbsMkT1lhnSfj+6jLzeTRrd9OpuNXLL7Wh1c3HUrPzz0syqR0CIni8iYhQrO6hPRh2qA
d+iEAXRxZLLXvZxAPvOEoQ5fMGqTWG6ZItesYE0/zfDutCV5wC7oKPMIQPl3XsZiTqDQEP/5OBT/
8S6wFfU3+eWs7GPmOVTu6Wecwl40GBfif1bWZD2BfA3alUEh89i09NQbV1Xuq7u86b/fqg+CYCxH
AQCombT0fd6NWPMcYMHZZlQ5OhzjUVeSNXCYBhVbsfJDUl9htenvild+hbG4YoOjnPbtoqOClFqb
OrGg714ptj29JPUPEKR0k09ZtQCC3A6PMNTEka02Fb0MGGwBiQXOXtOqR/46yfSGdF/L1mWRHUTz
QdFFAbvaZBbPDNB0leHU+/VAvCTmXqQ66Mtpm6EaNV4fXHh6HAHHAHtFQt8vhKF/qXBdzoLC6SGX
Ah903bI7kaD/v0lBS2phZT3NB72gIhGoyx5huCFXe34nzsV/5Y7DET77D+LCWeBTJM095F+r93nE
qOiqlR2Sx0ovnUQ1W197hmRzjwjP3Edsti/jvu1uP963nJaPSKI6nPX/fjCivk/YVAw7oII3SaYT
4ftU+82mHanjE1/bBTy+N1ma32Xcjk7Xw9QNRLHnHdVXGFMmoqTkg7MFjUtISAnXynLE3dzEp/UG
Avf7NrjUASdn4ZJkYjWjbgdUk9jD6TEV58Jf7QK4SHQ8SHXVrYhQRutD1+3J8mIXljTmLd5nKbS5
lXEOkzIRwn3DiNw7Sp0FLjcLzZUbbZjn6E1S72SBPycNE/KbXAhoH45E0ZuFbFQZy8ff4tK8ZDoT
tMhIyHVt2KFwoDMcX+mKvSqama42GkGe1tw1jW0gDNfrKMf+8TZklxES7ajlaqzJaMOI2KM4oSPV
O9Q2WBu4ijgFpD9yqtpTC3v6JdhJV/f2G/xRRMUJO4qXKEiGJrqzayruLBIoe7kt9RWo/GFB0MsT
+gzWvVNRRtjBdhtIT2jrZ12IwRohi7++SDgA64r/6CFrx/92+9jboJ/Xp4jwuK0wdW+7k21DL0bO
qyKWne1rCO/iw6fBtdoBw8Nc0U7fvj3sJ0uMtYQG/2Q3V0C0U1fIV/EeX1n/8lvZZuWyP2tGo5wJ
qFabagiD9RafpD7AuEFJ+ybSPmLesY+MtyEJJCHi/EAhijHZxFF3zpsKO/DqPmld4uuAf1ZE/Cdb
RqQtEP29L8PNOdqZB7TFnzIotK3Mb/ueQ46mC0mOsltFZHNfsjUMgNdByqWb/f89GhEwwNOe98I0
r7FjYq4rjtJKtOhSoRD9EAJ1lwh659y1F8JcGEUl3crrbAVA9vC7un1EFqt/h4F5REMrggk2QDBY
1gu0vHCOEROKW3Y0N0Cr8lb5/N2xWvBNUavxVmWrh0Rc9jLbtYoIAq45FuC7IuBalBiMEgc9oSas
9CzAc4HOraxaJVQDmDtVvOnyfaT1SHZPoXfvzeX2Axso1am+u5Q3pNpcrkLmXaclQ5KxyB+GR63K
sLEEMSTsLmdx6sUjt1hr0lHXi4C4dlZ0jmx2lGZLqldaZrg4Zj0BsyscIY874pbwdwQZxq2KuY4d
lFAwMfV+j4ZSx3rGxK2nnQpPbOdS80zqepMoMZ4VyMzPmXaMiughCDmHn0PipojfOg6BPyRj3Cfv
EcHk2bzCWEUw6wsvXuCCptMutxtsMJisAsLcosNBrnGdrMBBubV+ouR+COxUd600Qi950CwhP0Q6
AwE5hXvzjeZKl+vSWV9bKmOt7rSWCeF6xw0rj7gH2rYfCpmJ3Y91oDLQZaKLq9i3FBPglDET5fBe
btvR0M6VD7QAOrmfhdcrAg2Xl7Bp2tEhjcMF5J0k/1PX+x8egD1aRkJOBGMok4PABVLXMbNMGkZ0
WKn512rU0gg74FNpUb8KWUrcAJpBzTqsqj/5Il9/l5QTTWAhDK+i6z4JH36AMTNRkpMr0ZDCUZTP
kBoBAQGd0qLQm4jZ8fTQSq+hbIBAqbx/1K4fr6uhyCe/XNSAX0bL1XlkCHp38kruDw+LKIQxlPsP
u8DCKX4dEJNWdncLhWtHPqBWBBvKRMf6FL/uk9Q0X6jtTG4OLXEHvWwN9r3acrGmAr7Q7BkcnL7M
95FUeKIDq6hYucAD8n/faWYBgPFFruVTilpfoAXWZmN357o1guke1J/vEwvGIAaaU8q9CYlubIt4
3tHxtn1Zx9Y91trXpBXWxJffjAf0OWca9Y1BkWF6afIzxJ5oFxAS+NcI2jZAdFV8qBUbddb1UG6O
q+R/saG8Fgf2WIEB5LiPKjc6ehMTh82r+9T7RrWHchkLow8F5tcqcCyU/PRQaHJWLUcRfktlzjet
3Uj1bakskJ/q3+7d941osAWwRJIeAV2aBio1EkaL1BQ1KdLCkR0exQnm87aBIKKOag1s6tYJvTB0
Icm+FJy91fhkke8jTl5RJU6fCDQFAIX+yrjuEgMfRgdCkYyzjZgIOrczH6TPPMv1SlaFFUD6FXg2
tB0jMc7z1zCbkkOxhxBhzCjt+CuKptCoNyqSr8cY4pAh+sZ+Pf4G63uGBvZ90rb+wJ5RSjkI8xSQ
Zdt1rWlNWGQhAc+wInN9m/CwCgy2VXmdCXKUC2jDSt3PM8M3CyAdJ+qXtcwQimjqt4p6U778LUTW
v3xbrM4IvSemnzy2schh2HMDYVt3b2W1JBARcQsT62GRFh0g8eZFPMi9YbD1Kymu30pCgv6GvWV7
Xr3kkAAM6dmtCiDt7STqb4Owcfg/aM5V6x/w6CtetbnHM/ppT6Sq6G7ZoZTD7Qx3rT+dKJoZlAJr
9XfpYh21yoe0UcQyDjb49czLwyEqY7UX7/kqKRsk5MroQQpjzNldShzQzEMAUSMckI1j8Hcs5C6s
GMuxqd+fwXeUnIMkAB6Fggcx2CqamI7H0QuCC6t0tUCS2Fy/GUlxKKKTtexQN3LYKO92IQhNeZYh
3g8Y8RImb8euVEmSu7gafthuPSVleR4CuMv2f71mye0dobbgQUK5eRkgFGZFrIKyno/YJewYn+5F
X19OGJI57O+gTx+PQmIgRZQ0ixBlAbuOkoYrqL94CGJfHlswExF/RPFK6aFWKybhGJIiW+DF9G+Q
mCWrgF/p1nTI0EfZmgvHL7xL0u3Ayh2TIdH4bwz/OOdulDGHmAoJAwU9STQdVVZE3rnkO2J4HrnW
CFomtSfTtiHm5ATPUDg/go7jyOPXBWpX2UcpiYCeoDV0W587BbEfTfjXaYd2Ir44pMEMcdV/xtIl
J8KzEIkpvq2h/Ssls4m2T2yB0JFPuLnpqJldmSR7zr+QFZ/EkvkzLWBMlzu7u+Gfx1vVaOEArFuJ
x2uM4WS1URfDhpQBoCItTIYXhwhqLslhU9g4RHkEBEKGaz4I/7kfvV0ybk0Uy1B4Xtw4SIa3aG5/
t5bfuXarhMeXzwso2HlLlndgG2adC2NYxSw7FOgX7z5djm0QYwWicg4k8y1evyGKrOctYLpltpKO
ZAF2Lc9iev5LXxZVOiT+9vAux6UCI7kT9CiWQ+gmc6ht1Yok8wZ4Xwu0s8ctXAYiAI/fvT7BLEvS
GELQyjgaHVoeBcfV71VhoWr5diSEb/eZQs/0AJG+qj8LZnjY6eR7VIH2gq5R1I3hXWA9TfOj1e5f
Xvlqbov99HJOK17I8wsOEz4LUOsu9a4o1P0aquJx1MKWREjpN9s+iqsyJkvp4t9GCMxpRRth8w+j
MGawNNXsqUQV3DoftWmjToYF8gVm4D/B1XOX2IOIXlu1mLI4mQ35YUq2M5SbWFHudtsWftQDbMJO
+R6cCrCsGEi7FS+3s2Gu+zEoWSNP/ml/Fh20kAzk5gcB3RAJxvLnnim2KA4+s963/NrORukVHnn8
KXTTL3O+olt45FsUMfMsAelcaxmeTFkJZkTc7+xb8u+UsfykZpFD72RQ3fK2BSzNF/fjFOCB6L1q
GNrM7etM+CRRtCHLJTOOyf7b8e91+vcgZX9z188dqs0rhQK9oCcPWCb16sz6ve8CZP1x39u6mHai
9F+aDsls0ApSxAm8QGPyI3jhErH9iozoJAstiwCSyQ1VCtH4Q21U5mkG0CQWmnNzsdMXCv/DakVu
RY16GoPrtUuWcH8nYrJUI+K1dnE1vfLZ4kh0SBogp3q6WGt5IIvTyUMyKCfMcUYbUkhNZx0+zN4J
WiO33JgjKx9pwlnQgFUzQYAsrIIh8TWQJqirza9objkoFH6ug8yCMWMZUiil/O6tEn96gd7BFZTb
nnyTUpzF34LSOkYciqvipIKY78miYX6IBxu0mMqbiwvdJ9zV/yTP/SllAMuHBIKStVmNiWNUOp+k
zBgN82SSGCLwPWp2xC+715WbBKssxZbPKIXbDXlV69sIMeoLCo78OY1ID4bawz5Qx2+iT4MdPZCO
yAdUsSsaV7nyDVImM3KsP8ameVwEOjZEJ2hzuvnJEKQ+6hrNL967F5DcGzpc1AMLTRJjM+10nK77
mujnlFda/uhcBw2OFuqf9kGjLcIys7Q+bkTaIsxGJiNvRI5FRwKNApUIMWtaQoKhambMnGaDkAR/
j1o4tsqKgcCG/rE6vhvyLhXUuTOd4YXV+Xxi63vWtw2YDd4eQufEuBelscZagpd7IjpntoH6+/Wr
1qs65tXjylt7hD69HMNueUI/N5H1dzdfOJDKIUMxgZyz3V7cmtw8kuiYxKlk5a1jrBUsumMVBGwq
D1WBWxlyWaIQ9JAY4p7JAkHN1bH/1RBm7OTTo09NsCky4fWs5YXDJomBfYRZOPTBQhl5GSDtYS4O
n9sAaG09TcfYwmTVVmt+02QVtoHlliYNYFe5GhdLo6IY5YqYrkaaO1kkR+G82hiV4sBiyDN/r5Oo
uz2F2YXtG4YAnJ6yscezAgJA0WFsp6XCpg70gcBG1NIsTiABFlYqp77lbTaqcmDw4ki9ghaLiT1M
L8wCyVDFVPZIP0w5OX+dd8zx8zcBs2N356ms7iqtqY0FkYgOyRBUrrOEnwYiAMOQiyxumXIoDw/x
Rif4FbroZ3DbjcmvcRG9+jWvq1FZsXqR2C6i1/uJIRS97GZXiA8vrTM8GCul2uHF71xuPOgzXt3v
JwO8rEcl6FCVMIKOARE9VgjrpABIhqp38P5/LWZ9cl/bnnoajgmz1YI5PqgHFgl/nE3aE5Psw3lO
Nj6lGfUt2lpPVD60yiLP0IwGTe3Yq6o7DQdMK9qL+j/Oo49f04Z0EAObtAzOQkgKA8mlUFmeBNir
T0R9/pAlW7n//YACbJENC6w9CvfQLXr+D6mQiAPmR8kLPrOB9gg2R7gsb3Ei+A+SqIYwkrArQTmM
celPrM5Gtkeh2cSpDdGJuWXqrWv0o8wGQFuKdZRIzb9qZypr31TiIiUsjhTBu8qroOIbMrYaZ9tA
ncTjCfHEcC8pyBt0dAfvWbdZjWvJp2GoD6heOdV5HqJ9bmGsa7Cml8L9JS3kfQTJ9xpm/W3heWHK
25moat+a6VXmjCSqzJDEMrPzP5wXY0pufclBAi7Dfuez4qj+2djOWAs8y8xi720yMC/GlQ9mBOly
OBwezW8+gzKWZiKq0zEHva4UsxpBPWAmOhRVDLnUaCTjrVwWNggTF3swytUQF15tjCJPTLUGHams
QYL9zuavG5qi/f0KNuea1okp7tENOP3u5CUHKfOJ9l3HvffO3AmJnfuIoenvHUNnjyahfoR22m4O
46ErmvJJG3Fezc5BJZnek7uZtBdAK8783RvAGRUSNhSdNFyYbjrD37t+yfyMMvoCWiyr+6bJQaOz
4hydyNk/edQOC4QMe6E7lwuT7xKUMqsfNfbey9splabl6xQorxqLCrWekBmDx5gBw3ljBoqsGVAq
gTzmC6oHieoXehv+k/I2se3z3LZOY1pr1Ey/bTKrFFLFpYV39cFsX1RvHw/2QgBy/LjHMNr0sbRw
uxT/mT6WVJfZTAHG1yQyCott6Q9KOkGbYw40uNXAHpL3Rt9Uip7wlte7IpMW6kvFnJ7n9d9r+w5n
OVqSSVbMJJGUqUq2atK2ms/IkU4qoXxkCW53MsHkmc5pfOmmDy09KvnYzHlNd3jX0ez1Eidn9iJC
SwqmdlP6W3eWDspPqPG7bhpSE64mAr2Ig2BFA63+HwzJHOT4puGgiRvUAitChwori4lIQ4ygtYWu
avqK3YGEgn52BGnQIhtfkQE0UU/CPTVzdVXn3H4ZN5esacoPxFYfo9AyUEDGmUIKVx+JnOCTd0Z0
7QExS3NHvEwAyYhy4yOgZLMoMCuLCVfEHyR39kvnNVKYh8p+qcVolFe00mfGo68GXz4dOaFBeb+G
yfF+dU+ZpWL+IB4zrHMF9y1c9omT3zFemHZIV97CcYEgEpTWA369WmPshBpcdEHMYppd9vK0F6DN
9exeMMHdi1qmH8tDGs3aye+U81x1QaSlNUWv6++d+S7UN0aPrC/gJs36bwEhCZNW4HXVXPix41/0
dbGuacbXIOj8DR7y+4GXPaiOVk+htiZsyygI/3JmsrCysgfexcJMAcNY8wUaSjZwc6vAZZYpe5E+
GdkqW0HpUU3m6dXF/TXrhB0YZzEcmMK6/Ud55DQVKVJgw47xIMoIj6C+XLKgNyyWYQxp8bdcqxWn
qAsX5sGNFBchGU6RPi+CGhK/qgOSP/7K78ofKsTb92b2hfq9XM8/BJ14zjDTOFDKsfLqVouFGEpj
M/nEPS44soCt9OKXixjwsEDS1N2zyY79Qw4sPzb1ZEolNn+1WG4yk6WA2g1kBgAEIES5CejkfJ18
cH+ylUaaqr8hQAvTboLOW2M1UaxcFFdskonkCSTs+OB9pat1yM/Kf/nwu5kDI8s4gLrl5isUffqt
I65qSdB0kQ4wA1w3OCSPgpwEf7brMUvhhpo7OTMv1OiW7D8+PYE4/2JnXjTAqwUjz2o/U+yWBvB+
w5wCslS6twqihnKAbNOupjQYBHt5/nqKJvC/YDPRt9rUBvKq14/0/sJUBb8tj91rzankA06qWei/
MQ/tRN4wz+6Fpf/08tykjOVu/rm1jfYOTkOHLr/uMUt26Iai7JFExRVV5z0SO8Qu5Fjqbib1ZtNy
9il2CZ4ZXK+ldSrfgNfCWDMuVZC73l5bwMGrDzaaSXIpQ2tRkaFmNCPvrtukQRvfv8JB9CUveo0b
LOs/8hMNO6sveY7pIllusCnhk0Y+HEu4MGpNXl+63Rmjyvwl+KPd5jx7Yi07IkMY5q6j/Q7T4N/l
KUmo4dZtyLR/1tdhAgxgp1Z8oNyvNisbhExGbuOi/45ILIITnKMsu0SxaGvsbj8tHesMszFcPY9X
FjlCogJBuEsf5Q5wZfh4SIyw7n685EQdiyuYryZ6FGAxhCwfYw/+k5VZ3EjYwHVp8tREarlYmGbf
xvitw/iNsmL5kZ56UH3UofVm8m/pcXxLtS8K6c9lQxXR6AQov9IyOWohlAGVPn146cCkH5g11a0l
ZWjCGWLVs+8qsWLGWV1jHpzv3gmrMVAyhPjEEuc/36zo1MjsYVSwt+QsQTi/5GDmOfbd3nAUUYFJ
+XPLIVor+FioJre5/ALsGb7g9tMwuOrgF2kvQ2HP4B5UwS9oZ0HwPILjuSS3wjN2uQeLvIvIofx7
4M0dplL8UD+M0CXvi4CvGfEZLT1YbxQULkBbsTrxy81dhpNYqSUCfZNByBsmGT/bLXMTG3ZA8PRo
i1Nsa8q0+s/ADEP9E5n6ZqFEmAXomkD6aafovLml8NmgdouQJADneYWSgyLFd+sYRCM2KUjkiTBY
wwBBCipkVZ+JDeSlgia08ppvYPUL0pJ5/LLnIP9mrY8BcJu4Ka+4AUuBKY7Y60fTVrQEG4oNBqgR
qQ88ud+ZjObbHr788SXd/tcmTpKPo7w4my4KOSCS5pDRcgEY5sPHETihzUqWVx4ECngc7Tkfqk8O
/gqirPVTWg5O4EsitLKHDjSFpKHsF34DNZpLjSZOsPAIzmNr/6/O0KFzy10O74vRZE2MhQvVonQ7
9kdTyZMP3vfzquDUxGdNTYVdNHl/2MAU4omxMiAmd8VpAtvFWZ/RpTVzvWomtnNAUo9a8774waqo
w7X4utuiz+LG7QduWfQs/r6JTDWOPKzsWKQHAY03AjEbWK5zKHGEUUKWl79jUtRuDqyqsZmNKXo7
llI4hGVlyQVOhCovneVzewLJlXjvtTtSZZuwA0ig6+s1KWV9URzvANXet+KnbeZlbTs5DipOf1zO
oM3S0FLCL8seAiXJqgI0mXP361gKNb2BacOjbyhLHDnRyOuDMFes2L7E2nyRLvJipxGAIJb9CaMR
5EjZ/G79DRCuY8nAFs+0iHftqqbhwY8qxu00nzb5iTBd3xd+S5o3nvpSvAN3EjlUd+fnF19z+Kqa
38zLf5UHaMr+Inqy9P7PVoEYolILefa5D+YN2slQoG789jrvS5g5ujJsdlA4dXsHQDj0qWcN6CB2
QaObHdpz/ZPXxA1HyoFzZKyH1eqCZPXmS4PGg18wdS1DrjwnqZyTbxmVWc/9VoS7tgSGiL6o6dCS
cWGPOvM4gDpkfuMxllW5NXtBE1B/c5hmhDD84hmYXAxfhSaM15KWkyR9apm/m56RQJZOBQaj+5uj
jtunhtZ4VinVIBojOxAJDYu0dszLn+Fs2TNdaQSlAJ0TiVfDyR2PpbGxf06Vbbk3Voqsh1/DwC9s
cDk88FyvL3W4e8YG9xQX4E+Lw/R50kMTQSajnxlHAf06T3d5jTVS3mNDxQbZql/88c6SlhN7U68z
KOy9tydQkII6BriDdawv7EHvNToW1joD1qZxnlOiY021q1TucnKJAY4OH3Fmuf1JWiAcjelOn2T1
ZrWkGKENuxfNfBW/jcZDp3RmZSRTuJqYDhOc+YNUG79KRz4lbqNZGC52nNQUPzq7+lxJ4KZx7+5/
L9Sk6dGgoLm2OIFCXcMGvzr1SKPeu+NHNcz+hCxsZgvH4hxZCO43Jccgs5702GT3VYNOkSEqXDLY
aPrdmCDcJmSoAQJYP4REtP0B1idwF3vnt44iHjj1sPETVZZdEwol0TdWwcKcUHoOO2p7GVI0HDTJ
5zkm9Rh00fc7wwVDFXdIfLi6bjHnjqZaJ6Z6mPuLhi6lT337fIu5AJYHw5qG3rtCAzRNQ6AZvhtd
O+BPMQPqxu4SEPXj96JN4WAB78zfWl3ARUG0zhPYGgLFrETCNU6B2Rl5dTsZGnKLajNCOXH0JzAG
+2fcE79XAxwbbi+V1YEpSKIyhlRL7jHov013qjfeOeSTx31556J0aUJNoLjs+giKtPEbTgUgZDHR
b8n9C0Rwgrl2TARib6tfpdXECo4ZVB7jU09Bx2CN9dYQRh+QBjmUW3lTfwHNBPBEh4YVxWf4cZy6
IMG1SLFTdjOMfEYcSVvZcUdWgR6DxmJpLxa14rjh+gKwhXoLYeP8stBUtsqDJi75znK8KesHwz1l
T5BABjI99uEcYtfeNI1pjSVlX+p/i+IIkrQs9nwSXK7wQLDuH6ieUretmx3SkNQeuoafQXNY5A0y
SrIXXr81NDm36F1ZW5QjoAvWtrGUCz664kzdOWdt2EucQ9Jhi2mSHNvTj8OUFXIOShDCZG30AeKP
wc5RBu3VUcxNyqMOCspxF5EXeUYs8b1OtmePQG5YPUDhSAqAyKUE3gRtuDbGsAY+vFJD3neZXHnJ
cDY/DtYd5iXb31ZjjA3X6mkq8c+TB/ls8QFwZi1dBBhrd7jVRG5nLY9PiuP9ztgpsESYkq3cHt39
vjXiI0RpGFFNmj9W4KySwSDv/fb3nt5gmuSE09OQvHw//67p/aOH7pVPDGPfN9keaOL9sW3YdbJ+
jWtN+gMxDwt0BGyFsoXdCqVqEBfWqhMELJMNkdvoHdRzr0qinn94NXluIDd6ilpUBfM45ypqmwNN
zejAylnIWxrpsyzBEiyCLASpuF08PZTXV3c//n93SlY+PCwVQj0iTW2EMHx6c6dtcmIXM22ivoGo
CDW0N+8uM/bwp2VP8HHduFZHWACgr4e5kfjF6ADUFvIstWPpbJYTwoyBxvnNAl7jGFLrqgVSO0eB
rXp213BXu+zGfb/M2vN8g/ewTqbFd/jlfZxEWzsiE9WSJ0UvC2NH0pVJUHOUIwbDhFSPsZE9ujiB
dcacLID94aH1DOzvqhWWqY73bWzpIO2Jb4VX5CMhgxoIU2hqdyfkEY2wxSgzK8HOtwtbvZ0+61+i
oyObgs8zYKQE1dGvRK43NDt99q02kmppatXYPIhhaQyzj38g9qu36/kAGywji6HLDWYf6l+F+Wxa
Xt81y0TyodrPqedIVS0B/Xs7EpXE3eBfatIUYA4P4QokVhsuEX/qRS5t0NHqLJv7665HMVVidmfn
25hykcpWsXGdzRGsm83Ucpy+v7/LlCyY8zLO8Xy8cl8ColEYA62qKmA8IvazQyGeDQKs0qNkQ8ZP
/6+9bm5cck5j4x3nv1ceiLGKc4z0LBiGG49W786YN8MwYLjOt1tr2S+D3kMSzZuBYmlrLS1zIpqn
81trHnKSpeewUHskpaJDogq4ofxu7hdW7VdPaEjWegdn9r1dt4WvAxx0Oay0MaX28+lGepLl9XYA
UPvWS5uSd/WTb6r47/TCrOOtpE4/kvurqBDLC1rrVpP9OK3G/vWmGR27AVeQZSkNMtCmD0kmOqXJ
9grE4ZDNhufT3Q1S4diYMaEWNOHA0n5BR8ljZEECZ10TLU3ZmPK51aO38kOVPq4TlMmuVfGJUX74
tVONUKyCCc+8tF6UhdUaBZX0lrmAre1Zm1ELlL1tJB+tupZ3akdKl1pDTdZY7jyr3e5xLn7fy0EO
iHZmfivVCjRKaRsvqqd3v1U2pSmktkTfMQchRB58kI8w3nImYVUa5A6bO83pgqCqJJ5x8iKv5OPq
gpX8bSarnfTYBQshCsvzy3tI819eXR96V1x68z5OMLKedREUpkChGQzbvS6r0Dz8OaGbMVtvLfoF
5WZDaRVXRj2YYuK13X0VR1lYnuajoaFXkNuOG1nqXZV79dEcxKy/qJbitrUa0TISreVDwwhuh93L
BJzm26lyH83b3QAPqEj3Rc8vPu9Os6mU7Ij4pQbT4XTbRfiVwQnPp0wP+nJugPCd6B4F/3KeGZBb
VzGx23TKGlKN2awCSdUN3FNfff+bo2MRUqPRM2dm69GbGzclW0aFikormGwpZAAU1JDFajB4aV2q
DCbaAQJXJSy+SfQWy2UMZTML7wSenit5WXpQDPTUVyrEiEgzaiLfbhqjJhcI9B+gM6IQEBqcHaiN
OPVIqTYHV7hI8X7H89SHHxjnb1DU/KDgCvmfNFkHg85FI9kQRe2OHM5bMdNczuOaASViZ18XQuk5
SjLJ9PPwfWvpJuILwxn0W5YF/NItftmseZrF99ncj6deoPRfRUSWAyeFYOvztWKIA7hlgtLfRGb1
Pz0iTfa8tR2brl1RwMn7pP2tfjulEji91reCPP5zjTqxTnS0Otl3BkEEXl0TaTf+OKtHS3op4odR
Xadnvsjr8YrAizI8zmbqMVFMlCZgiWKlJvt8LF/regCnnvCA+Y+Jz4UbQdXfRx5L8Xq6Ub5c0+3C
U2QIjATNHGFv133Md7WdQTejvdn//KcKgckeMciCC13vilLIO/gziNuqSWUU1Uezaro+a21njQEG
PYM8xmhi9OgHdeXgfWwTlBWwpmYLOGx4HSPPogKSsgzDsCmM3ogrdZHjr6ql7+Vlg+4k17frBS2R
7hSE2BPcdc2Szj9VABn0WsHPwtIJ7aJAGOkAgfsY4NhBetYrywcskiQoJ1mlqaBkmAdz5q/w7C5g
GOrMoRMIugT8OGarpFsMvXk+Z7qT0HTuOZgEKhL7MZyuZoTGCFlF3BLzYVolb+3Fv8SsCiRFgQc0
N4tIFbKen14ib3ZvT/AF9dJMigAQobcSZBv+/HcUjcMMNOGR8xwXS4MGiJUgg5FEShZKHDM1m9/o
djuDwro+HGzRDe/TOTrxNwaP3I4RDRTafsBJxEHq7oa9P1nOCE89Or/DRhPkxxiXzvKphDyD1+KW
TFEK8nbDQnGf1i68ZI4Y9KImNlyUTBORO744gZvcfuOXmyG301bzUWulL2y2JwD6AzLqAhS+jliG
youUpNAIrR6XMgxiHGScHQTdxRDNcbxM58yLjM0+BlzU+XCSkgM+h5L0fWnvBqrKIsQ5LSaMQ+1S
+GBBszjQpuBClEEqxJl70ynUGw07ZmVrJ7zTDd+kcfEL2ryagM38cRdRtkn6pPKWeboT3tetBRkC
wQeZpEjSVNOCN57Oa6Nr8SGG9NnvlqN4hP6vvteUsE8EvIpQFXXiW07EhztCOdV1wt6Dwe70CmDg
+x84caODPfu/qQvLZ82xuCmYf9qUvKxT+W9LzVfBTLo5hT7wUci3X9F7AzX1OQqEcSKxfLZf0ZQ+
om9to3fI7QWvfK9haIV2nuhD6b5bCSM2rXJjrwY8Uhh26ggGMC864MHeOG0YIynOFU5JfGTTr9U0
O4/kujBCRUCe9ppMH0JbgoE3235LgmG+Q6asHTus9GbaRxsOZj+0Qtz3oY1PAKIbfhN0q6uazKrJ
SQvdIyFNo/0pkfQXdEEVI9JXejtqCQ+PO1Zmrjq0TxZ8e6WeegWMz8UEfHFN+8q8nqON5u19d3TI
W1oINOff0tzU6IizGUeb9rIVris3u/UfwBqKdhUuQn2FGoyiOh17Di+G5v9y4q+F9Mmy7Q2r3j2A
crtWQIbiQLcz+/qsCmnuM7kdFR+qQ4cIw4nBsMeUMbctSaWBIkxEkId1a5gz9Ujk5yQKE85bTcRx
ht/jTFDT1ldWmM0AXQGGiWOuRIfKfrMi2+OihETiXsHZIRHrt7j3165BwplGGsK4PojJMESQrf6q
ec9FmX9NywVLInGmpPEG11nQoI9SnoqQ/C1NsJuNLGHCoNNS2rwkXsMa49hLm4Dxc+MXZDdbal17
bbzHj3UpAXfWuOwHs2bSMJWpmvZe/YKWzvMnyNmdo+rIEcJGqwk+Rf0aiVO6ytHFQK2UN1X6fRNW
Hvph8tNWXZMlXfgpeNhV/wr5Y81SznaWYrxgPt1chLY9n7+yv+V/G8GpmN4gHxkLbI9uViV714W+
gzQQxVBMJNU6j4wV46gmcAcek1k5hzCx2XwLeYH2kyJ9ls+xSzxqhM771dira6RfK4v+uxA4xOk1
XeKqTe8UZH753T8iUWYr0F5NW6sQK+Qi3wmdjrIPj5oJ2bX1Ly7YXgWEYjcVyde7EL6aT8fiLd9T
RtZpYreW2VEWk/OCEWwVIqlBAqYZblIy255c1IoDoG20wG3ZijTbI9mfBf4AqwKjBbmZeeZ7dV7m
uSgdwYGTE3HvcT0ZcQz4+psThLtpjJcvc4Xs6bloGC3DKZX9jucD5SgilvOqae3PEfuO5ALYXEvU
MUDYeySRkMK/8RgREAizisrtOaETyfz5jwpzGQhmyjdImiMum+AdFbvAo/laeGaunDm3WiObfEIn
kqgO2mIvAGAnHxEjbWbia78FzS6AQJhfqeH+DqcHrkWn6h16/xpYocf6wjwSNgZzynY0CwO6QHXj
8ZGYHecTN/FCktEtYq5IPv62l122DUrY8YDyq+lnkYqZfkhbNYA0P6b9C1IG69jWqOSRgPjSgm9U
XBwcCong/Pyl1eFozKhX2S6gGtUFl47/EDCobXwv0PBhomyGfG7t/NrEmt2Auu/ICA2uKd9V4JkL
dhy2pkyvfYSW+i0dX5qpV5643HcBEUfw6s3d/2aYJ8fpxjpdE6vjHwLSJdEHIVHPaO6gEOxEEwkk
/HSKrkBEvRsPaBWV3ep0YT+RG4MPBkdATHZIUK+JvELMr1vcDEn0KxG3AwfAfUSHO3pSpfqmuYP1
3+3mAu2IKbMT4VjxJblqXzhjzWtOgib3QQXjWsTxZwN08ftiThQUqnCGIoIwsN0UUVliUUbA17zP
SsTUgSAOV1Wabmlx/tlS8nIPa9Ndnc8UHleouxpgKOmoGdsWFKizzRrUEbGGGNmZltE5jJsYMNH5
fHgMvV0JHryV6wTgbKHOxg8OmQisD6Prr8s14OPx+CN1sU9gAqMZh1jnDta3BEnaBsRMA/qZwPtz
RqJg6NA8mRvk6GF1UX/dyOnRx5gfNs1eNiY4fLHtkevxPxbiZleXyWNfMH/IS8wV9CD30tEyF5Ks
0VsRS24OdBTPtF17OgTU3jZZ8k2ChPuaYPwPedXODiyBCmo7/H/jHd0D8DN1td/QLXNMrg9iwheE
Mw4995YYIPA+SYBDrI/VGecstT5dlH5nis1RwzBUJ2XoLOlDNG1d+/Os+tjbp6isGiQQXHOF1N98
ltjEiS63Lez4gONCEbn7EovHgJg5M4jiESBMaU7hMFMr0cJewblukWlLfagrfeR+H8vJgaiu2M+O
kA+TLllP+OrZqUcXIjNoYAf0DCTrJ5L1vr0oIn2As9NkePdqTeSTlRoLH8XG/F6MAwgeEtaOyEFF
tMpUOZltMs1c/X8u85WZAX8kNzmzjyoZ+M4c5nQeCMQYkK8i5L4507+CAfpmKbRtweUH5CTTCc2k
2NEWc4A6RgheVZ8nDEw0D0sryD+zuH79NcEUWcPHayyxZYVftSafydjfi2GbIyo4ViKRfLPtniSl
aYI67VLqXTj4OmIOHKiaUZn00FX9awUb0RE+d5bZnayKiooEBIrJ/vtCcFaSUckDVvZ9ID0jN1QM
Dq3NPCWL6wLA95BVnLo3m8WwwRw7lreX4n9v4Pcqeyn5dArdu7QqA1PtMnuWlSSP1yjMt1iyRdZr
dUdacUQiDXJdWQM3exUc9c+3/BnfwbUgUJFEAtmGE5Vfbu6IyWAXdVI8DV4z0Us20cBK/bjY9cxm
r7rwJEAa5vAqNmp5uZT9Z2uTq1gg8c9P0tuDuNZKPGruLUjXP7oiZhOk34vltfd65osJKzOd4MKc
I6ZXPBTMJZ7YIRJzNdsFLBajbIVzxd/x8NpQcRXoR/3kD6uAkGS+Z/lEtjpU1nXGJqrP+CiWJTyb
WVUcHhLOMmzyNVE1S+8KZK49l7ZopLGS4ndczcCpcmeE1M0+puGnlXeZH1aDV4XRVfel00KTLiKb
XiZ10uL8cRljMqmI/YoCCyOQRm6s3BDt4YIhEV4jqKt4UtCVjjoXX7jy3oMPO59HryOZO0KH35Ya
hWiPjOSN7AwWgwgKPENf/+R+8dk8jkC0/WxB9mEJPEVNmw/inFww06Jj2NnzL4Y0xdz2q/s3I3SZ
6iG/CbdaLwQ8zoq+gNhYN9el7yXl3/nF7dphwUEHGayNwSzRPutKFYA9ZoiRzzWqSr+03lrQS/ly
UjFiEygH5ekikio6IPFRl27AHKpzpRRyBitPndJaE7dVJPPE6FZEYvlPpBTvVI36hZcf+5/LVVQo
Qt5aQA2jfcTCKQmiPfJbm9UUDtTqSCHp+tm/WuNCyC89XWmWVFMRxPiFWyLMV1g9qptWQzl5Ocvh
3+GX9wVGDwHyQMMHbECDMnsGNoD/iDrqcFlEVYBpMNNYEhmmMzC2k9Si95TQgQxxqMByHuaTlKHH
auxmkenSzMBg5zNgWvfrR2LxQB2sKufkCaydein11DGtBiCE2nZQpGGXARpJS2YVxumq7ixHz0V4
Wh7DME7nTTsR+4sLJIBicZiXojEiByb0ivOmxpx+SQ3PM3RGXiXKOZQJ9MWLbFwco9sseB5KlBwP
tRVJeTZQ0SqFtH3tTapHi/197+64GM3G8j2knRQFX6ULP7vQ/sB8udM1n68UI/x6HkDs9VJVdWky
c9iV89OAZREWxHxT+z5N36a/Z1xoC30S5B1hf8OGSKPaStjI3aH2n7GnTavAWqydTZ73zyrYOZhK
nQ6rGvIg3zWVuwzkXBIpH+J4TNixvpdKChpdi9SkJdVvykiS+rksTEfy3UwnoV8S2eLSEL6bTfx6
rX5rnHm2xEfp7qPLrfJ5i7auIeHGPTd+llrCgzGQQwZZVgvCFQhzeiNnXo3YMxWdsBwqZoL07FVA
l5vqOhtvsNzna8XKPV77XZuk7O2KsT7YgdMqa+NwZSLMzRebpZre6Uul+W/6AcUYsNhxgUQexPA/
TNmX5vhH3z4sk+49uMmrYeysGU282HDU/5g4NnwlqiHeI4qAuu3s8W/2tVPntw2nXs3coLlTUOjr
0t5vMphbuORfMDfeqUIQYozsbopeQN21Xen6+OOIoFlboqRzxLeT/zLgG9ql473mQafX6+6BESd3
xvz1IFv1X2TP79+9UkEf8dncShgnfXp12dgA8Jevdwwbs+KwO6VqLIr0gNeYIIAlYrA/4qrIOtPL
6XCMM5WdUTKPemOQqnkLggSszWeh2X1+h3//qeNHOFwn73oCmxYhPnyaYRB1NC7j9gPAAMHOGu7w
YjPKlCogNTD9liUIrFDzgKuiC2j7VXYqrCyIEbB0Ccv/U3ws6bnQixW8Q7mMxGbSVKXDoNIoYn7F
mCIecflfJ9+y9cITi+7HY5Hdvkwm0cqeZvvD4HQaPmoKHhtGZdSbVElpEC2L7nGuiAmCEq9qaXGQ
bfOweUnG+CtaU97qB0E7Qa2HprJQEVKThhhgp6lhEgWWk4Il6WYidnzFTDu9papPQNM6sYvvlGuU
2t78swc4cqtMnOtU+ecGeFMxYaGxy85T1VUxdxsd/ZyzYEO3PG/Z+bKIs7InEJJ8+sFjksr7+q/p
nzATMXlD9a8cEqOSH6ScGjvRF8jSGaHfTEtBeXFUoITd0z2VTUh/5Hx6UyhuQYPdsFgpaqciINJ8
KQrqJEuTrwfUIMcYskWiI49i0DCbJYEJcRShu+MCfSWdCd4sO0ziooCDt40yionmHIJCz34XddBj
zGaFcLOHF8ojTay6JFDiBRxuiVmY/8de80v0k0IWsTv5YASGvbFzVxUmLudxSP6GEiWXlLhNlAh7
evUJ/Yp/iLCJutirzbXeQMSztWwTtyagvBwW5pNmgP7Czci3a/FSmedEWb0Bhou7HPUctQ+/q91e
RWxB3C3uwxVEfKqAqyM83LqouP4k4yrwBmQhSuXUoAtE7pPZFMx9MQ+O/LZpdhK4WnXfM4Sx2KKC
4HVohaK4rcCojQusAxQbdFmD1Qq7yJux2i4bGYDu2YUcbheLt0miK35kRov5sLDuQDb4msSIlvhc
MjaokfDC4zH+v0SQpVSU2/qIvfs+t2ijZgNkfoo3GFjRZ7/Tlm+G5QF++vyUrSAP8XqPwbMBJX5E
GqtMGRqm3ug0yNpGqZTLPwgQnaXDx8EZ8wLfKMO4DlTKtQzeReCe17nhFeeD5GAdlAPwxGTG8m3I
aOyNVizrKomJ17x80B6ZMcVVtrDRjTPPUMiN1Q0/Lcni2R7SAP9eNF0VlREAfgVCpMm2vNsgZJ5N
JDUVXKAZuYVa12QgC+W+7dRNmMUCzRFUg+YWaxya7GmG4d2mTQ+PcjD1LD7NCI+AFTwHBLm35nJY
Q4zItAF9TnGLqqtUaYNEa3R80ALTFgddYv4ZmZRLky7J8XrxhCIWCmHXtLp9cI+lKn0n0YdzgKVP
e6dexkM4iKSMZCXZQxerXkcQ20SEsU1vn9cDHNy5hmGVyIslC1qPJitO9PHUWriNcPjSS1DpaGgj
vSxtYR2Kkeg8F60PLpRQGdys368dW3G0OaT9vz5tnbcW5jZWh4DeHo+wwK7cbMPxowAUfHydLOST
43t2nGtdWkIrPENtWqVnSZGd3+NrhOCkW3s4G+m8RREx/j3Web5nBTthlO5lo18CJRmfsKQpAP9F
lHpVS62ESIDNHRwoDlP0UVOpRiTN6aCypx8WI0O7kJs3UAPvj2pjVbaZejCvMlWVV6ejNc5W/2q/
nApN5PTQhCaPbXuputAFNRXJuwG4CmALPhUGzeJAo/cxsY6xQzA9eje95oVGqKoW8Xo/SDO3ZFkd
jDK8o+8kLmD6UkZIS0NtT9lUymis0RUJoy1PLK7MNzesXMGySsPccYOSAkQj02ZuuN9QYLahsxhU
kxNAZ07/q3qTpDy0M4ORr7Y67FfCsqimO1XR3e/iVZthmX3+fQlZu9TeFbBVV6/3JIPj+eIrLZtc
m+Y/WJh6yKAaGMOiYsVPkHBiTBEJFC0IZZ4EMmwQ8ll8frjv1WFCBaHPq336ATalNLAAcy5eqk7C
pkmGrtAq+OqztapIquLXfWkcJCH14Ys7mC/WPDVOUJP92Arq52s47b6HU7LXDfxWMGuqYHPzGasr
3aqvA2ZQvFC8HZF7yH/NnyELkCAgYa40pSP1R/h/HjBQaEoX6UuHKNnzKP7BWupFsa56CdGbsdag
yT/9efdgL1HEhwWueF9vkC96K7ZzlEv4gJxaKNWwl81x+5V1AIf+UY8ADd0oB5p//XM3+c6iAj3C
b+pqT7FNg7USJaVZqdGtRR052ncZajpmEAbIFACLPbaewurPa9sXaxovn/IG0uOJtZOoKdf+ylB6
jY048BA6WX2qAQCp88FfDh5Zgm1qqVSGPsn6zcRLr58jO6beeScaIQUZfbR24yTdjY7tJ5JoLS+n
JdVJl056RWX1ndb+FvkoAHvzMnO9xzDjFmuupRs+rV1Ozgp1e8BVIzsDVQYoZ8X8Th193h+VDFpP
ce3ZhH6MVSLvl+KMFaleuQnS279mbiWdIYrr8L/viXCrIcyiTAqn1bJQVwKsb5FUpm71b73iclX1
juLA3zX0u782aV0EUKBBaG53BmKlG9Qao9Xoxd/x3qzZ6VCXXGQGifQIwS+7p1XsE+l56kOAivp2
q8LRLU+Q/QJouic/h+nnMKi3QYQrG5chsHYCc889oZkNjW5jaHXYtZDcPQ2O482LKvYgUZinqYHr
JyPKs1VF/IDWZJozfSq3MorJ5ZR5OJq3YBt+Td2GNYaqkYBRIQqyT2VeZ4p/MMWrvu4t1eofc4lO
exxU+H6S5osNiXqK80A1OmznggCasOpiJ5iQ2o2C/USTZGLdxU6UCWZenOAgHJOXD+wA4JT3jCty
wci+j+pb82nFrx4qwz9As1zOAFgBIQpOpoOQzhEuNL0aYlG+ko7WCUTPv0BJp+KsIT9IQiNTDgLd
ABu9XBB9GRHzc/mZ6iHKcoLkC84AqeYmsiQ8UHi9oD8EyP7LgWXIvETaW0rbkMq0JokLLrDmACgE
0K/ropZ5H0Y9U8W+j5G2c+bu86ih6wwx+oEmcwsdzkDwzEyaXCDP7r6R9SWWGpB9VbPPG20HckkH
HGrosXvtS6q6moX/VHkBcrijj3AMcGKPhx9Z6YEepjKGaWWgg4xYJ4Ktbys0unoSLD17IH/SXodf
+cFodXQfy8P9olRCoHszLNnWMT+ZdFyna4G+BeOCBDqybXMVEcy1zybIjhvuYYj9OOrgwpsk1WKD
OS8m+7PIPvuo6TMPMA2/S5KSxFVfIyTBTcZ2YTPEatBViwp6V0zsDfEbaYOe3kpSJ0gAkc2YrNGu
gBrwqeb4DHjv3xUlp6VX0RGLo3K9nv0CH2qMs0elB/k21b7zfWiHDaktUhGytYCIXIbLxJ8QawyM
stss1odGS6kkXRVaM/X7/+Rq0niI8KQ/A6Cji5QINdTlzCat2v5IkzUnjBzywOA6QnNW/4QBYl6S
G02F2+sXCoFhW/AGSbW8/9HaaY3XABJL4ER7AiHvF6ZBp83sztfErDlv9GYxyQbnMqbPZhcDOVss
RSeA7lH5RkBVdzGO2AZnCDM9aWEK+W2QjTrlU1uAVmuT83ZsiwLgs+RpHewxtOXJ5h0iZum5HGv+
0ZedETZ0hNBCNIzyEXxC0HjUg82hcEzNsLvxBrT5Zo2KiCekqzO76uTZcjlsDm7XBHguZPhqogOq
nQMGeswjiZI2+y1K+PSHBRd62kYdnGGAWKLl3SVvUycLrahpVYW2m6uK1vAM3Jq/hRvnCJFO+okr
Kekd1ARredv3MZhgIjbYCUdEVcSYY5fqCvq11psJrAcql7xtXnWTh2LHozg1ET3m8n7sglq9Hvue
Ag5UMCsW3C1X2+44aa+9zM7nLVauSejda0AdJERQvlQ1keab6UCj3mI+pvtdX0iPnGbO0BND4hNQ
YD4pAqkxPrkWWxbrQDPEJxdujRNUMifA9r1IO3LM6UlSwAOjEmVb6FljDslOuh7Z3xCrwoNbiPXc
CUdlyq/HBKrNTX2PyAIX5Q65IIPfVcwWZzkgPSgGJQlff3Z3cwgyu+N+PQYT00tvXKkgrEnvdKrQ
oJzAMRPIx+zDG0Mdpt2qRY9T7gJUjMVZrYtcHzEwzyCfSEnFzHyh/HJjHv+MjMLnqErXj513bMJB
Qv3T+0qvYcDwLkykTh4HMnTwXmpP/NuJXgNGhZcBeOfbs0P8f2NiyD1w4qdeYhDOMSo/Ei1bKdZ/
djBHCN6vUbBa8JoMDOcENRCWIDqFDdfjtFPdBMsYH+vOLVPMbDc0tL3LnQF7RvWIzrMFDEWCe6Ik
GtsH29O6TYJ5guOAcR2unQHhoC/PZILsnAv9yciZwvNtovK00FTGi6UZIup2ZPADuvVUDugZucbn
x371GePJk/k72DJx+ah+Dg3F/Y2ImmUr9L3KsDtXwUS9TlJlYxf+ReXxbdfy3cbym6V8o2053gWr
O8eIBph7cGs2NEuavoPbebkiBtMBU9XR3hYk/PyaZDQqqbFeYGXIQ47KXG69wMc6v59v0fSuCY6n
m1XWXGflbyOQIz9n022ICFCuCV3KOG54LSZ/vgnk5DwHCWT24k9mDreCXIW0i+U6OHPH+A9A0DWw
T5MIexkH3scjFQB85fBiRdyTwsSWUsXdiK5thV053/YYs87fJTYiqVZ/yseQEeP71auQdKHRfHpJ
ZtoyILq5j9YI2hVtXeRM/5uVhYxRclJS075xoas5voicQuHEjWQayDsKby68A7zPbtYocRfmVuZA
93CyYvicCgfhq90t/stl98LY49/WIrj/Hr3esCrN8H51XeNxv2aQOtt6HKPjwf50ZvWoUf4isWSR
g+XILU1bFF0Rb4r9Tu933QYmt6gH6mKkhjuVBWvuFvRwjrTgBIePNkNydNNyUJIjLAFQUIzToQXl
/ELw2/PYlVQZFCiffofmy5BOUm6R7tJJhudBLOxQxHHHW125MYYzr/bcJNIS8DvT1nTHvceH3oPv
pVsPQH+w5nKCdSJk80QeAFin6HXNjnxWSMeFYJq6iTM5lzHTzvIKpGbbWPvvA/tBOPjHLz4gw/h5
uBG5W2pyFjPMI6RaSqvX3FJ2Qbm19687qrOm/e5mtgPo5crQpd3lwvmg0VCa+sWVn7yCQJL03Pii
kbCq/BLJ8qRaDwXL9B0kFAQPE/kV3r8MZTAvfcjQpG0KegQ4qHbZcY4rAieg3YKNtv7nRAiwYk04
10l+HzHOcFLsgqRJXmm9MnX3xEPvJVjVG6e/osljm8DB/hUVqI7rvw9DetiWiyNPXOXm6T8Ghjwc
Arh5j5kPjQ2zlUbo3GdXQQJ281AjduQnSgfvlQMpSNKNcoRoKB/yfqac40mTlUI4HlQBjtUsXRCb
m+MhzJbyTQTvs3aHKtnnHZ47sh88wPN+6U2SzCIZvqNn9B7HSC36MA3ACxeiFt+GkOOgp3Kg9orh
DI2CmPC9xPvit1pRF8gCWhJhh+IcUf3xlQ08oi877UlxQ06FgQXyiCIRhyfuSG7cYigS6VBLgTdQ
270dOj5qbT1lDE0xdzkSQcxSNqmJPhmATzkEDfbdRSUQ2ULksJygdIAfQ52xkj9NBz4PMQur04RJ
KgYLapXqakhEszJAXL4d/ZuCTyqBea8bg1QafpjlI7soywODs2aaaeIiZmQSmbZCWPPjrr3ydqz6
nVqmMFu4xTwrtviCae+Ndq5O1BFW5WF+SxGxPkZfgeP9ql1C2y6Kftm2QCCyMIb4NvqxMud5mpXW
g/2R2rH3t0MFYeW3tpp3jogGHGE8oCk2jqotTl3Ca0HCrKtPdcoLmmV2VMrs15F5iZ2wX0s3dXaM
FmnjBxnZgDqpJ6OAZWTMW+vThs5dFOpLczRpyI94+Tm1AoCcpHvNuxg1fxz7ynoZ5kf/DWF/hKdf
ZMOpewGeEJWFgwPqjYpLoRy6niy7cqyp+09trQfAxu2Xf3x8DYf2j9Hgk6Ys8jyPS+0AIfFRUBHi
hC9M7nq0F145Upbo5oImAF9wisvmnudPFqmWWNNjlcUt3WHIjTRH5Vre80dZTzTbn6mloVFW5Wiv
1aNANgWH3rPujW4RJ23Oj1dAeoqf9EZ3CfPpixDQC3FuHnEPanbnQsDQjGfbO76kn5wT26WgJt9Y
4WRoUzbu36+N9BjoHBcvzKY9JSToXj1RQ0T1aobVuYJR053ump+u6gVixZ9MbH8ngs4MQxkXMnvM
g05Gkqkm19U8PGFT35+edRoUsTo8E4pgGuWsOagij+YVZ32Bu2W8eHYvXfE7GnZvuNb9yCn19Ll9
FYIbzUhlM/b6demlWk3iM+izbGP/4GaxmmpXaYUFYewANEMczLFfafI1+I3Ld401a7MuF6yrjX4H
Sx0gnjyRDkDAxBdlToAk8I/Madhp1XtjxxFXsRAWVuornJ7R7tPSY4NNGC8bM3RndXE/MTmls/h7
vTxJMCnIwAskEd9ZS/6xClVGueSltht27KBcgeVHmFOIlXHgwgbUZ0zHZ4sZFhjaTE01X10yWTkW
CTRbpgv/vSP6tYtZXY55lqYjtpxJxiG7eiE8neQ2MKMjhtDN0RQKWnZR16UgOWN8kYSqZQty0Cts
XDFiAd7JeIbdIngRkVDN5jGm7QjSpUmMJL4oFMqlWA2MlcwQKrZF323v9eGEvJ9OsihJVrxprDDA
JIZKFs6V1WvSlPE92xo0202JEqScIraFtBTaX0hTghhHgxdjEiMbIseV9M147qj305UqSjRkXvIo
z9BuLT6kRg506toFMz2fqQppP0NzIwCo78/Nl4opkLECsdzm5veZ9SuNF6k90qglc1IoZciBn10v
46Lzsc0UNbZYPusOUjONYSLEzVr3PDyOy6z7kJP1q2qWZ8s2ScQZYTgqHVhXNngBSi+szgZCUY7V
GUS4F9uoAKUpTTFqEWzhO3JPbdMpCGHpQoTVxY4a27m0PmHlpEzKba/SzC2iPvpweqfMKQQplLdz
r70K/EDF8GxwQt97N2ELFfpD7Lu78Y+h/RXUcy0ljVxxJGZn8DFXjHeKeFXfNJnAMZmj9OgtfW9X
jAvSXirUF628IiWa6GkIpf7xHv3hAlBx9e2udQJyBy+J8NLIC2Pb7y8IdrdGyMDNm+Ir6Qc9cFhD
qrKAzYTEpLYoXssTBPbB4IhdRANTXvFo/lPwMVp/FYREXVxBTLU5gdXP/XX5Wnh7XknRo9uuERbV
kaDgfhOJAjv8KpPKflby5otYZMyt49WLF7+fxSmR4iHAzCjwDAoF6vMfoJKS51U6tnsUegjW33To
Fwi4tkZXeGLiH3amx4jbEMSBPyUte+uEPTbTtQyLmscB2pjAKZE/YY7GU1pbSufIjRTIYPyUPM8c
OtVEZwOIQtRi1OZM+jhU9VdBZT1ahu3WhTYvTO4OjOQwjMf72qQI5Sulyy5Fh80aysbwxFnkQD7l
lwsuiMf0Vd3Z2vd/VZTA5DToIK0tUFPoXSot6jBXjyY92f3ETP3CWfw0cErcl7y8hl4GkPERmO5G
d0uPgbv12Pu+2WvpoyOgjnmO98sjdWv9HddCu/eLyXW2l77Tr3Up3f6n6qz4co2FhDw+68C09Ag5
X/FVa8FNvsPBfLXvf996hriRMBtYCXl/BkIUGG1nyFqEd+JsXmg4QJFYuoQfGB1YgA15v4EwTUUt
aI8/Kl5kPXakv5fwGuQsHo8ZN9SbPk8AbRtkXawQO0i7/l4VUVvx8dWzSraGFvFYGTG6UV7qWp9+
BenWUABi4ncjDrK+9/ZtAImNfwl1qTYrW5KG0zgibTfTv63ZbV2khPGndODU1vFoeKm+2LBTxzpd
G6eDyh+yRYXU1d4COiPKixwUOR0vH8Vb3f05Z3PjRJAxeme/nDXSjjsOwR5I1lDUfIsmfyk1dIty
VyRZHVPzucIsFQdLJRVqutDOqFAabuUWUIPE0WcxCH988cZgOUTcPgL6hlYktyIcbJ+vflb8eFpr
T1eCVzhdlf7hqPeUVaqAtXZ/HtReIF9JZQf/GdtMirqd68trWPaUb62vj2hwSuMxvg8dY7y46/5V
pw6h+DHVzEWrpQxi2qSfpjVQooCG4SubCiblhCC5p0Xte9fG1Hv/HRPu7RwqtGezf1ms3vE72EKO
0cVVxO41mq0TJIkgEz2bXBt7fogjbHCWuc7zBHsd6DiD3L47xVOo59iHDacsdMP0u/9EPU4badlb
u2tONnzc241HIaNu5oBjO8pVMrAMkgYxDUJf1zhZeTEKPGoehT+9hRTTX9va4C+Ktw7O3JTQ93IZ
Vn7dRN6nHa4wSCiqo8fxJMDwnJH27V6K9OZs1zpZkdwkZWLK/4FD+2+qiK6n/usUNW1ZGSJtb+qH
lc5dCvFBt7AREctsS+pU7pBtWkUTJDqw0KuHgi6Gr6jDV/+vLKqP5I8QLFXmiPt3URF/WiNeG+lg
cWScJ8K9poc5zViCfcVubKCRjWYxXLOc3+sRjp7T/q0+kQu4W66+8D4GESxxKOkiwVturtaCKBLB
Fr9ba3TiW/EYLNRq8vEBeD9rO1ChYf5m5vGKkEBFPVp4iPmq7jenHxxuIGBjYeyarIti1WPmI2oT
aWVH9+hHCjEGRL2LJTZIwP/sXLgVD30IUCuXNHkbd5opCwlQs+ZEKMlb32P3YPKYytDHKYLpvy44
iX0dZBo8e6miC7ole6pNXg9z4GSKrTVZ+t04doD5eV7lGE/CW6tpF8oMhXvlBPk4mRaWPjTSy3Ts
zLo3HsK3QTRs4ii+Mdgyp3uvmaopMEHvtK7bSo/xGdnTqFoc+GwLUNWTsuFvPxBxCjPgGXMp12Um
JYVkjZJq+RD1RfpS33KN3nf+tRVeILGe2IPjzbl6Nz5U1d/s9R8YHTzS219pwFAyWvcQJHwIPO5g
vcnj1b93zeF9w39Q+iUfQEWvb50rHhn85aoGBy/KRaEa1MgYumZm11Unvly70cXqaoOK6psN8TAE
ctNsn0UgWYWl9gkOiwuaFNEQ5urA3kBVdsMHfKjzRb6xKb6gsiFnQEeFFNdgMEufH//a0RtzA33S
kppOMyTWJ/J8QEqljOatvvGEuhHr3JFyDKTtexLNNR+Cu9sO6IFUIMW7R3z3Co7VYEcgX7SDM8yU
O9O5trs4hf5zpnzSHZxh88VD4bHdgC5d3eNOrGNaDCuvbYT0lVCW0bvY1yvf08g6Sr50BUJ9ucic
MXFLFxSQvyDl5iHP8XX0PPZxhz0/1x9DL4WegHse6aUQ+fg5mfkMgQJu5sfIo3ml/EJyeMNlXaPK
UENUXIo6F/CyUTYXdkgdXbimE+G9+I5UvrwB31KfY6wDUlpXoJ9+gOHQjoIaxC8EPnsc2LEJ1zsg
2C1Wu6mhK4AhwJjcTptCb/mOxVfdANSdwb55osRlMzHOAL3icAY9RE6fBRwdgy9UAahLXY/yxJrH
Y3GKcFi8a61aYkQqUsgAT6V6PvKfTFvf9hKeY0YHThOHfhJgFzbzpOgxKEjMA3zZKMucKXoWpCkC
akt/7MSF1VLTfU1C/XepmNMFuZCkgEm8+ykOEP5d4p8hZOEJNepnpI+ACUG4MSiRJ8s1cK62SH1Y
a4Y9d0MjRxz+ND2yLe9CL8SoY/i3lg9Vfdr8U9X1Ui+wtarYVZeH+UmmxUtRfWAlujRodkXJaBss
Ep139osEIEfGPE5vnt4HJVwrmPVywVIgM1cjvdxWrdZOH11ybPpXxrWoDvOv1Zo//BuiyQdZqiVN
65MCWWEDFk6C6KFJLEMswLcnTpnWizxTddVyokPQjbZzHekavCovi12MHrwsHAzfcs7J1SLHDDj+
7zrxlmfIStDR0zFXOWFmUDZur+nZ5G/xHt1MKSu1HecXgTj5f8hxvqU/0IUmBHVoGLHulaInuaTR
pAvyafdmbiwhC5dGgH+HdAqAjhw8Xq4KSFRogKD8zCu5PC8qXU1+IxKwIEuJVowJ1R6eH1gyqLz2
O050Ib4zE995bZ1iX7iY9wfmk9jq6ClUAVpbJnodFWqVIio2RN/6kBGhYtWnCz5ridTSWViWJHw0
UL41wGedG05y8hy1exe2D56rLiq08DrNJIpCpPf7J+U/Mf06yMC2deE+SKdIEmTAdKHd+R1OLoio
kYWyf7KbiHxSEdn7lu8uMQ3c+nLEZzD4Z6gUK0x6+jGyBAZdLHLNtnCPdP3cdAllAoDJ+T8tE2CM
jTqb7RTkC0doX0bLMQnOCpWNz5+KZRxpzRCvkJ7osVkWm9BnI1eMlg7JkLOoUifWeZIGXeRJTTza
8h00rWPltnqrhjggo/qVM4rniAFE0hpNAHV86R4cpFssVouCDJ8CnJxOXjbklSjyJcW4++ArFy3t
wBlMQnL4av806ljT3eaVlsI4robgCE0DmmKlHQhSmyx3fNcXGIUwLP9GsvLs7IUR+/z5pihlsi/F
2/2TVolenOcYgLvoK5yIg31jO2KP5LIO9LrPFBEKOvzwWI1jOhSPI1C1xJil3CQEf7CnyB53qVfO
cZRqfWPYUwv1tklqzfDK+Sxh2RO4vOiqkQFordq+jrxs4/AvFXWIpByFmERCEssfTDrRL31xPA0G
m6wmWB+10V69VHyVxGAALn34Gtia2yguI41q3Eo5wf0ITZQQ6ZUCA8Yih7AGBhmCoOD+JRj1HAb5
WIQLeZPhkuVeENlfGuC7pofXsACG9L94lIHGmYjCwgRJzi/3l1XTBwqoOnww0Tc6PDvul2wwmgu7
jzH/WzjYCB2t0O32YNbgeb2TlSFo0g+SsecvEaLnImuVdTKLzAerv2KRcxBo17HYf/tOwG3PTncc
5xjT7eS3Avyq07j9NEnWb30X99IhRM6b792dwFFnj/I0n2q+XyueF1DvGEkFWHclrZK+KEp3Awbv
gz8Q86+0+Y5MKFElMKAj96C3rLLGtYKdeAOue4qA8tcphHOE1XnXbHz8M1IAKbVdsUPctBRF4SEM
Qo1+vDyds/Mxtix8EOGN7GSEtUXiyh+XX0IXdjr1I1arZtAs2LGgWM2EcYMeaLEZSJzTY5vInHDN
Pl8UGEOYWBYu020AqQCsvJgsQXYx34N8BskeuYUoO3/T4hxOKx2KpQd9iC6q0YPOP1Rki9KmVqfl
p+p8PKwX1nMFvnMKg5YbB1C49zv8aVFQhq556IfaYeRrBsolEakzdMp9LV8G3RCq6k0JLiiznpxb
BqTojAAYljKOzaAsH3fgNNiXj3O8V2pnn4mrlRWeivn042O+dB2fS8EtU5IQjBYi5Ojap9yLkaSp
+wuW9tjJMxkyt74K0ddzhbyxsKOPhteTOp0OV+dlJRJp5/wjmqGVM/QcIq89CpADTDWsvGB3g8Qj
dFCrHm/URM7VCiBJ4N+P+uJlppdpFXhfxKI6J3JgNFwxOJJqcP+ko6tkMkrpyfzt2giRdLKdKsTP
j5kwIKzQAITTl2oH0t4bxO3iMTFyEDASXsFJkrwUsSb3SAy/nREkbqAtSHygYDbIM8lKyaABBU5W
pIGoDpRQyBEUZLxBpDDUlkloV1SsV6YYsaR2lpjHOhSDCxpsu1D8KtfXONC8IQUIjsHGz/co9Fkq
+RkDFWjEi8jUggR4+QYzUAKoNnVlxnPClrq3UOsA8ttL5omiIJRo27vBicAVHuZWYn+f1TTgxjSt
k/L0lgbvRBLHJTQ61iJLbsADY4HAdg2KDOVCSU9+cM7qdwEPCjZSYhnMDkqjVPaRj2fwduuerkI8
qn7P/ZLpQq1E8FnW+eYVH7ONJB20SnM7l0A7GsFzfYYuP+cVeRUB3QU1kUbRar1oSJaNmMCSKIaz
MdiRfBMs6NdL6t+AdAeqWxGRVmKdnSEGLf3vybZBjdZjv9arszRFM7GUHLY/q3JfaQyrmlLR59lk
GUmscLjhaBql6RQPnVlMzagOXhsC2F/fIcSy+dQtfDw9YRM+I5TPKVx2qS7pHZQDMzbRw/9kKEeo
DxOuWQkwyF+QxkgLbKdnyZRlPHJJpjXYlmIxgx3x4BE+pWuMR84gdP5y4U6x7R3WkEgIZ+KlCE1H
snoJguH91lbJGcYK6xrsdpszkUkbQSrSCRd+gHyeWDo8BtGluzEoXg0678jvj/koTs1u/Vy1oAgM
QRb0EfJRpeSR8HOls7paouYHJxgqYm+a0NnVy/cHLrixbYKwGfmhatnum8vfDOozKI2Pv+qHqt3Y
mur70Ea11gEyCOg3a2ZolRmKyeZJdMbHZZ9iRA8XGEcEohVw1ndNXHlOzNzq0Ku88uS8xaa31aJX
p1FX6AAUtH33LEhIh7ycPfZyzpCADmmM2ZTWA8ma1albytP5VMCYFNgoTwuizbQVEF/VNPTEAr0X
7JLSuPQ52TMxdr1ZS2m+SxnqiQk211nXBlmjNr62xSjunA5AaCcmPyfa2WAgpS6ry99j2OfxQqSY
x+DvkpVnWZoXDkGV+s5+7cchs/9VPQeb6vZeet7m/vXlU7c5ToBY4gbqlrS4EeIbODMSwu0s7EAC
pHBsjaCyv2eKXwnyLFyV2UdLXHNbB9y553vvjDEUOvQpDIEDKFeUKoy3dEmsa0IWOAiM7hqaLzj0
8dVD8clUxXk2hdtXuo+CXo4TQksUjeJkQCn0EPWxhfzB7A1jlCHxcU9Ceb+2F/hDdF88pmMaQWsT
TUoki97B3+BeTDX0PnyhTrlAZEmfHqHADqpY67y5lX5GJ11Sxm2Fao9K9OtL9M2dxBtdGoxJDglH
P3zXCDUAbf3ezqA+gVkXlup8MmcgmsJR63A+0az9bSC+TMmSpN+u0+cVPHrRAmkPL1nuJjp+kBnK
l014Z+VOc9gpN6wRdTDz5eXeZlgBntjose3GFgNv31P/hE/Zf6UDXAs9IfUJSl6CilLcduc2weKB
B8pdFJ+/bxiyudq0lf7MXW7QuIGSjGtBBzwKFAqpFqszIBCDXPQ/7nbLeU7FXI/GzW6bxQDUdoF0
JeD4wuWLR8v42gEjfu3WDXTMFwcMsaqabfdBzA9/n83JtL0OQ3pftLIrdccN5FIO3CHN4WEmIIp+
9/IHRyZCI49J8DFiNcELP4JL+8GeQJoYOI7FxbAtXkx3DMSe8/L+7E93QPVp7GxsTFGL0R7WrIRi
rPj2B6D8H7CNm56P6Dx9HM8KxomHNuGMO7x7tlamknLEaIOQ3I9z7aMTqqKMVLeLlsVG6JL7Cdlq
LpWOo++Y/gMmaVZC6OOYJdxdfqVRhqQKgGRIp1kkwWGOAi6ivUwBChHpB7oCPHtQOsBiLzhlCoG3
KEPigf2BVNRCB/ffIp9qqHoLbtSCZLr7kcpi7j0ew9lNxv5abSx6CKdKxrw9qxTLPZKZ9/VPhoJC
JaOEvZBWi4GG4V6njkKswokeiv1ctYCHiTQ8qd3b8OcPhaFKC99DpPyqQ1w8nbYXUOyPGJ0mVIKT
eVnG+a4ueCo0n6vEMga0dtP8GhBudesB03leU384wdgXkWtZAs45PmQcL9eTbX5bbFk8rc97j4SZ
AgXezsmJvDBVRWL7xbHTnf+HErTRqXmqCk2FiNJCjffm/wkAizzSgZXwvW0qdCZUvzbZv87iV8Dx
jYRh+/fteSOBlayeDLN/JnJRN9xmjSApZZJCL6sYDC05fKsym9JEbFTy7eiTJiZWvkhCX4cpvEvm
EhPZUgzd0LDhUrYxI6Lu+FVo/vfOIZAcjM6qU9bZ6dOtWVAru+5/dq73l0cryW8pEuo3KIzMwEU2
PeEryjhe965MaLaUahO/J/BfKtDO5asvrWRvNvJtRXNZhR2/QbIA1VMcj6en4sMIjRRfLZ7kkT2y
q4GW4m+8KWIrV2C2gPl8vZK2LTgpofpi030RfSU7f+nj8iV+NpSln/CMwNBpUfjgtgDXCK7LMP8Z
HgLEBpCeYmUVUUVTKhlBkVrC2r8S5aFNdS5Hnbrt68poGbHIlrC43yr+45R675KmvnJ05Mt8+MIW
JmawpPZnQJaC3CAGpvWfIAQJeWbSPpHRbsHFx1T7RoD9EBTjiyszUhd+Pa6TP0KFFXJrw4Pya2Hh
r1M0uSH+hygv84hzat63PAcorTjcZJ7aJ4ySPcB7mERFznLQtALd06c3FDL/mkGLpqAo4cQnZLSR
kH0vTHZopcl2AI5pIRdTJtIuZvtwRT0P8VzNA8sG+gXiiUeXZKWZepvSG4xcHifPCgm7TaFS65Ja
GYLMVVS3iOQhONoxukb1POqYAoglQUW0Xa3Dzg6OqmNQBD8SdgV6jiz/OX0CQyAF3wBxS3m+y7S+
YgaCdwVA1IiP07XbH3AI1LjPVMzZ/qt2Swr4Mb9pJOHNVoPQ4a7V3MrYJYk5ksHoB5XVHHD9zkJ1
zZJGvbIrjJm+czLiGKReU57vLYqL9D2+QtLM7fvUiMQVZtxmkfGEyZ2nKXrVWAbhle2G1subWf6u
bShJNFH8AwPAHUcwN26YRt+qaCJSIY6Taa9K/xraNZkPtqBihj0OO3HtdcbtLpMt8s8Eaag8bj7Y
FY9RuARo7+qF+ZBxj9evy6l8QKGF6zsTM4mVgxQ6BzZCPEnaGDAIj6YNsJ3vNkc52Ils5cQahSEK
N7ZMx68t7mzeRkfbfZIZQ/f7pO02W+ptJclzsnrBOmx7o8jpm7qzS3hf8cjjJxWrymbtb+hriFY+
2J5LAEt+JyJ2XE5+8gI5jyc2k5LBZxW9XwmLZBL9UPXXq/ofFaWPyHe4/su3aoVq/NHil9UuA4WJ
pQVFb5oXKNJPjo42G5AgmltdvW0j1van8KDcbIrGO4Hm/qjFct6x+GMoTAsTO1CYgixMujvOSgTp
iCNDoxWL4W45xTGvygPTQMFk2vlVdxLKrSmDm6BJheBYPBMnbO2bQ2qYsrC1E+PoyxYY038zpk6a
phVm/ZG1Ui0JACqgp2plvekYugk4fW3EPUVMpjZ5jXqOKqb0663jcx9es1KdW+fx1fXh8FkcZBF8
9S8CuYeWy57LOPDme7IffOAX2tDy33gY8OCb/i9N+cDpFt5R7mwXoKGsLRE0IwRsyPdvVOVqpN6G
Js07oAVvkI4whuuLAHH1e1kT/mXOmpEeDnmJ+eu7/bVFaud220RchZ2F3br0sdYLCms+LmQk2nMC
sAY8XLvKQR82oK4QMJWQdap9m0/G8x+3KnTuTbDLXaKO6++dGmGhGD4aUGjGMsDgFE2nady5X2qU
3xRMpPy6uapQRIAtNgyNhAkgejd3krikhX/TOqby301q4MzWTZsWrpAoskPP7sgb+Xypy9F8l3fO
oPd4w77k14hXxYREvPeSWrN7U5L+6waMGArACCnMIzGcAoBf5u+2eiNsJ5ZWSLUn86moSd9+XA5j
aD3A/BijnR0qXiLHAhgyuKChbl60UKCGtoinoNZ4GhuHWZwb6eKU5HIH8uqn2/Yk8BfBtrYVHhF/
DkgHVTuDEiT1/SeLkVqjQL+tZqeox1OW4aZYEX1hRNsrF0siLEoJOxRF1rpoBvUkKSfiI3OtdCFc
WNgJ5RFY7JXKpNkKvoGooEhD79r4Lmi/g8zMMkUurHH/oTtLhb4gYPuW/f3umLpcd6FijtBHDCQj
4PhqF8pTxz3o6ljdC415ZOnbRJzoCbW2p9i8+4/NIwHcNm9wNj4CvvXIwTU8bOYmRX9XJSMyNAjK
aUdZMe89XNmzF9tGXl0CpMdK3hcBDQKm1aIPGOyvz2UO5bocZ/LVJVHhIyMLzOr2t32qj0/lq0ZQ
KPHnqzUfs5OVRFrCUlVCyoDefMEOljXVuBsEGAvJPhVYb9ydlinY8r7oeL8sxf2B6MbHl8aGR01S
ga68de9MnBJl1M2yHqRd1aqsgNMT+Uuxu+cJy7cLl87HGiDXiTGbLuq2OnIeWEV4xxDmlkOGern2
veV93xcAIDFZsk18zjskimgouPCL9EeH7m7iYDnC3iPQttQvdtY4NMBTihaRSF3QU7ZJEWCho9SY
I9F/sLBt16Tw/ozG5O/IuZVRwP4iqmXvvNN4VBmrtl/vzrJVxZd51lqzJMet+UWwY1pEq2lZM/AY
NFtdBF+HVkJW3vQFfH5nT31yOx85ODgzh3AnjL3gxFgFUkfbpZxJxLCaxzI7ZEPwxqVE7juxDRvN
xMPd+E/BrqA67ZB8uTEJvUb9NAkmmxIjBRykvDTE8pram2+KTafLZS0tTFk8DR5dtWeshnFp9e2I
9R03337+bISJ+vvcvgDOKI4gZtbPic9RTKe0hquiyxyVBP4gAIrloqXameBCGL/IssJ/8e033YZt
hAlmOm6Vnru+O30g+sYU/75RiUIS7dBI3TLwWbclAqrczVE95GShMPndA+YMnR/FD61YKymGEjwy
25SgPj7tj0v0NRblkDnm08ekN27MfwPk8jUh1053a30viZmFTzedR++/ZUmleSVCQFnrDRfesQSP
8mlitI1Xmr4KPocqDn+h+lJlCm+5jqdiezULO+hhLz7xWdTdGaQAr5CINW906o+2+LyDH95UuJ+l
Z9hg/2SI7DuP/RjYpr+cHdDsCIaYFYKGYYwNsukKKXcLf9eMK+WhaRhbPiOmbnwajBpenCEelvPs
SRidbTyn3zz5qBSYG/nZP886VDsqX6AljQwVzLsQ+3yB97UKKIq1b8C75LzEAW0ltHQsfLioWCs9
KdWUTxon1PxTFDUDOXhya7wGPG/GFBGI+nbS0enRr7BZLHIKNJR5mip5+Ad1B181Kaa0xbe7gjKH
mEi1sTKE1jUHut2jOVQSYNVpUBxSDgi6u+zLXdmQgvaRFALgDVh2PlfPmJ8j68QmW9y/Y52w8A2M
VLlPCC8B5/CF1Hpw+l6try4XZ/E9HbjwSMU0P41KKXh7AU3h1ILUpQxd8VNn6ckPMbvqxeBrquk1
3RBcbMO80U6JJ7Ezg51bTBC2I3IWUnrtu1LJo9K7lUlmWC2BAp1RyNciQGL9EGikkASiRLb90sNi
ExvV3tULCbT4Cjq9ZHQR+Iq4xAT9HOPink8d0c35wXOP0iOWiG8nj4fKFfS4/ngWDwcFOp+LmIF4
Q4nf1GDY7lQxe92w3JtBTimAdolTjpL1UiogXq9sADnWStFiF+5fRpkSC8hU78WC2mrp9s4TvaGT
AZEwq1aKWbWbM/c+WOiO4YPqfjOpy6MnoX0coOkRIC9Y/t30l7V0u8JDTplkKBDqS8taB71MmZgJ
+jxAzKUTCgtDeYDh//gfeKiQZ86FeYKwJJMOeirGajWPe4pAB+ROmIa/XQlMIAADti9i6OSYDvkh
pl9gqIA8AFXHQLkBzuDkoHsQf1APM8kmSIgKFMH4CvtC+/n/qcHLoXahGuG6HKppE1gPHT913s2H
LU/lW1uPfF6ia+rUGBuycbMGLgS1yulGTg36kBhWzkfQVIZancxRaeTGJLabEUWyAWUDfHQkhv48
Qrpw1Pm3SG0rrcAzEPkC6ZM/4yA8Fh44FWVoiCPfoEWmeI1QIJkO6dL+9JR/tDOLWEf12nFV36Sv
cmLDm6AZUYDklf98csPaemI0zpkYKSduGMI7uJNrwmGBCOjAJGpbejqZeeRuE5y6TBA/a5tAQbln
lUAL5Epa3TAzURMDTl/dENzy6+8WrHr+FVEIKp/lSKlrAbod0tnfUuQUfn+VxKVFuCsRtVFYpGF1
+sfcGkEgKJqQACFUq/OKA+qvL7UA5nMTr5fdUqkXpQE8cFwW4CzTlX03Oxo4XsYXoXHhBni08L7t
IyQfLmSYsq0mzDA0GBGaKYe5Nbvw+mCyK8ea2l7I9IvPYM10bdZaKhwxBH2mldqJiddH1vU8/frA
lEi0sMurO818fJtnBAEimeaF0XcmCb5vhxe9T77MWVS40rIwRH+wTm5LLMWejB7syUHqPkZz/s6T
6GEhVfEPC9VgG9hisp1e236OtF529cuFV85CWvPBpDC+T2iKRXnOlx1WMGkENpQpLhwRlMCOiKb2
VKVidrx1DYMnliJ1oHYG3i0kkUqyG+OqmmUWtrkNB2Pu57nBKRvBMrjSTOrlBXSnJf1kJmkr8kWz
NeHRRLY6JQymPTK6S+TEbScyiSyVkcm5n1/hYQvOx/9QG2kASO8ngxB92Bp/2eu1W/80N9z4Tx7D
lrAoraJuyHJ1uqs3YO6KNTBmF6IjQipiSUcI058SMwefd8hI566vDhtJOB3fepbu8rIFsAxbg/Rl
5FJNNr2qpDQT6Zqt55+WRJtZsTsfPoxcmXt2tnTp5oNFZeI57F48ZpWYGvV9O3AOgA0X2/kC+FER
DQ5nFuIKXoFdvo+PTq+LWPM80IQkhd2T8gBSbzA2RPTk6akEtlcxEhF7EzUpNw0fccPh5/2alC+L
8PtD7cwu1F8SpG1/2H/VPUBD1INMRvyGViIr4sJdi5ues5cc4ZUO9dtczDCln+3LhJ7z6ug/dlXH
ZoP/PjPu0ZKKk4gd59P1b2zDivWrTtX6s2JWZ6IDdHsyG01Mqn2+eM2umHXt8T86o283UaR24hPm
PGG2TD+Pm7Ql2DiQmI/CUfD0m/EyUBFrbIx21kDE92CJZnI98cjqgmWTl5DzRRRIkfHF9qq1Ic6N
IVjo0Unmyxo/CUgzRJ39ZuMxcLpRPIHdrR20gHbN7w49upUIYj+VSCBkTBWdZcxg5FcvMN+Nt0/N
YkIFr4uHc/Jb/ZaZebY7FsKA6s6a0urmS9nVT2LPa3cpFOhO8CnMkxBzVYbY7UKX7egKBsnmaFf/
HYM+HbWoR51CcjSD+9soF6/Gv8HPSetJ8pg5uCMu7kmLfwahb6V4+6wGE4XOlRBA67nPRPVzhm0A
JcRqTKRiDDuNMOWS8QYRR2cx38WX91/xBbZhb0V0R7qHOoc4/UcikR5wCNXWIDx9O8qLaw/Oxp0k
0+PVQyKota2uWyppYcTg3/CAOGCWsECeFdykIcK0n8aZ6L3N91GaeuokG3DkXrSUclhquopQIHXK
FFTsxK8hHzRgIkHI2Tl4JpCnIuz5CeaLtzJGpevVNjR1TJVnlVeIprOZP9+8ETsDIDPehm2ox90M
uDV3xUXf6CTVRym/DMke3r9NjQ+sdmTjZ+/+dk/mMyIPGZCtrmmt7BK8laHaeBJLEVjCahU5u/DF
IIwwcjOt5r0f6hy4IZI5Ukbtp4VD6s1RLqgm2f6zEPhfWM+6Xhpsi0gPj3P+tOStl56x5/oHCS16
cjVMVi0c6DkQWLCtolYh1ZRo1072s8qR9O2PdhLPXP5KUy7jS7BJ00sYNdRlWolEgWXdjeY9Xx0/
cXZx2opjcOpYU4S8ermBcAl+NXH7Dm6IfqdPucCD6Dmq4lFs8bbWFBVKQV7KgeKEAoJ4bgkun7Vd
oaJf/PEoa/PBp6q0cfxdGxOR1lgrErajjiOwSddVUq3EsQ1VPBvyeHgArDxj6Ki6I63ix3K4A3Gw
v82XXTjjWbsOADq0X9XnP0Jb0g9IdYrRdUq80RFyxGpBq2rcXSIeLoEWo7bJv98At9+rNNJUNOxy
T/+pN2BmAdtfWPdSS0IHxwEK0Ev1+Q2lY6VcRdmuxMot2FBdKiXbVLCz5Miq9WdI/apvZmV5cHe2
/iqeQnNhs2GLsShrk70HchbJJTW4MreFRBAG0H0a4mEbUGfGlXhCM232bgkasAcTL6YRMeRN2ebk
lttZdzl53TiTZezG5fi+RWF4MEa+3T8zp0HH5RQnMMs93ZHtUVh0iqLvEmgDiy//ovSw7/fLYxsk
vWBzKkhLs8zDGD8BXkfQaQXXTGe1TcjRwzITcAnBZ4hCaHnOTwGnrWIhhgcLEOwjxDWdlfZuHhgq
Z95ncpw/UzPiLSPjkj6fgSflXTouYpIWp9G5rOcdcSlD2AqXIhkLUMC9eGTdoY59ysf2DEgdfDcU
hexTnrnR5oNGljPX36gbZrC+Px14D5AoTv11nlbFIatcpypciFlEUlFrNVtSdlHtM8forr7fVu+O
76N0E/gCYGuBjRI3dZFay8kcObxAQD+xot0U6qIpXE5XILaVLFP7DDj0s7WagO0tChTHtvaNF9h7
GqntygINKeoQxCIuB71J0zw2qa+IBi9yLDxTZUJcvDg/0iytFz8RXkxn5dMMclR0fp8kD9FrVe0w
VSPfRKY4PRUDE9qhF2Dc6emWP3Iu5/89z3tCdHiK9xvBDqViUA1lZ7XEUkCpRA0GBPjOBk9/6d3O
XNMDZ2T4ZWbhN/2tiaWiIyIjcBVRXIEi5Y+O7UXRPOxLcrWKiiW2Z5KbH76dv/FYnNQAEYc4kbQO
gEp+bKzRHQfLLdM8Hz3saMaloGK8HwXTXWJHLZhgBdfZAJtpv9GjJvZHlqrLUaSkJnxG/5RXzo5L
RnYVLmOmuMADIYIV8kqf2HxlYjTX1+4jrypcVovA6cTSLPeNXpBUIvxd3ur63kN4xaauQumKvaJW
I1Ur0nSSKf6JpKxPUil98r/31SNdGxQwTjfUd2Ei7pccmQBpVDY2Of36ebIlU/kjjvcGKP1hAI6O
bWiAYLEifi+8LwP/AeidbACThWvH51qEgH3whLcPa/Uaur0yTZdy7eHM6esqiffCQ/OyRtEh46H8
2MxuFIouRV9JEna7Z1rFe+hfLWjWvxKzLCmSoaU6gGHh1qSPn0HnWaPB8qKxJcGAqLdOP1lhYxQL
+x8X0hj+L2UF4gRmSDu7gUF3sJYtAzjaPVxA2qMjmXm4F+4qFlHaBUVb238MSepFfZ8RpVrIiW+c
ZTHvMU8c8enY8poyTqc3n4EZIvHOoc6d3nHywZdUO+BOunqpeWmq7VRfm2bVRzUD9LAdeiEcDfxZ
Y+MAwJChwT6In3R9Va6bKSCdmL98iqiF1Pg2uE7IFLV1cVIUmI37+1kSdJ1Xyu53WzB58Ww+iopI
iMC1VQPsddR4B/ZsVFGR4Sj7kR/hypJdCKxCChL836k+71Al8pcsRuOI1SGfhSh2KzW9SxIclIt1
y+GkhcaoDEfEu9Q5xgWkHbTYn4Kbvx4f49n5zlR7n+xP7NkUwukTBg6zojigyCJXyzbrwM2+5afK
QNkoLawQuN+GN0yPHzRJWUaN7PVxFCCnJqRRo5ut12rn+aBiy/WjVb6V/0KJFZJHgw2BDzBo7lKu
7ASUAobj/xdKFP5VgKbyUd3NbwwfsBTZ5T6tcsv7T5Ppj2kf/SXvmNIhZCNnDVMXeQhqkYcmBwgA
00P/DIVtNMkC6isw/Sr1zxozTWNNbDMTwUF/juvccGHJYp/JNocIk+1yvB8/ENBRP33Td5hQFS4S
T3OGUEcVnbCh5RpMC8N+aKk7Wx0BIg9M6ShG11n4snJRKhIIyeYyL61zolBp/UTJMg9E8tb5pwKM
M4tcqP+hlEP//pbgK76rxH04cNIRCo4TjsZANjlRidc4H5YbSoACjWn/SPyUeBaQQispV7wLs9oN
0dr8elT38X6KKHJGJd1VABx8+5c8f9yn3WxDWL7qkd3ebqpjvHd1rAiNxVAzVD2ld41J1rJj+m9X
6HFh85C1Xfm9rFesukB8PPpHjkXKFcsgZ+QVg4Ugb2a6ho79i2RfcWQkG6gf7rzp420qaRJYESED
KsJb4V8orkPE4RRX0RCOTtIXgANyLxWqFgOadqCdk5TYQ8ynWArHJDwr+rLmD4MmKrce4pzXgGLQ
JdYezNCNPL7cwDqUTW753NjT8CBoxWz5QPq9PEB/VHAY6yHmGt7chN8eEvT0yzhmwcgrBzmv4mYD
n01v6bEjmPgzX//aUYLYlKzb6kL9ZAk5c1owJBme9uIWTvNXj4rlpBeRmybrOOI7AOQxxYYbq+GN
jTWYl+QqaNs9UIAeiJah+MilRls0A7pPFDdZnUKFOp/+fUefJTVJdiB4iECPy+wIqvVQwBUoB+rE
2rabUwdGo+l29SPkSbXp/u+g8PAKun/c+V5MoB6l0lYlHXe0oJozhbgoS09Or286+LLK5mRvS6D2
RTMFOeCkFkHolygR3a6XUr3J0xk38qNPQe9PfKj9waaU2u8yQvri5xNBOnytZsRQipYMn2CWMff3
wuCLxhcTL45owdfUUgfoJ1rpy/uglbNuGTyr/rdWmTGgmcHK6X4sSql3+6FbkzaaeVMET/dFJLki
EOJY9t4H31W6AKJ2mv2KxVljh8H9PeAGgwwZ8qVMEkP+KZtkOlGy4HsUhZdsCkZWbl6mxKajet8Q
ZBDwPyAirurfk6EFbnbpGDHk7+bn4MnvoB4xm3BPKP3ybFrdCVL1M2M4f41+unLPeoD5ZoGrTAc2
uKCmnAbc/Os2/Nn+9wflyyr1hJUnKsKPhM3aO+yOGiezLBN7pdT8N0ZYPaubH4AGV49skjTeD7U6
t0zDo3cd8++IGSmqta8I36FIxBenghNOLtyb/7GkP//c9St6gwN+uZvuyH360Ls2kFPgFWMNNnEM
TaYQMG96ocgMd6et3+UpWYaioKYqoNFORSKaNMVU4+b6ASYOapxtnP5e8Rox5fS8C1ReegN8HwOA
CN0o2zl+4pAd3Q92Y/Wq6Ww5AntB3zOyZNwjMt91Y9d0Qtn/Vs9OqTdd1k2arKuq7p7kboZskIO7
buITLRA7tDcmNvd9ZoY6D9egJU17LwAQz2w0/Nd/rrR2zPgfcOaT+GZeBFqPCkRREyHJYnnVXp/t
27nyBj/amN+9/hbICtxsypGNEmhcOleBBNjoECbnC9gJryJ4d+Z2uXgIOtfJUotRxw0sz5nOITnu
CBRRDByO5T0WPPGMZui8RydqJWmB5PsT+d5x6rnOnKlK62t8aE847b9oNNUR+2/zQiWLT5pqR3+i
Rz3jG+8Kr142wmq28XjP/57xSWlMoPSnQCP9r0+Y66IO2miC6Ym6fBVf+05n/VjrF5s9BcD9ZG7/
I30orHUYqbRLm9i1//DahIcTaDxMiBQcnN9zGM6fPKlr5/gN2NjpvbHzo9JJq0Ho+PLkOeLMv1vm
jXobBUvqsApURZ9DF1BWHwGU5mXiDstjN+Ya/VStfUirltVr23Ttc33ywSvds0tgE57qxbSmkOvR
N4lMgwqhD7fQ0eTOA7TnKZ2I5PFciN4bROdCJEh7/sMPUrKQl50Q8NmML/fEQxrUd3/i1kmfCq2A
Xhmfyy65C+5Rnnb4lG+CxolELgTAjweptD4gHJObCo1FgAC+y0oXOzJjzNdUW1BF+MmWo8yAEs7F
aB45p4n2y9CcxsbVdPldc4Aiirq70y+2DQcEb6lkJ+JHmbuMpERmRdFXYJ+uEXA1bEFYlTyPBOYg
XasBoQGUNcwRvY5GdwTTaGEIkZnu6vrpkxrXKuxGulNnLkx37PgB8D43GvtVed8KGSlDvFEMtFvL
YlniBgAoLSAY46ctLDia9jIFfU6L50lrjQbOotPL4oWKX1hUZmEECeb+nB+fN9ijSxWpc5xqVgnq
Gpxa5qGJslRrOgPhectOEVIfdEjIoeZ9yZiCjyOWf8JFy4Jgp+JjD65X9+rE/BJ53IbC36dJUndk
QXZ3x/7sGQ0d4O9Mw8i+bWcGHaPOxZEa6mMHOpBrJsNqsI3Kr9aqTnsFQq6RI9r3jyaZ5s0K43xP
MXbyHS2+XypsfD27+0xCSIzZ+AK+i7xhiqN3+uU4YIuuQuqGuvktRoP2AZ78Gzh30SkZ6a1U6kG5
N0LRxZZGAedbjKqj2W5v1G2cpUs3qRmzuazuDHQnxtzTcxThLTtSSWml8KvsWPNjdgMjeoy7Jznc
rZExeSaJZDQxkjP5MWDOhh4U56D8nk0Q0s/MIdgfv+xXx0D4SLVr9sU8e6llChjBkZMz/e9U20kR
9akL0Jzb2UC3GPMSuIKj0qfySZ7IUmZ+zTYqV/kPXXdvQiP8mEha2XVnJkQ0HcAvQ19QuHRff0fl
fPQGMLMDQvwYbsNPvme4QY36TczQmoAdWtmL5MR9L3A91QHU6g5dL3JAKoWW4NocGUac+72HghKY
gFCU57YL3D5arkcOPLqGOWSwbrMl+v6QTqQr3+FjnrwKq6hPRTOtKCFblvJ045kNHlECqNsrlvUJ
M3tDypDQPrJ3kgTg2lB7wRoIE8uHvYZiwXSPIRko3l5xcFSYqIPQ0ia/DXNu2LBoUJd9+mXAAwBG
ZOZO2atAhtkf0SSq11ESMeNuWf47AB0Z+nJZ8z/B3C8A3dZkmTt0uzqQIe8DuTE27QI9Jg0Km4o0
72i1P4WmBONKbfd30232cWkvfXG2ZZcGkNMP0L7iPcii4oqkkdEOb/BPxCipS+ED7tA6rUtLVA8f
6k0rJ758CbyKfeKxiNDpz5oavNRnGDQcD/a3nbRBEQAeeO1UMvFCAe3TxiDO37UfI+PQKR+cJrIZ
qPjbFxSXqp5HffLL4FSvbRMHzQ59RNA8a7lnefHwtTXuQEW/9xMtY1tvDry6HsMMxzNF2m3sdOwB
LjMWyRUqYMWcjNoekJPUtc64815rBYrVlhkbo/QqO+3m1gEfz+1+/tatr+NYXCs4hYHZ5Fk4Ri9b
F+8YGRadr0SY7CUCC5ZZ9kK3JZucIW/IhkKmRJQSNMRjwTx2C6WFIGPC0skmq5CIX8zIJ3jN5110
7lZ362S3G+YCRKLCtvXMHcLjE7EyhcD03OKC34qnw+AYjwx+MBgYCk1s+Hp9qFVoCNv+FXWIr1E2
FPQ357HeEqdKDaded+9Kf4UUaLDTO73WXu0eMHvRsLeOepbN6v0ibUjnV76xPxCGgRpzofJVV5wK
2+C3jbd50IfkcX68G5p3Lyh7B862WMT8RHZJXqLIy07CDUBT7wjjzKnQICWFhV6Vi0E56EZvr5nC
nykHDHIHmq3Re28DImHqZgwZ2VthVzrshFlK+s8bO0VLXWCVDXodXkpS5JmcaxyVWsEytP+wm1LS
mNCvHQMvebzBL1KWndq5oUIs2bzHwP8eRtsmo4s0BZy9lyA5CW0/nf9veogWiN6wO1GLWzDF+Ak3
roxV+pkWV7mFm5UJpTJNug+yCtFXBrzRnTd+nQXSPGFAhBTtQurBGNse5u22YtYmkTBdK+T9DvwO
o4dmZxNo6lgATAacymNjIzmJ9fRCJLkA0Uh/ESdoS2AaRiME0fs+A0VHXzH4x6SZpt38bq0o/v35
ARI0ssOr+eHYstxT2QponRUyZ+JFwoMv+xUF95mCV8kPwrjignY63K88h3zTDQJG5Qq9jtqAMkHK
FjT6r11JwgwaWfX8XK0pJtYEVS4kY6kqS7J5VwPZu2tXJqs5h3N1L0iFQBXKGKEByx7ldMweqgiA
aak9iKd0bQvHuPfUShQAjx6Xcl9xd/bgarKRzNYsMH/ELlMJ2VRFKPlC83UQ1Pn15L3OGBm21AUC
7wm+cTS7IlUKKAm4mz0ib+7W6LLpTPFGNLBBCcUw25vRv947dIo2qbbNDzB5Rj+04nQNUn4ZIMcW
B0tlllmvt8CtIAfSoeQNcC/cNKrhlIqxa8ssRGq1O8ZqmbsAjZ3XJJ191SNXPDHrh7937vdYzzSY
SNq7VW5IukbQqeHOdYXX0Y9pmdN8vrc1V5k0Ofwzz2w0YAUxUwZe0cYSSgp6Bxft15M6E9709L//
a4HQECx6SpFg0HXm/dBCkUTaZmA+c9DAx0wPrqZqhQgTv12yWn3Onzi4l74ZLIc0ISNuHfzdX6VJ
8ToUYSj/4VN9+1L3rxw5rp1eH6zB6VIjuhbUBnUltfX+pywBEqWXtj1C2NEa0rfdujDNeMSAzIUl
IcNgFukaSFDRXomZbOFBh9eDGwUiyRxkfia84knUmoXQdE1hPrSPZSQXMLSJQ4R+mQ25eFQhkAYT
+0KvicpLgoseUPsu/ja97uR2zoQ7iAhAd8W4H3YxhaCXcEOOhUjev8yRseYoSWkTiD6ScvPNKExx
JOaBFnofuD7ns+MkhVzZxvgAxXq2I+OHR05NWroA6qR9LnVXkYXoSL+KLpkJRLMMHYoWEb/poY/E
ZoWPGgJlPJt3kAulUW0/jntH5aFhifsTRSNd7sdbtscdSUqIHWeAJkUZBhSJRW743bNxRC3BpVR4
Rou90U/qmd4wXmHx4AZCZSYbZm4uuyHhUFm10cr2+eTfZ3Rc/3hbCFxrxqCp26+g3bhbHaNWOe5d
TgCkhLsM5FWChafOgaoWY7u9D2UsLcK5gOIOyXO3hiyelt2EwdGHNij2x3OdT0wLP7IYWcFWmaU0
kHdbfFU8XiX6e8LEwcHtPlzK/LbRf1tltN/nln+dJgaTsbS3tCKn4qgyNC6AJanug5m8xZcjsXn0
wVZFyY9X2oT8fZt+IMR5zS+2vMJPb/1r0N4U3LbbInMPHy9pbSsPrHAR6Nzi1sA2ntBnTkCy38lf
f9RLsfDXByL/fw968p1bPKCQQfflsdGxF/1DRylT5ilE5WDdOZOHaK7JuN8Frpg9LR4eHZ+HZF0V
WXGPvfITqRgz15KOnrLMCaURYFpb/n2Cuteg4NW1TyYh2RpyHajlDKti89HuNgQhp9BPgmXhUvwm
N4CK8+rZPuF4V3lo1rfkvC4Mc6PLAPgLxtvWZCEcCnpgDK5KJTOSp7S0iQAC1lH6CtF6Z/CapkNT
2X1exhaNCs2GU1P4LpaezERJ/iot9nsw61BXGK0rhQgpZElGdYbiTV7pV3ns8rxzslWCaTipTQ29
9oBoZ6b0fKNKSuZLJ71LWYtKh0SqrCmSbB8g/ipqDCigEfGPQedFB82hPff8O1Os5FkVHgGu+UMz
tYqBc5gwYVVpUqYsCaots01ORugS44dOsMu+jhtgnz5io9Ilde/bqwhdXjfwyoYwk6Gat+sYYBQ9
ni3a2HGpiA+9a8CCT+gaAp5IRKW6bgUYQIUONNsO+Mm5sxM20+L2BupzazpyaZhyS+h9vydVdGWv
zkbLzBn/RjlDkxjoatePJxUkVCkIrfaFFjupiSvu6Lmk7D57cFkJNMsYtDDnbOg7djJBJMjAHYIC
2R4R3WLx7hkkv1N8uhvvoT63Y3V/+W4Oqzq0xkDwWiMAd1bjtLsez9QW4Mhv8mwjJrrbK6mrwQoB
wmdW0UU4B1Psj1g/ymSQ82yIne29ALYiReRwHv0k338uhgNWgEMrjv4Y8c5aAxHuruZe1aG4oCHJ
q+QwCgBSOeOnfTkvIp4yctfRNBJc3bHntK229rY99O2KhdYEzpQX2Xk3OUQCIUy9T0el3QTyjtUv
VvQl9LqHua0v4d/HjFIElKSzUPmRiLHGYcWWjNqW5s2bEa4IfH1/AA+T2pTWZYc5PBGvuQZe2qB3
RPGCRtZ/OH5K0sqvox0TRLqqV+mUXnv5SmshnBAlkp76YcybQyedv0uVJnTipwS8GqK886IW5pXx
9Zzlbx67XgOtiR1EWBdC26+OGNjOn8Hd5LbYZnl9hExCLuF3h5W4f1ekcN5sQbuxDEhkoOLDeDQ/
Mf+GUpM+gXX2QBXs3QYJYlDOgo+uAIYnA1bywtfiD2PX9fCSBRL6GNM7VNs+wKzdKtWD/77NIDbJ
tXrrSiNYs/QfJvvn//JVnKCh4sPYgg6EJarkxOqsCUHHMGH8RCgymm5q5QXfkkHC7bvo5qBpKe+V
/8O6+hXjO+ai/6hqhbNoMhONeEQ2ALKZLFxQu1aXkE3BwYLDj7UNE7DCB+uvr0Zh5kKejpCXz5ja
leKVuKAEMRCtrpVO9l7b/ePEyriDw3NushaMBpTb6KVkQvdoqnU8O6LYotxRaWWEVafAIe+vJWdY
57UrVnwKpEgEyyaMxLbfU1iq+HacNvLh8vyH2lT9YYuUfZxgUrHgJviXx4b2AU1DvyWv0hTTgoaE
D5zGoIHTIEKGHG7bDnXjtN/BwUdVBEe/L56V2EbyzmpbZFEWt1ZWG1Q+Jijp7+b8z44icC3GjJod
p1PO9tAhumJMYh7hZIaR3wwaI+Ha/vqgYco1JlQzuPndIK6pMAHR1KsFeGDlTthd9XpCgORgWAZ2
Vnhz64+u+CjCLbA/tUJPV3ROtx5iSp8geOIubMwz4CtWiQj0xIvqYVWVX5yn+e3kDibP3t6ILDHI
wf9RDEDjwbFbpuoij5aG4O8Jg9qpLPHHsgURkUgpePY9ZedMuNnwEmALdqp1lJ1pjoE3FiWfk6hu
KSBcG+yHbO5wIo+/iUN8whmxc5VCkjaPvOJexZVHc4+1igW973qKbCXmsSnLd4nQC04tEJwhpXjB
/uNjspvkozHhZDAwEm9nSszGy+8n5IXHGtqa6zhsVQqgTLYDog1nb020qgiPyXV5gl3+gjeodV9X
UqY/kcS1pcy68yqL7o5Zqc5gslyr9SpvYgjx/RE78BJm5CwGpGCo7QLyj7Qy5D1vxhUsLJVIHqfu
JsFV+qYYEmW/Mn6kWB7Ye/FlAQITVLntnD6lEmha13XTJS0tSI6Xa/z03N29CaO3+Zo2pJUS+q/i
1C9rrN3v5j2p2Ldm9W4NParT3GRe+j1H73QgMQb3f8F4MlUaiHx/X18FImuIEufOTE78mONJd+/X
v+8ZUObe+Or8cdFgZXFgzd6wOyVre1wY5MTlWA535pgHl92fqOOetUwGwDiuZd6JeZ9oI+ksJYCQ
51psBRDhwKnexCHu9FiIAqK4Bv3TCLcJKkUlQ5mswN462TZrfdE0zE0LGWz0sjxlGWJxqNJ8kROx
eVfiikuYIdgt+pNzSZ1rXfUEVRt/1yjK2C1hyMshCoMrw6W6ljpsUYxqmOutJQPnmG3nhjcj3eVx
dlYL/fZm92fRiksajMeKDERT/CEgOGAr7k6yGzQYkdMBzK1xif+nZatwn+QqtGxb5TDnInmqJMeR
doS3PpR01dXJTa2NuftqGoTKL4uUbvRFzpS8DPsPDRk5oE3zb+M3mE8MUcyGl7VKcZUKzynAJ1fg
6pEZOkbQmeyhfLHBNFBMdsRLLLiJFsSsyVHax9NLorx7FYK0MNFkYSKbOyKFivGxzQc9In4KF1pl
pa1KqrUHflXF30tnoYV8JlG9ctpN643qlbyt9Bvd4RZk/IASlymM0E7jTyalYbZ6Rxlfp4VPzZxy
RISJ1uf257rE20sab88ZPR1LtRT6gsHKJpZP9wRS2XnhMxz7bBR3/+Xqsvv446HKLf/262+mNv2S
oDh1YjP+v+dRuoawfCyUVGDHkLcHRy225XpggMk0jQLMD/s1+4lzDoUJbDoM/j6E5va8YAynPiZP
JtWSA0FaVk1/hm2lBxK3ZLGoXmCLdQ2hEeJDz5dNWJYP2VBXkIXT5jaM34MNHZpTueIKzhmEBiAP
fGzHV0OSeD2B/YHxElbRbaTDhrghhMAaVFXini8K5QRIjHv9ezY2wGi9fPdIJVntAM7Tf7k9yVl4
DUZRmlmEUmiC72EPUrc6OOoPLxBHe1MQIkHCj+w5go4oULFyO0Xd2dvrXPUj4emebNZ9dHSxbm2Q
28ZUC7N0FZ8xSody6fOjozfASL9kOqoCp9hQWWYgt4Q3vE4qgrGezJvIso/mZQAlTx24rYcf2I45
AfWgobAH2cAofC2AqIOXWsxR5A4jOE7ft2NS9bNRgeSjk4paSRP40coP6ZVmVR0lfSg0yHK8LoEk
UmWJqORL6Ry1cLmmC1gzSAlJ09NJ+slfczQ7jETmojqMSpcxEZwfy49aYQBJstXw41o+Ogti0gwr
0Lz6fAdC7eSeVqxhHuy4XmBO/UrEgf2qaDKpp/OlH0uXv8ipLfdk7Mup8qeALiOlZ8KETUK0cdgE
9OF7gjYWD00yl4XG7ajBWLtROpUlU7jnVQxrHio4mvjg067A2W/Hx0WqmEOyTFFcwfNuYrlCt2iz
cAnishO8pcXGGx4gaVC6PMmf/SLfOoejuG+R6lFIyd3S9lrdxWBGqVKEsqFZGBM6G/jre9UGdRvb
xVCarMen96iCDyw+u/RmVlTQ/15DEEF9AErUPL3u6fEseQKUvfYGCHuN149ZjUUuOyjtRbvgnlOI
hnbr5jaDeMY/TspFg2L2q84OkAVBfhU5nCcdvEgHdKiUU9ev5Lu4HGCWaL+zkRkjDfCl+7bljArC
kMbmA4TFC16AxZBuMsifajUL/oFe1t94fAxzjzHxovY6fr3tTkkRFBYt30MVPiSlnfiQct/C1I2I
8oOBx9SeiufLxsj59FdDZxq/d1zym2EwEcpy3ItrIXay1iH6xYQWZGGwVS0DBp/g3D8HNpinl9O1
W7oHR2TjHd8mLcwxAxHhMQcm67A8qw5gYMsN3+opo6nA0Kg8qX8zem9WXbCPoH1q3usjhnL3RMkl
nQD+Qg6n5lsHkr6hBMTLJendUhJqUDBELdyYfaaWD3HLS1Fx65zIB3HrS4JUwBzQ9IYR9bFZPh0Y
45fVShYDW6cKIdMvH7FkxgClShxuhIFECGBIPL+vYebvfaNgFiyTr+6iKdtzBwcubQjs/WqvyzsC
9C2nfMKr9x51InXkfZPtwA9/aNv6ok6YJiCEVEB/iXudoiR+SNIlI6fLGT/mt0n98pX4Ap/ov0LI
uMYM8188sdQQb5AXSx8/noob8JRrVs/XgHF3JXhmY0hTWxIJeMUoZkTkMPcBqW1W3vPWKTDpiFiq
OQIbz5T9wOu9+a8pyyxZ/MosxnwVhuYhvWbJC9iZHCJfQ1/uhPDPuLUweoE5oGIqbu9787pnrOYK
OMpLZI1aeIHJbeQdkDzW/PIbNHXIIpz1MM3JUaFRNycF4kgDvWEWmbD+9pgkuwG29MzBxTTM9rxP
sSoztzBV1vuU5ctXKDeRgYJl7Q5vvh3cUwv5qQeW8WdNJJU0xc/D2PUoZ89TBG5v9g1jOTOe4/nH
7vsdGFvUYxYcPkXsI7q13tO5CtJgYHquRiMMnMfpc4Zl1AFoPXebjb9kyNEnF2cMD8SGypA09eip
L85lKXDoyYGlE3TtHi63pDCiFgAxCuN3TDmSxWinpByb8s93S2C3N//BcdzbQBGbRrxYYc60O3rn
su/xC9Y1Y5j5oYDToAiOfm/RTOogwV8zP9s4aKSutsAdfQ1nMG/Ex0wuJehLJrYmoDyiaP09sHpb
1QbGBeVxM5+2smFiJqyLWJJ38xLSXQD6Vrs1RgAwFZDT6vcFILz0H/WslKS2K0a62yUGmXY1UcEW
szEehbXxmT6ZL9PeXuGBGnMyualY83ncknHSqGRnieK0A90HtwdB9m6pMdAH2peSexBEMcZA1c6C
+kWabLuAOdD1TMDECIMvVhrK10ONP1Ct/jc9MJVqU+SY3+SFG9driepJ4QQEp1WyE64yXCwzEdXM
R8GKBmmGg9RSBVrNz7eJljRNjxuZEg7rT3RvOtBamN8DopWIV7Os4+qYptzDKH/gisGciJT2qxl0
VDtjtWofqziYBdQ1vPOGBSc1KdTAWdPLBSD/q4UgFvqgKLGQq9DDrenPN2kO39ji7bOx1QMAuqiM
xOrCcIJ4Tm2naWYnNapGJ/ZGOETA2dVbFNP0tkkQ1Um+H9+crFeqSRKmnHf/1JVz4hMA7coo7gkq
xa6ZktjryrDP4YD3GkWWW7cQypBNZrPoKuRwwTHFnIFudKVFBr3PrkHJf5NJYdzW26BIY6s3tNK5
crUSpgXdXuG9TokuDrMgKXzeM4uXO5LaUo0qFP7wYWOj8e/PWUDAquYNbQfeaDk/JtPYTb373m4u
A5LwQcfVjxugCHWpHeINeeqRa9lU0P1jjAeLe5EyPzeS5AxW1ThuMkrK46cFtB8ZdwfHZ7esXTJg
xF7lutcnnx8rabbMmAqWBIXW0CpStWsJLdfDuhDLROLZ+hAzGTxxEIHpeGFcyt3cI1gQIJiNDmzH
il2PijwrnGa7KqTnd2TLsJ/pZP8h2i9ICKGMYbBn6YHThLigMtUJL2bdyIQoduALcPf4eoDMbRzZ
IliwFSbIbflUkkRLqg8r2zx1aOktMyQp6EZHreP+eITld3Llb4CvsOD/mJ1rcbN89UutsCBGEmby
DaDvGeTO9GHjnr2r7SgYt2T01C4y3OTwvXSe/gaIKb4tCvzacFzT8wByYlOO3um9I7kifCUE5sRa
8/5BU8TEzkvzoqZL72EWbg+tMFFxvD9jV9zOZB/ctrkZqN+ZiTkFAqdfro3rkDvRdeR8jxXc/wOJ
tRZ1VOajcGjLPVWO1cBJavZBWf35BTihkPjUOerio9x6e5TlZPWkLb3m/DggIEJn5XP1lPGSnp6f
3qG/i9A4SA8fdje0Rw08eewCNMCdaJ+VKhd8fPhuVmBK8w3ReHe8APsLfy31ntVzhKragqG8aT5C
a04X1nQQ28Sahpw+AxDnR3y1ZRZ2bAONmtGH7Mnn0r9B3Jq/G5oUZ34wri1XVy0CxrSzZQ02QAcj
dkwiYn/dRdEnKzfnGoOrJbmQbJbEzrQMIdOGRwzoZQAbL+bMImJnfEsZZF8510y4jVNOJf7lIwR/
f2Jjebmu9wb7TSbFSHApZCzaSn/4NY+mBBTtGmxKRABQVaUXK5uP8RmRQcaqq4Ef3/6XfOtFeKiN
3Bw5tS6cDh88CZHxP0BcKFU0OKGnQtLlx+V1OXx3qAPnsrVUhPAfo7FNzMQVomOmhXsutdDbT+3t
tMq09ZAklbNEqM0azjitsIP6QdPN+4IztQj8flqX0U4B6gi9DURc2vSXC3gAIKDxzkvWQjyH/g9h
E1Hea8OL4CDbdM6rlK71YVz7mBxOHhiWTylUpzm7Fg/OZekQguShg70vIn091rJEcpUsERa4nEIR
9YLpioSIPEMCKhEDZp/q4himrjSmNBvpY0J2CJLwenzBepRpXvesbRjO/ovfEjROOQTEFfnIllJv
DocOUpIAeb+JAcxr/MEk3f80SWz7e+NEmCIqf/0Sqc6Mn0S76QeQURoOc1hY6A/gH8e0a+r+9uSf
F1w93YnsnmmV24SvibfohNaZlehPxfvkGiPXAD0bz3HNjZQ9v+LLSj6ipOCDYgorZJx0vAd7WasB
ZqVBLhxpdi0LfbU38DhjORe70NWYTbWG9e1A0V6QC68dq6FzsmAXli7FYDMGsNhonJ7HcxnaD7BY
odh7dzDBVu3Kazn4nZS0qn1fuj1ZGFH0oQ91kb+akhOXllkoYsPKpfcyi+lvSOX08QqKuifGrRB0
qdSw9rAjKibkimC5CBg/K0Kr+84b5ZhCXR5VlIrjuwdtipgvAm9ylI7DWPcobD+uF+GIRFI9iGRV
8nWakhFn8Jcsx7NZAAqK+cGInjgiTZS859Q7xeiiEtyEbvA0mOWCYa122pI3184Y1eYck4giMeuG
M9cc8xVKO1+7VgGHUlGlVdwlhC/AHGGISmjEzDoXvGEezeF3KCfyWNFyoStrELNnBkBKgK1FnTrs
Jla2c4q+jlX5zjB6wCeY3ERirDziqiZu/7/qHH/OGS54PsxDqYsCcfMQjydEwHMXpH6hpqZGhkPB
d1f6+qR74V1dXj8JUr2wu+T29mU3ofjKk971eBrje/MS/GIqMQnTr6totJCzSKFoJf5GM1LUbiNy
lGgK9uRvydTWRcU5G+31U8GluunmTalsu3JbryK5ZJrjQxI5IJa47DZkf2BZZANVcDvvpdgLjSQt
bRWuHYgZZeOpz4qCCCHhCY/LYyP9bmntmOlcssUa87Zf14/5fjSPuQkB//rc5opLZCGW8/fUTeMH
10gSmQYotVc/SjtSStVfRmAXwJBs/caZdFT//oMAscD8EYf4aC+dlPyzFO/V+vD95nky7J6xsdmw
m42AExfWqtw4gg1gZo+UiqZ3D2n/kRSaIWN3Fn2bg+6s0CDnxGhzua1dHRz4tiveyjpvGDBU+nAA
OaCxcDRyPwoE7Xw6ciUHBfhL6nfKRd0vm7qBYZTYAWaY4FJDwwoZxzoS5WAdKXJvb5hfswQU8Y0r
oKCFz1NS+W5wLTTdXJjvTECUUMQGP3b4M9Tj9ju3/ggL/KCOWIEm4gwMFPPDliWnYcJlpgoJdv7w
I7K9kTJIOhUu9rG9GcPlQhlGa3E9h4lFhFImkt/Uk2vZk+7mKnQerM2zfWj5tPa/BHo1ieSZdnMz
91TrCrmIJflRG+NEWEF65ENSlGnJNFbg/3dsjxtkSPJP/W2gu4gsNK/JIQChJf07+BJV3t097sff
tidUOoQb67tqf2FHj6Qrb4TimrhRMgEt6uYU/utXTrZJ5856r11rkLo6vmHqHym76+TR+KXNIOCR
4ceBoiQ/Pxwjhxo/bqCjt3LPDOvqQ/HM+YfQLO4TWhjyA6eQKWaNhltnS3JbITDS2/iRUBpHkBpd
VG3Zfb12xmhFHDeb7bleG8ZbOFCU7+t7/cbTCYr7WQybBRrkn/ZWfb+ELfLR9qdPYfA6XsEoTpvO
q+x6BZ9YPT4snkZELnz5ddtuB6rw7deuDSRoJhcWzaBdzXXsmBT4+R5pZL+gFZyRoSu9uIGveFZJ
tYrJOPWhAxtvDCo6zjkNCtjojLO1yl3JN/5ZhnHgL8djMMTKJGQt1vNhbuIR3jUwuimbg5gp+PH3
3FHTIPbbj0XZ8FET7xW+ZHNkONv5sOhbNfAD1lqF3PB6KeS4xMLPmK2IUimLPoYnpnxSqdYThQP5
MgySLq/cntj/osrq6n/LqGW9GOF2uM8ETJqmqhConWTkGxNCP+RQQP0qG+U1A9ThpQlfMRY2euY/
YMECjEa7L/EqaaMX3oJrZHtviy1PvNloSi/zVezQyr7bR7YhNucllcE854N+g0fYZ/JiV+OZoAIf
IXbom1C6GlCmtCWGB0LSbf9bCqP2luB5iPUS4o8grT3FpP+wSSrq7SEZGGVu6mDhykC+4RUeAH99
mPoYzV5Hc7A5KYVmUIvaQ0aW/bYJ/SBBX2RkC7HwkPh24e8XhcyHsPbL4/w2zu89/16UPp1Cr7rI
FKyWsULQl0BCTMBO1noF0cRKCmlEJV1i2u9Rt8okB8w5ySIskpvg2/Iz1jYCF84+yIwKK4x0WMbk
Spbito0Sz5M55+kI4baEkqrCRdDJBICNLDuSEPZU6jHL8Pu9LVFW0MgIL1ETs61xEOrtmSn+G6cK
NgnN0CPG5cz1bGP8wTYYpz5EN/qP5zJcOoz+Dh75FGCZmXEykpA3QsAO8kAMnx4AiQbFQN1QkJ3f
bjrt+G1Fbb2QZQ/Sp7ueWFhxxo4u2DpYz9AUXS29PYLje0C3JtpAL+KQERDl741V64v1hQWY10J9
KN6vQNYyOwDdyolQCDcJCLgXAY2luB9aiywvcBQLZsB7kTfrygjXQgX17EQpbtDCIPE1Zw/Wl/ch
DgCcRNfM7b/PFFkffjQg1gFao6BDa9bfEClmfwez6Lc8KIndZmFJRdZFuy2/In+LzaqSNQh6zQbX
4BtTFdFasrI9rNJhvpFQfdPsuS5wAxFzsE5ofyECcXg7sYAYG7774qqEWFne1AugjYMy+WGo8lzi
ODUm2xxm7L7eca+ydakwyb9mi3sa/XRsUVOmrW4YEOfFZrcPiQW+0QpZ1C0HJ+V9b9Qnd9rFBSsM
xvRxcidFWEtb9Ge89ha3jUe0tu9b0fxcJDWfW1zGVuBPQCiuJpvQrfDVtEVXgPKBo3kPaqjPMPKa
5m2nFjeLyc1VnfQMV9Ih3D5Ai2KOtVyfrErd+MgY+g/y+yazQrc0fzwmUBoQhquXqocI1sA2Ltlt
kpK3kINw6sjUcShFHU36grnmB3WH6jyy5wlrJI46P5QBg+UyYQ7yhNg5q0aiekz0mAnJWv2xYrxM
g0jOL1QysniHHPIn5cuRkze+Un4D1NH+Cs5ciiU5wirQp8YuUEvuJ2m9GB0y1qvqE5HosPsdNwCH
D/SKq4dghABEUgT6p03mMGrVjk7kixbB4whLpwqDBO6TGL4G4Kc/ZmmU2LOYJ36JeQ5X/0CUcLfa
PpcHobCTAJOdNugvj+xwvWTCUta1x68Sll8ILiBWZSWvB9aP+deYfuYY38gCZGzzZVqGvTwLgHO4
Gog5KKlJQaBn8gzHJYBkEUylA4sfTvy5wS3VpJVIOANdEXTX5RA9PP0uk1P8nMHCVd08pLv3n/4C
hoE0Vf5XCmhuh/LyC5H/y3SZquYoVtTUy9WuEqY2mJO683ZqyTwPvbD44SilpDWqTxchI4WdenkN
gYrXLhHh4pXC7dM1gzEUnz4GEwhsOxhM0m7eg83hH4HXqZ+numuRMzVi+v0CKPh9Uynlf3M8cAGR
w8BDbTXUF9oy+PYFzZDQ7jrCr1rk1MDe9QAx1ANeKiFAY1QkpWBQxFSOPyf0NHV332FT7BTM2sRr
lG37q/r08sx2Fz+Kcp3q3HJ2x+OixySKBj7ZviAk/HJH5r+d0WGfEGMCx0MZSHjN4jGbjK7j2kZ4
aMpPYcCY7h8UekkyLA3/NSMaKHNmgFXcDTr4uGZ5GBEniGiD5YfJAJ/O5Ee0lZplJJdQAa9IQW99
XfMZ4N5cg7Cux4H0WGZecUyqfLbF/QInsceggsmICWn/RO07NmxcTKtUlCMxLobrPNQdrh0eMvMs
2FOeIekW/NelYEaXHB1g8kAFcH4J88GUkjMCRD5P+Wa8eEWo+0+Gs85XEiNuH/nEKfxR6kZ3oy/V
/IjnTm/KCgr5gsq+u3PI8aQYVVVm7cMk2+c23e0lWUCLd1w4Vk2tLJgc2vmy9xmVQPGINjpcG6pQ
cqcFwkzS74tjqc+mo9WYwuHg5thP4xJXUWXKymUUHY3SPBwzRNOecaIVgNP8pz0kZzMfQf4hdvgK
rZN0dp3xd5TXdNBfwwirYm37CRJBKMLbo2AQ6E26jZFSz9gEKQxXKEtoyXAKIIveYasc2eNa1yMG
twZD47dwMJuViOsTP3NZQgHOlIKV6Cu1pYquqV1TLnbe79O7XHdaDy5CizZhI94hcHJpzEp/a5hA
hHiAnw0Q0cWp391cKvgqoWN3gFCv2y0tydMRdy3LAHIplyNaov0V5dHzZ+EqTVTrlQRBsz8Ve6nL
ogckaW5etN+apgFzz2gQc3sMFjfxrb+/BKN3EjLLkrGoq3q5kZnbD6MRWhQkLLwyzaxaP8/OwZHt
8593KXZMD3iHp2qul5wlGkbNca8DGFCyM2TkRtC51px26fnCyA9+FDDXlOwbKKX69d21U5CkVk/8
MfNSyC19zUin+yPmL/C6xmm0UmbjHoxdr3+TuELvTopXNAiahxzHrYC2ZyPlOJr5YyyloOajwyFj
/bYkP6NAHZZu0OiSY0/x/g4PbfEhJxlxnZmMKgCQusGFaRYrecz2BVQb7SOM9mo81hb035xbWWBZ
S3cgpG2AwCK9A9R3LpiVCeRBB4/1PHzWIFZ/VTW/HqA15qVM6Aq78l7JjYe3rSjNAES34RaD2Fzs
QjWwixV8opc8dlZJtiVrDeQZYd35e7o3KJ5AJy/SFzk+CPyImUAOTxvbtO47U/L7tM7ESW2Tnu2O
59ILgoRFX252leIiPFpgLZ42BZenN7wZQBnUhtg2dP2Nu/JGeF/QUwEHZOveQrza8f56yRHNXAIm
mNmDDBg+uOQBSU55IvXkJOwm6pAMb15K31HNyy+R2GpJKiRrs2HbvHebUHrej+Fdm8C7/4cuXs+d
FOS4uc7sq3VpuAqhLk3z4hRrfc2MTUMH0Shl8UytdNAl0txfvWdzt4JbL47zZdEeOIOSxOS3EKgq
KM2l0WPjdQt7Eyu0ygvKJlbeZBf6wwYpT9St13Sjk3+S5oO2+rNwJJgYUy3do7A+d9Y2kEBUWm3K
UPgi+0z6cr+r62SeIdkn4lPwrbJ7EwWqIKcwFl0PjwE+XuxzyKlTuq05FY0vmwSdHTbo1nLhEE8B
1KcUqVmCj/9g6CYj/G0tMdgsT3obImf/SeXzOxkEw3Z5w3amgcNcW3z6TUDrrcL1V5Jfxs91/WEk
Spdljqdl4gc5RQWbwGf3IHub5xPNmo/VwOuexh+3tkegkUZQ5IjmUJJ1naSWnqg/IUW15kJslAui
Jls5UfNVVM9pYgepP9OGnK7fUUIT3RMp8sA5mkJU/7dy3rsNDSH2JnoF94+3rZeLkLoDkpmYwtDm
1mDFvo4MA/CQx2j99yzVlNRgM/4zHCoMC5DIrgkDnOHjguRCGeTWW1gt/ufaSAMiTd/iS1t32Ybi
UB6bZZcFaJp9Wx6+DjagxkjxoCpPnMjbCEBIDb2IUn2puM6tqjXffsoY9Ohyj0z9Cyl5YQuw9kbQ
NFrVCtTWnSrNBcnmOBTOXPUvGnslSFWXOweMa4vKw7rxofhEGaM88vxNy57Aq5vuNv56ssMNUBLn
9M79biZdSi9V7DltkHitKBmZ8XU/analL1Go9jxiz1spmGoY7LowdgG1SBwZ0eN3RM7ES78R+PJo
uPDbenpSPHgW1pihOjF2tb6pQYWxG2VXSr8M3gXSgXjt6xRRiVH9DD7EEJYIYD/h+XHh/Ds79MrE
bM7CwR5hRhozvwhQ/dcmHZEuQq2fKg2IDGZYU+jgtGK61eLi+UAoEo5z+ppoPJulnSoOCs+K4r/f
vwHXjJ8KkJ1vYGB9MWS5gJU0ZUwO58sB6lEEhIXu1ZYSh7SCNtAt/XsEOdezRPq43AgMBMKwdR4b
Fer032GX44ctYnlvlsO8gt5JRmDwyCqlDex1sqFRm1dBYuelVW9wwg9x6VM9HvuRI7QXyvQ75u9Z
2jIali+pgflO0zwmDeLeWtrSN1mfoHwQLf1PQ/UbIrBmPiasAkoSvRsTj8wU8DprrZqGmFNFNP2G
buYkScA/50aqTRhi1n67ZJoG3UGRamtyM9DNyGQploQMdHhhQjAwOccMD0qj06XQECaWcyc/1KZB
HfQAPf5U/pQwi03dziMmUOhsaQSQ1DkIDLCzfhHVYpGqTPgHcYGmvv27X8tg4y3FdRONMpkA4jUp
SIRWNhq1yXecV9eoAQdKIJ0e4kY4m7db+88y5nL6nK9bc/zOHv1OztGCCplAtvhgMmjhjrqarPYM
O8jb1VjFlDfHrJwYlmiVhpH+b2nlIW1Lrak4dOCmjT60kEPEAj3Ce9dZaKw+LHo5QkwjlNXXtlFH
AWA4wtLOWWX698x3IZSRaHeuN2nkvbQOep70Xt6b9Ib0QHd9OZQlwXprqF9KlajSTvg8zDj0LfEJ
cp79qIy2kyS/a+Q9QGsatdLhG4BRt7HB4nA3OwI7DM8FdmvUqtdOBOm8uVcGrjAI7HC+dP1R/sgB
D6fxv8gs5LfpOLQTzOJEYA0o5yhDHZJTxBxH22KuPsXNFiXdTdoJq76btJiz4dcDdD+usScTvo8p
ASmlx1LFsIlZ6JUP/ZMMcV9d7BmLBbfNvoODK5qzwbgKw1kWNvZXq7Ujr4IP2TZ4+nG0O+n1s2zk
rq2Fmk6B9rKdMxjKAIDX/nPdgLAcvGmFFIfdOtfdev2Prpqv7MRzBhahrt4bX4L2B0XjyBqj6XEy
AeBe1ST0DSHaIMMcbKtO9Ft9n1g5haXtSJN3fRQQdqXFsm5ZDb6+VbnjNOQbEQqhXEcO2Okd3jro
lFiit1cjdiB8O3qJ8DtR36o+WMNWMnUJGvFvewJlW+DiJw5upIRjRpMABOkyl9FC4j/0o0OeI/KL
WcXncLzTrdrgmFqHl1pmFTH0olmcI2yGqgYIhBmaOToH9631+m8EIeI6ZTucq07kIaE+02mGGBnY
4ZkxMyhlobggY8RzhO7HhFIe+ysGDPe9fCkDLPDqMy/0rv4B4P/QTX9IwG2F5jONNo8pmN8+b6bi
eg2T8nbmPaqe3QpfXJXKm3XuvF5OP+7++jveDASY7xSJ0kDZli2MxuWbf9JfBNl0Y7gLcf9IkilC
czZI0nUuqNTFbv8dOUcuy1YcKIQVNDG5Dq/8BIlf16RI6Te7WQtrwMWx9D+6XXYN8nildsRNw4R3
THQHyWvxP5zoCzcpOtcr5xgYqwfjqs6xWgjfTMppmIU+Ex7HNsiUMAv+EAw1cN8FhhWjcDRnejnH
8arrPD5fT5b2Ejg6BsuMFp8QCPAzTb3QI3sRlAaGjIaoEd/nvL1zRtc7o9uCYC046U0GmVrf7oTT
h+M1wie9XubJO25d6sW7XjCLPzKlAdpqMd9dFRTaR6FDf0557g16ss2L9GxEzQ30xlaX4asARZa1
QvI1JG4XnAZ/LERbdXgSrP9TKZMd2TPkd5GhKfBNbGDiMkZYb00D0zCDc8h2KAa1ypmW3G5Du0rJ
Q7+736W9sWIVQoXXGH2qacyHkc9gbg7XDb5Hfnok6KDneLVPLxlfli6DE0oImubuzZjBrwgZmrnz
e/ryjqCu1dVdiUYR2wXmXehLCbRtmmhTGdo1GTQt7S5id8i886teggNl/p3mScjEqfTtK2F4b+lU
ylBCvA6JP9fLjmxCXcbc1TuUNQWS09r1aXE+qJDnMriGk5qt6DqecaA6Uh9+OVxgkyNN12kcsb6S
LGSLNKfkm7wCZlUkgzSEXyyTaH5Fi/ECoH4xwTtM0dRnincmfjBIzZ9FE9xWJIc5EOXanlYYYgBJ
OY0yQeESNWotlWk6HL2+yDDSbLbo397OfMjP9fpmjhQZIos/7EJXYHQXRKcI0BffqgGpIICxpDKA
Omdi3Q8gXA46oDcTPWJnOnQZN7wjYqptC/e0J824IcahoW67C4F7nfh+ZkwItgr/2bgvJ9MdCPDy
hbts/5eA2PR/ENZVszTVjQxxoSDg/XtvYKzVxmAIYjgQlZPZPZl9cfJqJXsAm47DiqK2FfN47Av7
Wsjy1ejgBbHOBGFIamNgq2VuJOFTKHIguAU5d9tWngA7z+GI9buAsQTt0ScCe/4vZ7IJiFsFyAeF
MLjTOs9H8xd4solB7tvpM3J9VtGbiy6l859M/J/gPUGInaV0mpS2Zs7sUc91Tcrkue0HkVCCpvlV
zzDwx65qj1vArAFOX8Os4d5I+tJ60iiUhfVBfIBeU/8BsyeBipKbfRG0B0HqWZe9KSdOzRGrX4R1
WnOeWvUU0dLRsHQfLR0kzZrN9it321/YguvkvFih9Md5Voarv3FEf6eITxOSi0u716vpoHqXl2cv
5qHnd2zI99uJJqiK1Gd1waSwEYAgtqOuV6xYOuwYXukAK8pxptItSuFtw1FLiB9Td2eO+h1esny5
ajkqbrdW3gYeccHSeyZd/7SzFbOXdwT+DIMS30PM2oVVg+7PCWt2AgsEi5Hx3ehg97L8jmtzORzA
+dE18fq3o8FZC88Q88jCT+xVxxtYGpEdok+VCQuap2qrYoiGd/F+xtY8ClBJZga+pXjxeEUJ3O2K
O0RYfOLjX2goXnsq4TfCEqND6KTH/LD+vS8ZsxcOGCo1Cb/wuywq94ICbuja0oR1CAmfx3KsUPa5
Mh5U0duJR9/gDbl+rbkKfy4k5z4d+TzWTw1UJsriUGvOiuf8NfIVOdLeCm1X+gQJYM7Qtmlzt1qf
/tZaVY6+O1XDJrMJHuX+0KxcFkjmq/HE3Ni0Y3cvbtLay1h3DCi8ethLmzZyDYGnjSEWEQ6imBwn
b7x+0gyz+NAh+I/9ZslWMZzQh83aZqc+giDrJApzFESjGJ4mHL4oV2b5TOyABJCB15ZubxSY+ifr
1RqpCJSF6MmjExS9UXb8K5zvgj45Vt+8IqTf4NUwPA87Lb9Zkaka0rLcQWnWIXAWmpOV/uTKstOn
DEuK0s3xXFcaFQJdi4OiqaY5DN/nYiuI5D+STuOj36EdPynmQqvXP78J0fp6aIiTkWrhhMTk9S7w
9ey3hKaiafya0FMq4D+Z4ERTMiqEFXjG24lcwXyOWfggJb75C6bjbt6W6j6MZe/yuY5hN0Kt3A0P
PLNSNXq0EvlJJ+04tP8ZXt3USu8SQeODdaOTN1NhsQ0O5/jfMine3HnF7lWFpAHRTLPX7728Fg5s
ZaqKBtWuDohTqPbZ3rEzexi8FQEyXuXdbQkkCJ8Q8BT5AsL7nSQD865E7oA0YSsFJoSLQ5mhEzSO
4MnRLX5NNNWMqIiDeUBDGbyxnrDrN6L27dQ8/8DySXQCYTD9t576sI4yaI+Fdw1zp9t6dVsdskCX
kit0+3h+DWUM7nB3PMj4Zj7ycbnosZGfCwn3w+lDh+cI2NMbgU7pXAm5x1JwQq/i06nZdbMOcQyM
YF/8s2ObVb9/WS5YTL7a4KRgbtLZVggrneIU7W6TlSankY+z5kCG3gE/VtU69nqKkvHXznZw792f
kYQck8iHUKWYyUTDKqVTdY9RYTAiF1RF8SUC3OBhlJ0BNkoB75yKc5hRg9tWUwCSXEDJAK/vdqFt
Um1KNcKCIbw9pV5BLVvtJC3RQHFKya8vQmjlzIop8t3gTJy+FHBbi88LVYvh0ZSwb/T0IhyO9DHd
EYDtA2aZDrk021+DWKNLDJCAJI0YkcYRRv3maFrQEXeHAfqiHH7BogKCAnLpgJUEeAoPqyJvvIzZ
CHKgqe2/dLg0CeFULpH9Bz5q/b1wc9fB+zEZnVPgwQE9o2tuVA319psivqBxmTh9HdJIeWuFXqAd
DMnofq2HHJ2hIwhOYodkWf2UwXsc7QWMl0rcREZHbNqjUmAJsAeCxJJ+Xlc5VuUEUpJVLa7onJyn
z/qKnmJao2kQP0C1Ep1ULpeXpos6vUs7gBKJUOr5j18B/Npsbgo1tqWg9D8biiMIn92v/AmTQuId
vHt/AYWflBscNeyWT0ZUXXpKNDj+HIekUZwLPK8uNlhPMeAZjaykCo2Xu0DNL+zF1Y6dZdvXU1tG
NGdJIs5dR+9gXXXHwUHAXyAs1RGzFMuBHFkuBXmXDC/gawrCorJXRUbSqYSez7kr9O4Uq+J6pUYY
20cbYQ3wjLZc9L1M/XCAp5k1CNI8yvZrQ/F7Dl7Uu0rnMxggTpL65rTLoXI0KBaJbe6GmjMxHILZ
Esth5Afbk8gNLadYliZo5P7e1Tu36bQ7m8cCRtpywjkH043Qk7wVxJyWsuGjbMEjfBTQk1CS1/dh
6Pp9K3gTGzmV2crd6lff17t+NVEWBI2YkqR6nC7JUDv2qcBP0UNL0PeAXqy5DI7sMwenY7zAH0uc
sW/HFHpQ9y3deCN0NgKgqkceMaefkCC1UpvM3mAIk5WWBhr7JERDuQLAA71tnyurnT/LV/u8VHCX
CXlErsfc6uZio507/xQqbozbU749U4GpC/vWQa1E20VvOqViSAq3dyv/g+0ENqe3YSKGPa0CKs9k
H9sPhd6J9IdMVuYHbYRGktFCE4zUTbQyP7+MPZM16TtrIeoGzOrR7fV8nyRD6xKfeQpqzevl+Jfy
h3WUya5RjGinXhtwLT3f/mko4Vg7l7KxzM1Av205L44BPe/6tcACqsLFx6AsI85LaAg/ULEJqi5S
Qh8ueZAcyuPH6Ad8INenloZGO5YyLU+8L8NnX1Cun1AwK0Hh1drLjephPhNZ1MErDBBXk8EPtFyd
25852sO+kF3CRXHDLrIg9QD+01n/oUFSf9JB/I+uhoW0isClEKZqu+mt+wNfyzDxOHji4AL4ok1/
sEayM5BdRSwtmRbIlmivXOXCtIZzX3eR2rPxFi74gBnpEE9Aeq7IkWUCzVRqj0ubtH3521MtVSq+
UD90YULMAtA9wfwL0hSgF3kC9zDKRk9uyNYHAuLaSW2bgEmsWSEjcMjNgnFmD7xNt8nwXJd79G2w
KCSnchJDvVWxn8qs0b3VAx0GjH+Vd3/FBrfWPJxRAaKxrdLAnYAK/ujzVppsRJwqhdIKEH2iA9tg
ck5OrURaz6SolpGGgsHNICJSzIWdiBPlLHxs6u2BtcpGWyC1EbcFEfHBoxbcWcFHpneZWMBV+SdQ
W4ub/3jSiDtgjzivYEcOQo/1vxdBJ/VHhG/ydeDfZ4lLK2z6oXNhTe/YIXmUmcDBa8kRiA8+l3PB
ORLU5hnVuCrx8Vb+zZuYUdGhiyqbmRY/X7QW7pq5BxcTG/P5P+XSp/Hi17qjDhIsUP8MLvz1/rpg
+rC9G717yRxxSvPNOqbV3fkc85LjTmvU7X0umR6+etgzqtLW3JQMNm27UHpCm1Dw9kyIgvXkZV28
G/xAAvmPHfd6DXNsHGqUtXcCD/n9TLLdk+tB3YxnI9EPPilvB3lpYoNTFubynWdkM/blpAVtIhuw
xYq3XBNGz9oJcaIuo6ASCY1OVAVot45gvki6Y8c4l2RDprpily1OMwvBiPR27HnnBHkalUxK4W2T
HnQqNDkn94cgMC7M+RfRe4jMnTf9VvTAJZflDvKfUC+jyAlBOQJ84SqeH2vgcEF6zStELZHlF8fD
qmR0Dtdebdft5wb6Ne7BBTetjb6baA3ayvtkB1C6iZVW0npkK+E2ckGxNu4NO6095Ufnx/Uw9c1o
RuJLZWelearZ5Sk5+eeJJuQCfsLpUsDRqShMa+UAcKhcXDVE14Q19wHYuZuI8Y8x247yfONFejtM
hTf9MpZVyeufwPYmxTSa/dHcQqSZe+QYLy2RVNqCozWNWe7NI4H1MYRjVv0BC82sCx2oO5B6QV8t
yeTOZnfgkxLXXglhUvMJtMcUSgLMh4+k245B3owkE+78YpNC7NbByzoZHAYnCaqBqHq7s4i+wy3A
ILypydVO7wPecFsiUad9lvjO69KM6imFjCXASLLBb9FyGlttmBDWLYCLxVwVFosypIN2xoSQlKFr
PLmhfRSUnEA/qFlAXMAIS+yBBKhoH2IwTqrW7+MqBxSxkdVjpDNiMV4uPs/CDSIM79tlgwz8OToC
VRzSquwW1VlqdO4IHpYyulqtfO6MOgKKAI41jfytxMZtUbTGPzW8EE+HNEHXE/gnVmTZyvBViM+s
gNQXTQ2QCLT+87W9ZgehMa29WkpTnlwXysYbqXrqtONvJtYmaS3O6xPm1y7FqMRqwBTsya5umDB9
isLzPzJe4ntZB/h2sBfDQICfVgQsXa/i+NomwD6yNv/O3Y+O2psvvJQ3Kbdu795aoaKvAWQRHMud
G1XpIWmN7uDFuNcpACI7/g3BjkLJvFuxiZNQJjL9Vqi17X9WfBLQaRrsXt6UAe2BYIEYQCOAoEKQ
EDxqBAQBHe8G0DkF3Tx+EUWOK/nVA8rEY5QUUXyMTqpPYbxEk8MMZkrigLeuH2qSzvQBNm3i3PkF
nEtyVO6S7rOmc9j+xmuS/fWXDHy9QUfF7PCEBeaCBVozSWWA80NUo9iI4nDW0CJWs3UH/aT/2d4I
JkNQKZsguKBhYyZZwLjjiW2xVKaWl+KephUAsVP6ogOuB/8Ai/2yrSmAmI9r7Lvwejb6mounNnqD
2AoFIKmd0Mhkiqc+gLT4q5ASiZkrws4qejJQSHFNRLSUZMc3AMfAdInjLqJZ1IEyeqjXuh/dTlJy
VsnhEAB/GRqL/8lbZKCiuZ8ZhCH0NuJn60wtDTAUCZFHm+7WMcm20Di3OJ48jcxBSQqeNW7DaL3W
2by9pIXhU7GyBXRuvk1uuZtSGI5haPfcsPnStn2vgrbOog3Mtp1k0mDQgEFJqhiGqi1VxPYJ2Kvo
0tPV3G3KuFyyqWMklAhwqXupLRayvLb5vDar4eNbIYlJQcmvLyajS0yJ5bTNLOB/wwEOTcHhhM8c
p9VVIa3t2JHKgwXtAdoszKhnGsqGlI5ONhW5HAq129zUUiEvMLB1vWBExix3VliOzPJuBjjVs2qZ
gRrnhgsJmlvoux1VtJKsFe7bGuJg+CbzBrFjRxpO20eDMKgaps3+S/Bu4WmSLoFkcNHEXmoLFwSw
Ik5Ma7EYdJ9HS4q6qtm4d7ji9DGqQ6xJ0yss6Wm9nxaljUTHyOta/fO0RB9+xgvHP7jYC0HIIOop
bmKbAfO4R6hWfTGXLMW1+FACz1rjwJobDoXoqLjF2DAwHL2VUP0d1eMkKPdtmvy/lnEadpCAW4UT
Zhd5v+O2zViI2kV5TdB1syR8NAzOnG85PZxZeNFAK6gRZoVXZ/0YFToeLEwCIoU9BcHoKAH1kA1A
us6dTb4d7A6vootcoCBDB9jFc+EOMaYEvHK4iXaYgVKyxj10wfb+jXaCyBOw3I0R2z0COTzwantz
VSy4HgCP0UdWXnDGdLmKs5kR8MHGCITpA9LgTvqLyftVGROMKL9xWSTDK3pbFyx38olrAKoskLkV
UG3ceVCqO/R8tjXKopIhgMZcbJkKVDuzlNZD0OZ1jJIu9cuZAT36nk01merN5/Ns9WmfWyM/5rQN
bAc/1o9yjJ8CoL5iyt7TpX4AB3kvGDqzgm1n8yfk4f1aOUi23aBEJ9toFNo/wcdHh017MQZCICyG
vBoIZ4GKapgFbPUervDgDjFvkleLKJDbdNfaDemLFLbEGpzeoc4LYm+6jYay4Wb1fj7NfXPxQKJN
6N21LKmhga4HpXFzwcnTZ1nfPiI7c1kCVvpGRBjxgkMgtMt9d8UFqyyMTwv88PFZ/cgDmWilmwMO
3L6S/szLboJE5nqnyp7S9vSBIUoBM/0cLURDlGNHFSXi8OBTdbu4Bxny8oX8J+enAWv+SF5hEFWl
onlxuB9VUWqYT0llV0axdtLkAjdTLax5lIRFnfXgHR1X89JTYsXR0JGjxwq59v1WiA8TyraX6DUZ
c2U7Z+irGyoitQccBBxGGeLv68v7ijwGGcVBA9r2PnKxUI9TaptCw8OS8xzh5gyM31wpPdgssM7X
5+QEeFtXMtMN2/9E/oDC1f00iMej1g5Ev2dxdcwWSRlOT9bCicKaiIdblb1UYfsnTWsBF9RL66Sk
R2ZMZ263uVtOZW1qrLf4/IXUSGMc+M1YYX+2ppRnyfhYei6j+L2BJfHdEm1Cj71lu5DGUo2CxfTI
SIjdImHsbwmlhWqsVOrY4uepSpoYo2NH7EISYsQVgnEBdboaFO72LhRFAGHRzm65eSaxfmScatkU
DPcSAg8+EukAwwmRhocgyk+vtH1L3EG/KbK0SfSE4J25s0mxDVO5lypR6CnZC+KjqQDkL7IIiN8G
le9wfFsgT0HBluxP+lRTpSI/aoS93vrscZxd/Sqfl1G0HXe5ZdQ85DVjekNgzEdfdKZjcgS/gmCA
cHVlCCJSQaeZSEDxYxMuIp1Rmevv9hgaG0YsGPNW5sarqd/HL7AInqbcvNIn/B2SZeoOu772Bp5O
2OmyAIB9khapbVkRYldTa68dF6cBehQi1OBkAIb0xr+GFZ4Glz0YZbRqcPd9peH80oGM6SwMW++I
/QKnvhGVubCH3JBqxWyOZpuBdcvu/7xNj1wwaMts3e0PubM6cp99ADUjLmb7Xeaw88DF9XM8HxbF
ial8VVqfW07Dgfybphb42/RmR/YJP8VkrjhmLLzRezLabr6zJRNo8lIPC+VOYUr4rALUZzXPbtzg
5S9d1kAzYUhRQZ0XOBdXjZF3XB4DvmW4dO1g6Ec5FwlXxs638hGgPO0bd3Cla8Kb84Sn7VCalzQh
moFkRHEENDjMHxAU0p8Fiv8D6daIyxcotxvyFfZfXSl8z86w3/4xeGDydermK9qZMtcp8H98CwB7
HjlSUPF6PfSaGPHIdQZYTukVP+Fp4+7cqoUeD+r9x8I3MHSvJSPjUq/O1V6tlge4PAevMKOXOLrO
dRy0BDV8/SN+BUh7ogGZUr0tnCQ2iS+R+CgfPEw2oA8CosasEVo4qdrHX3F5O2wUZ2CARBEPJHG8
32ymC4nX8NTNj8Pc6ZRoX/uMzCpbWUYqXojXNNcMh4S0TNN94V95nfb8+TJVC4RGZhYx91CLze2k
MFPJNS8+x0JXhQafUiMkDByHUxk8vmxCYRjUvOqBwDBi/lEzBs5ViyvDzaPiKLLbxIA4E7Lrgv8Y
q8v0DQWMP4MTiynwJYJ2RFLp2W7RADRT9YxKMHAjQwW/gNUCQwJTKzcsYJ5ouGbkui/BHVm6ekdU
QOX8MSWxoB5MUcaSzZM7JvrMeG50RYTzEoREs1/vQARWD1VwdQK1ec/ntFkILEkbiaiObLTNIaKA
6u2rBpba2hOC0xBqdObSmTEcwI9/60pIe8lJ4T2rgFyUCoeBQ4tgnOY3VEyv7E8ZwX6ylBCWxEK8
W8ks62eD02oDFUazdqXegcn8IsAAw6+XMShXUb45WscX7+dssCBxZtMZGGuwNHNXpeTY10sXIMAY
h1HLZukjq7HEJuCFZsW7YeNd2sB1VRaUgO+4FGro/XLTzCmkj2w5kMBe0uj3qkMPudBGd4CN87vl
kXjNsXG6Rt0XG6IBKI1SXOgu+sfx1KMrDPJN7DxtFcMMcu5GpwWgfdLyuO1d+pKKQkfkyUpzp/4+
TsoaVuUPnWNEsZUVXTEwobf2TpRYDmTrSzaPw1fpKeqea4vWzvVFd+NR06OPJfdU0jjYYvisA7OG
U9/kITkqfsXOsMbTTWgy30xdi1YNkXB2lXj1SvypqwIiZRJhqDcdkMCT1zWoiFYBOENkd5xiHRsm
75ESFlLgHUPxkdSwUuUUPu9li4O5sTwdf6xISrSBT+YK+Jcki0bGpr7YEmA1f9gTGMZKhq7IlurN
kWLqoeNMN+FCUV0ljbzWHg+D0lwMkWROH0+guV3VIzpvIm3dmWgkjHlH3dKh5A+oUAtCPFcjXV+L
/jsZz9/utRDzo9gqpEQFHVey5Lff8vUxiwW3+P5vPVtqy1X44ABTE/+TcXZQlAyZhrDrpWBWsi9b
NcQOJh9Rq3cSW3NcJy2n7tLL/wQ1Wt6LKIpX0Ip+xPFkxlBWvS8FdFa8lyboaqsTFR56B6HAf8Fz
t4ugVXflWviXdcfzjlryLM6fRr2fvsP4KIy0tqYiwFZ0Ci9bQzorYtZfz2jTa6N2ejX1AXtSfxFP
vkCX3VrscwgLufbClFEUWlpFAnC+LKLZxairgGtZ+mEwZVXp5lD50fXIaj3KAB5oYI8ZcXxi4f7K
ZpueVXfQt6FDmDTY6jgfeiDeh8HuqKZmijSP5eCwYMJPHjfR4/ILooq67AlbeEp+9v/grSfAZpeC
TpApSKXaB7D//CWRzAh11Uw+xSB3OmN0dV5Pd5E38xlXQVYssOr1h9k0EH3B33SWGp195Wa1ODjk
1X15sconI+iJVONpvG6bP7Snu4/1hERvNrrVLDLeVtA7OhEu3h0SQGtTLCeIQnGOoU4Dai/QB7FO
9v3+FVqas5vwreDsj8tTiQkPI2jFPkHd+SoWfHQLbCxY8NNq3Nz9abxZ8DS06GsIDixC4f+DgrVk
a//pjUHbeoUiMnMkTP1nbPyWXOLHYR5PZVw5fRnF17AYoETi9THTclk2UgUxvPK3/SfVe73iOFmt
7MAEBtXEfWXKZv45P3G4wS3XUvGLEAAJ6XXZlT0tRSlRcEu48gfU5VePovDSaKUMH0/mWXGFc0jo
RG+j3FAR87PPDK2QCq1PEuyHPUIL7yDf3S9h/Q+2Y4JyaCae7dy2kY3HHEIaxvtqBy02mV6z/s7h
ROtEd15dS5TEOuL7rygnBWQvj7wCmNUioZcn7+jqTm3/mTlZBNTbIdhlpx/sF1j+kFmQcoVIvG0m
xnk7BeoT2O8kbQ//0JCcifkrMeuICWahVC3HLicANuaN7PhWmvy0MT8+exjWXsEO8jB8yy6vFOq6
hAuW9282dxTayqw9DCZgtPaofhXlCEY06AEhqPBK2j7d/JUux7WRZ1Gqq3whXI/dCGeqw7ZL05nZ
+YovaIjUDkoEcdVjnfmGaLQcCvsQHIxBsD5AAeWAAU+tUnANyPd29E/XdfjRj6Dg4gHuqjJr5cH9
k+wqpJHBYQA8gxnSJ/xT/IAOrvqGamqQIofJQpE0J38B81OHW9cL8ReU8vQggRAAX29PozPYn2nf
KtGS1uZ1Z/Sefe0AmVTDiXD0anNVenHEResCKLK2gbJYywuIG8mWtXOckWjYct8TdefvYCUBaLEZ
ejgew19mZoYkTaVw2mj3bCqQHvxnoIFYU0LJW31Zdy6caG9Dgylm+adW+XnOYL6oKBkEAuPkuvOV
bE/OhnS3QPNrZZXVXr1pvUP3X3IqqNEC3wJHOiGKUWjDjFqCiMm+zInQ7jKYQgN03spKtSxqxJXm
qPcoHPDIDDx1ZW/K82r8OQSvDinB5V6YnGf6/qp97+RlU8Do6q7M5q8KbzF9ARhVGIAP0UlJbhcI
EQmzwwsfL2+dgY11bo942gp4E6IR26MH0Q7xhd/04EAVi9Q9WXEucDIL/LXipBkGT8btmGEHkt/t
T1y2rzgnKQfQ1EEtR6C8JRF1F7ihxzZQQ9sI6PCsX/S4jGSEuxAE/QwJPBXoftS1UKoUlGlJcQo3
EYsxNyVlHw1cvf5tFVUAt4n/KPwrZUxsAWeknYAniTL2VVw1nsSmt0Ix4pMHrMdIe2HRMQpBgL3J
bRGUxZD7AlnD/DUWc8yGefTSIMHhl+SqxWu8nBcBuIskT30dw7oYd2UJKDYpCKUjaoM2l2yrXgAf
iEovYRbSMHCyYdd+KcfSnWxePgUEJV0WcMYfobzfhDElj9JSqFBjZOq3DKsMMjqGN0dOP142kJEM
8w0VeK8rnAIivCALEQp6B0tA7vqtU46nItFsakdaZ0yBVnKzJ/gTx5ySHIjs3dVatyWh/9Fbl2fx
qFugCftkjAptAAGXKLgeFXw1pIdLu4zbgobPxyR1ZAcWJrd/o+zH3+GHtNAHzCO53DBYKF76s6oG
k/PWwp2r9kk3JNpawCcSR7IXR1rwCAL2u5L7sdtniZk1zygez38HqpuAVRlQHjcjqVlyRw9KqXvs
SZ6wSgoRwAsH23Du4owkmdsI1Ya7JHm7OmaJuxn/eQ/btn9rJok9fNE1RkLHKsrsl4wDwGoReWiS
Y/6570Qxw5tGqxnPxbWmY4Py/+YERCSY26lAAPOpviEIvdvkSjAfBcBnrIj64XDWV2KzanFG9fPb
3uuv7v8SBpfXS5c6cfrapHh4Ch7WGiVVfDYrTXfFKnrrnF4bj48/JFwtg9lXdlZu35Yz+Etb1Fcf
FqB1OwhGcE19KYZKepRwoSXPw9RG1EGXeW3Wfn4epd3w050/LnFN4sXZ+bivHw3yBXckpEYoCLNd
o3FUcx28jXRaMLR62alm0TWFTC0JsrrVN9TEOMnZgkQYBRZP5pr+yXZXJSJqY9bt+U0/ZdGwnVcp
3hv2vdVonX8VAsAW8QSx0xrxvfQZc+hrZtk2dwy0GLD6IZ5UdgxhT8ucl8xptLm0u1JxdOogkmkO
i2+NqbrgOwaHd6wDqP4DQCD3nNJXgQZgepyuU0asDQHafs49CseN9h4VS2Ogd3VFTX0ZMJu5b2ZP
0BzU+pAtttV4QPr4s0/qpnRh48BL8ErNkBmgf0AqBDeuwhjLN9N5QZr/rcH4rwwuokUlQzuZjwL4
ORgyh9kcXXyd83YvDXWxGdZYG1LfRj2Of1QVLjG961L8yIwYXyAiwcQeJk5I0mzgt0lBNVVk6xsd
7Uvk1YpqBOeQJUlGTOQGmXo+ozyatEV5ohMKDqI+hkPoAv2NoIKrm+rdRHZ/JD0q7omn3prWVTeA
cGjZOMLdg68hEaif2kK0yixLEXD2N0w4pfgp+8rGXz9LlJolC+cWu89H2Jz9q3dXo5XLhKuZnewF
N6zhguI9OL0En26IcG37d2C5dCbfcdeGKQ3gwA6g2RCk2SeeqRWSM2UO7JRp/RymQVFDx/ZniX8x
GVtPw19lSfipObTWeMfXvssSOo2SOBk0fdYodKVGTL/0xwyrOxnZASoaGrlbwksA5ahB3i2VUydS
rjPwavrHnYCGSitqrXW4197SHeOrhJsY3Xp7qGnDmLCLbc1atDbWSbr/0eAuhwMa+3R2uO9k2kUU
ERIlQ2zBlBIBQsQGKVetUqemYHhRqG+ZPtwRzs4FG2pyVe7F/vvTfVWEzAi3hd7e0usLim5wuK5c
KaA9y8rwGxnuzNmrd7vOKtIbjbR/n0XUx7SSGUCXNo3Em/0quvWpF6zZ4NGTP2jcvLtNbcjjqE6M
/j+4n9w8b3mE+g4VVcygME3g+MrlSZklmwajnPbUh2OOBikh6bzkj6hLE8kO8OTC9uqVQluspL3X
Rddt2cJjL9l/604LyIes9x8cIJD2DKUvwut6Rb9E1dNpG1+VrNyQ/Um+gyi+MmZUAiIbared64bF
+b+y5MQjUDuNZtwRptAjwuBS+EqdIovhF38AAWlzV603vgKegMiDdOdlt71kZ0p3lZ8yw+FXDOJ8
2gFBgJkpu6P5hhCqfydvmO1stygYfgRU5jQGBApCf6P0ydIlGPJoJxWe+vBvEXIuagWz5AZNuDFX
3jd+ak8avni3EB/qbXz/OSd4nvwu5nPEwQXj08Y4jtShDgJgD2FjNvqjw3SupQC7zaon5EWqkQrk
rrjwi7I1R93mF4HNvV+r2IfKQqWaj7XJVA7sM383HIrm7JfTCzOKzqStxsHHcJgfSxAcnPHEpaoI
fCeqm19WVGZsIDlC/OFNtzbKnztxVo17f6kTYlvfEX9npUENLOeNFVTU3LEXQlrGZ+D2MXs4C9uJ
RZh/Z7gCJwlu9zg5Eo5ucLIg0FuPEz+MO4FcjdCqRC5mgAg+hWxvM8fZ2zZvQROjMSjvKO8vQQmB
YsXEYOhToIlQVAa4iipHNB1064EVi4h/Iv3+ZCTjHXVLno81obZAbt6Km9BcBZYmTkPD4MsjJt6F
hX5i67kl7Hv9rOzsPb9zybx96wTAHJB+V8NsC/iQg/K8pu799rXSlZFV+kj2mjF88DLiXtlQhE/5
lBt7FhDRwPqmGQqXfcN9n5ScvW+yUHGePR1Y8cPocUzkH3Hb+3ZPgt12oxDN3WpZ5WQLQ3ErRl2Z
7gkjpMCot7PpoYI3+etRBNG/pskG+uyPYfKo46F1fs3wY5xvj0rpX3Bh/LhntgsbNDZx1ZrmjW/7
Tb98Le/p3AQ+j3OfqvfzM2K6TzbnkNA458xsn67tLvX5t+rEAr708jKqVb2E7FgT6Si/aZVh3KqZ
jYEDm5B3GQDhmYOUq4HNpc/1UB6uYJtYhdSz2aZEMJKZ/gYH+u5jLjItE4w4Flu+mvGjkWaltAAx
/NZGTQXx5QV1Xdom74irBNHwDa4/KXmhj6LrjexcX1ge9g/ZPXPeaq95/+cbjPEv1ZjodQybmEPW
x/KOzAPTTiG2vjMT8p6Q+FEA4aGPzsa4paZm0wHWI9xFu7OZUKb7sK0/3TRlq04vqmmxwG4p46Ya
OMs1qqDo804dEKgUQ81sQL/qqLmqmd8HhRqyplLlCCEHgP76Ng7TCeAeLEgUbw9aS8V+dKlfiutN
DD/1PYNc/9Mssa8tc1c6yS144AC65BRnN2jYatozSxFrIVHjrUG+/X5FJf5e8OaGZ7E+LCpbip3i
6oF0X9owXCRTyK1ASFDgsVYnilmfkbeun/U6c5D6ERTXItNGX0RzojMWD1OjpxTsbP4MT3QUgADU
7q3hj68KzVYBEjOQ0aDiNPcAbU7xBNB2K6Djm3g0rDAulhMLcc3jRglt4Bd1nUX7eF+lKWTKiwlh
4vEYTYkYvu0UE4xoXWLfWPYlW6m2Asv874yc308Fij10bSvHhYoZJPcj65OIbYhV9rUUGSh944WP
7WhNIfOcPFpS5xH/2g81x9MqTjXDCywpXVkuC5vllGuino4GhB8yf0NWTv6ZJ7LZLS0oBcAVvqdb
yj1wx/NPpnSFrL2DVCuVWULvNEvTGM/+uhfuQNdh3XM1PCzQpn8YdkcMv9tWVomW9p2pYqkTyWTj
MaA99TNtjzwveeFk8X8t2fp/t5c++o7vMWPPaYtyL67IDGt3pdZxjgnCIaI7Vle7lDFPw1rOBExc
BCGX2UcjjSHFgCc2IYW8kfGASzPMpdJGJQ1bF1vpK6uhoN56OusGs6cnM/YEjNCsmE6RjTvgnjY/
URL74Fm6qrDSxWAm8iwDD4Yc6Pt4BSjCLnKXKELhz4jhxHe6v/H80mV22W3RFJM4y6sbTzqub/3W
0wQzNee0T1JNbVe5rHm0LV1jbrjL7hHi6BK49Z7pwgoT3rKq89qg0K1LLKVjNwjhLj8IRUovH/sa
rsPcj/4Y+QTZGRng+qxIOUaZ2cYQ9RbRz2unAjgHgioa4jB/S5HTj4wq/mv5idVEBfDVntWSYX/B
Dcpm2tkHFn9jsfDRCgQJkjbAtNMTxXD49YDknnZAa9PzXwhrEeTsnWbYUOOCydmXEMQluzj+LIZQ
FTKbvPNUNLdWSddau8nJQo3S0kdoiXabulK0zYhHrGXkCHxfQDVgUYZPsvvf3FKjX45l2pvIN8+u
yGc+Ww+7dkEwnsIqq7kCkl/sEpxf98DoKUPq0W4o76pBGxQkTS/InUdhzol5WIYnrHweXUkksu8F
ZHoTiKv/EFHMZt8+bZqDmMlhYeGPnI2nmzr8RL8oGkDdFRDcotLnka0PLmm+K1d8j4XytuR6MT1v
dhkfez7sy9CqVoSEPwk6M7jaQNxNg/gBcPvINCBjLtkZZT0xOtitjTD95h4KZvjaHcRsmYRzvc4i
hjiyQk+FMjtJ7ysg29igtP03etVSlaWj52MLsbfam6+gd45Dc/Fd0DvitScsT2kQChpCCBf7G8lS
5eyAPxupbWlzYcqjw/jDLUdEYrU7c3nkTLtF7aXPW9Bylg5GE0mKoq1BoLWUOHqhidNP9d2LzlQ0
LH/B3QAd/cHDT6ZLTITupGgMPI3PL526v5HJeEMdbqXOKJFy/UQE901He70eJyufk1OvHpUZFhcC
Frkq6Ic0I80fJV61XtLYZPl+dqVm4l7ggoAY4RLk4C9w+0ffkhGtd+2zgOhzK7Q/4BOPBRLDzMm4
DDrq8P+Y3qU8FNFAYPTZU5D56Mk2pIHs9X+JOS20cc+XO1nIbxX0NzIB9ButyhgERb/X+EgjbWp1
8oKBAdC5L3MBLUB3OiNL1Pw0HYyn7bc1DamjUeC5P0fn4qUEg8gkpEQBdkrlXaOLQy2lQyh+x4Ye
H80dnuNM40K9eK7HEwItmDhCbc4JRuiOXt18CQ6GgOqCH4TE8Ka2dtO2KfGFqKHG4T+VxNKiM8Dn
p+5CqwnoAndypYGNoz5WPybjBoC0jBQyjtJBfNdhAo/B2iDpsUBzG0WwP6ZM3+ZpTU3SMtlnib7Z
9635/GNBqTEFHvUrz+amQk1XV0P3NCRcoJcRjsrEU36lHku/+wZj56fIHCbSNqLSxDVnK/rFGtcQ
VG4Xtliwo6x1DLW7W7H86sLAtaORT/N/mHqRXgmtfkiTs+O/QsjsfpKTIZj8zKAMBeEEKzzIeG8U
DQr1qW7onU+MzG8oYwYveADBkqw/I14Bm9BuVSpQ3cJq0J70IkHBmZmQC9m79DG2jFgxcK180LYc
6yxm/4YesFXu2iVQWdm+tf7X+RNg5pGohjx26WXoVHF7VwehUIP7cROd1JqeU/CKFauApazJIPtH
z7ZyEurFBhFeTEY0PgXfS0owOMv+xh1gSqe7GVd0+iQ0qxxrD5/6mL9I2onIm2cbXyk1Os6Xopoi
V8VwwKGOJ3CRUc2VRfonzAn8Ksnijskl70TFyYa1Z5GRwv/4TF0xXR6JXvbnKoxjNJBZGwEGNwTE
hyEvmWHECOXO3HcPgYqwqy5j+2gDYJ7jrCU4zTzYnEFEqVkp91obXJF795+fucvgnw36Tf83YaiU
0n8PwtfQWpxAZolttt8PGm7rK4gfKHKZi/xpd4TjayvJ/UhW8DD6pxw1eo7PAojlh5Jg+1znGx6V
nkOU4AheQAtqzPKvHFURCFKl3Trf4eDX/mx5Sq11xLjbXStscwaQc0PZl3dfM9FuJIjYFL1NJbBt
UyxJrlmdgsX8rsn9PwS3dNQThhQmJtZ/1DKNtiyNkkV4uFNRUED/c3HakSib/fX6Aykc0XDX0qvT
+h4neOn3sJ4a84QamEDBcqdk/gxEXvj618yPt7M9DOOenFKN5rEfy4NNauOC8weZlIA+qB9JraZf
PACVx35d628qhZuDdORJwgOPwkPdxxyefGHkdznYKe949eGCzx+hzT/YBUCRVW31Q4zi5Pe565IR
+ztQcyBuvuRkZjR6+Z7WSPWmD0ckW/CCZGXlTyCPATeIibFi4kchbmb3j0NEqdPbB/JJtrjciJ/q
fSCZ7JRVpY1YpmFjjmBAvreP+Msu1HfwtnnEqKOHuxQoqvjr2K8n944olPvTatE7YEUn9XPp8+bP
+0Ytb4Cl/zD37RvbRMX+hHle85ZWtfHNbhl2ViVHAtYBl0Ow7jrdg7YBJgevPz64Y8vRdY/Mnisf
svkkpmBU4ytj7c39fX5bUJOeR1IWNLrh8hi1Ib5e8kvQcRhKMtX4q4MQpokzuFMb2holZhh9YElz
oDVw1TBkNChywosPzXb1gpLcwbgWH45uBUquLri7bf2nKFXu8BJm/cc4dJUkqUg1gTHFc58uyA57
ul87Crdp6ZJ2vYdYHW42VDDAJZz+mifVUWpsoI8enbe7xybMlwjK27zCdZ+Q8PlsvssVX2kVROu7
SGZeX7eb1iPsXWg14/HG8APOQW3DT28mRaf/LdWb6ylOp+Qro1XUPoXAlPGjUdQq4Q4jKSzLWAeg
zhhkopoqwU8PzblhmJWFsZcr1+j0SKFvQJHGybHAeS58Yizfr8Wlxlj2T4J89HNQBmoFIoNpz5U8
egveTiXGP4sf44qu//EvAm8I/+Co/SM9MIzw7sfIhh4xhyiKLDZm1kdZuYTWvCwkG0Cz7XQxElVv
ZCsc7nkM6OeWOjdp+G7NK0/aBEnfog0YEgIkNJ9YG6kkh5jIzlepH5FKkyxeDPxq1uHir45cpYHd
HCkcmEnUv0HwlrGSlvndGB5rVg8bxT6WocRzlKPONv+eFLO+74VxlYR4I4KjVbeeJLiRDP2o1qLN
CW4AuybiZgmwHXC/GwwDs1KgOxeCaxGvedhQuCq3Mu7bmvuZiyppAcTlLl1ZI48K4vEvhtRMdZjH
djJZ26l417tZZgmDgdck/q7YoZFEVP6VQj+Jry11heP3xnYWL7/KaymydKjvX5/1F//xxtT3/6BZ
7oSM7VyZVeBz3Q/uyG3t16Hzr6EfCDjBAsiRp+ooSGPxRb9k8wi9K3LvogxrgvJVpSFvovm3s/P9
2ZxcXrghzYRPk5muULSedsdgEHTM7cjRlImct02X7dOcOlGogH3G1Px+YxX/NLnHQ034YRA23Wib
JhjSkXDZFFh8cWXG4hn4JbS48wIIeMqvWOMJKQ5xVIu9XgiiDNEoPDLQ8PG/G7+VeuD0/s0LtE+B
dt2R7s9c0z6PdF49dD3AFXdsV0+QhQhQH1HUmIfvzJJfkHuIm0pHB+Zys01yddb7E6FXlvxpzYol
VNGBcsYpuigplOFvW/rUxK7Jq7s0w3jdKAHZDSCfELvBHOnhSyyYFNr4sxvf4PxrbeUS0x+T9i3T
F/Gv5KvPgk+J4r2Bus7CvMjzlJQoisyHRCPyC7smc1Bnfb14yHWtPP+ENVb6BMwEGsABhGNJYgrb
OwefqPYfXiRqgPsS4o6GYSBLQ2gw8QfmzjH9ll1pN3HLsb2yz4kBXgplkdbt+k8XquPIm4Lr7DWC
yN9XPrO9HViza+JLFOV7X84gWn1BW4i0aUBRfJrwyN1qXGRuiSSee4CoDRW8y2ENSSTwBcXbNIOT
XO5PUwFaU3X2y47rCmcPZlseqszyICxFoqstrQpPGtYsDZzKgaxoe2ON/jpx0JR55G/OC1UUpbod
8C3NPfBY8soY2gfNaUb8VYFpcvJdI+H4D7uZoazdYx0J1PEK0il/tFZ8eXUQPePWxdduFKMShPPb
16yC2gPt0eyZPJXFsCEJl6HNpkrOcxuiXyVM2+a/a2TeNG1RsDNBOTc6ccVov7J1vBkEZXvlFWjl
O2LQASAs7drCXkfPMK67fDBI3woUOAGpRbNF1xYwWru5s7uZ8dLBx7tWVoJFBVVIOu+iuHq7btIP
+xD6mxmGpnufHPpANlZcuTLea1EbxuyXWUpPQYysYOtR4nbXlooiyleBcctGc8HE31eLtUM8TgT/
2tzJpEJUxfKeJvoHmcFuRHXnSNEwBSEEj+1OK6v7kA0HBg9WmxZyAU1MEcf19zRBTKIc9Cl5vJmZ
D0WWqQRHJiV/rKje9yzLtmvbCL7KS7ehPawzYxIazj4c94zNXShHd9crJ7QEsFJBybb+8zukfhb/
bOi+ecyTh08zsHfsYSh9mwZ+at6RCc0Jd7rsetQbbImlHZ9cf72cSAVhqo56kf4yVtenIysBfs8e
DA6Im6eXDcoFyoCDke/fY6EbFZOzmwzTx0TAoP24ik2HMUowbfETzkNjA0yig/TOQZPXb9oe5CGj
JQtCannesFL6n5hmN1ECLj4ri0i7FuYy12pT4srfuHZGl2hrw3874Qlv3u03dvU2G2S5oro0cN3A
4FHK0R9WHikacD91h15NeP59ghpea1PnY3itXxCjZg01jft4gcYNG4jSFxH0M9Duyevmp1blEzW2
IuICe2mowtjRk+0hNyGAe6F9Kq9KhBFa1lVBj5O44KxB4X2o+lT+FR3PTn3w5Rwrvs574Eoqpf68
0R2nOSHfVvKYvv0cfjPIlPeaaezviCg0KeoJXWDR+Zr22n2Cb3jvKLHOl4ICD3DY5PJVkCucq/EB
UxGcm3lfEPOQsVnW/qEjYQx0aaTyrsQ9krW+KABZV2VVxxn6NsJM7zJAPxmi5kZg/8ZbVKJyqEdH
qrtJJYzjnhPvSYzAur8APQJ981KLX4e7U9MFPFRaUHvx/SNlqsxzXUJ59j05MYqPr98oLqX7sFTJ
0ejeLhot40URzdgHkj8wVUsgPKZ6g+BSg1JWKy0T1DVN1ejFZkrl87VaPvi9odvQSJG3fQUomLer
aP0FjqleUp+4TDn/IRLfPPYdlwU8cgY+pmRCx+VMV2aqpCkVYnq5tGo8aDBAsAOCtIuO9s8h/7Ya
dX0xSxSofVoCAQsdhN+WQiotwrCYrs1hd4IEjqv+iSHbQQJDSj2mOz1SIbZ+S8immWR3+1a30vEH
n9HioAGYI3pMnLgQIeSZkEvo0TIDKSDf83Z0FDxeEUh+BUnpGtjfnLbYzoIUus5CSriR0xdJYWPm
wUx2rcDC58gyYNJzMHjdCY/cSbro3/3/JeG1se3iPYvkW4UnEuZXj9hrA/146zjxCGXuwyP9NBo4
vjQyxfkDOdIJ/TJqnuFcR2A0wzEgPoJLshRXokvvK2/bbSNWpf0eh01UkOg9ExNj7biSwKIfpgLc
M6u4DAU1sCVDFZqU2DQMrO2Hy3lVR4ezO0ryABK7nGyStNY1G1cZ3nd9Z1lvW6RkiUYLbVtf5MaI
wrL9OGeN/jfm5JavVkMNs/uCWfE5/xYz+EHV63SNUCFNvIZIUR3YHZiyB3q8TfssV84iDzScibVi
ukqgpCi/iByemmIo2KPH9oX7AVQHSZfdaBJlz6v4xkg/iLWeqSpWh+DuIowsHJ39o0MAi8o6okac
NDPhbCBVlwti4adebGPPAIIxIE96azL7TZPyOGMK/EcDYmSFJdNaqeOPHQeBMagZjB/kw4rmiNOk
gdpPbcRuZpYULPGBtRCiVzjYN/M4no2AALxRafZtzcGFxojh+w8okfqcuvQ9d/4+VI43+tx8PQUJ
uU//o289N9FLbNSI/DRj+ik51JBBZr1F9AzcJSUWZw9hGRyn1ybIxIZXedLs6yU801SfW+VXdPYk
j7JD7toLNauLJMGMLEXzxky8OPpWxjm40KVXhcjw7JlfkrxjimlSnzk+9ynOLyaTSfIhmQSIo9/3
4mPV05295PQyOtkMutX5/F4cmiKIyjSyRSdTyTUfFV+wZQOVeqLhTiYT20Sh3NQGSbaXiRflIows
8onizOZsESf3Dy+TrRvB/5LjIogCnPjc3y3RTbzwjpMaO6yk0dnE+AZT48FRUXlDIMdst+eFt5Uq
xam9c148mo4vqJQHI2+z8fs8LwpkWZQhGb1f+GuXl7hyoAm2HTzR5P0W7AunH7C2XDJ8SyekaVmh
wo0EX4ZmAtUEPX69S67KOOLFkvhznv2M1FlY2T3LDamiQdQ9drRyzlLC1UcN81+tD0l7pJ8qOAqw
RiaNokCfXOwemMbtogMKk1ag/djFY1gJ4oKQouNpZjCOxuyoIbj/6JUOZ1GPNuiJAQhWwZ1D6/6v
Z38MtBzATeX/QAvrI6VTv4rI3bW3R+TC/8aApVNuJlxYGG7iNUsp4hhRa63gCoiaxdhDWu1mz+Tg
1Axc5zf+MLvJ5aiYp/OrQ8ZiGPuyUMjHpEuMCVSOQdawR8ZUAg5k54C3Du20sT62SxY4cw5JbzAa
NPwSxie+2StwPFGWQTgot/UDAHppYCjUzBwMGEbhhFKQrq4GBHLVIYEG8ycDn+4Jrn3XopYHwDZ+
+p5Xa1BGTHmUay/4LFg0+go5fYZaYGdvY515E+b7aZs09AZCV+4QcBasEEnzEp1Tg8qGFBpG6v8c
HwKzNs1S5y71N115r+/fAn4iXl3ahUV7VPYfcegSXiHBMJQN+3jFZGvXB9NH/kWM+JAohepi7W/b
HgXsLKYOR2knnS4HtXYUmWRzUWouD54n7CcUm84DRWWbT6BBL78QTf54MxjcKEpuLYofhq6xPR0y
2Oeel66PrBYudu7Ue4RPhwcAwMCBG17Fu4hnUydRqxztW5TmM4+6b5VTvY5JskeTiAnBHgGujIBX
wX6jHgTRA9daihKFAUd8V8B9pF01yE5ES2Hdw2PBEP2LTgBQ8XwFfUltsDhRqh+k2RkawltfjCPh
D4PptxCN1Yb1iEHu9w+IYgsbHng2vhjiFlRUS2ztYhXrIGB6QGUOHn2K9mSxu52SHi9g2tmx7tgp
hINMUcKK30md9kMbrj2jTcKYOP2qmo/u2DxUnaI9rB+DNK12eA/Wlkdt5vj3VguFkOh3CUgjXuNS
KRzNSXvGpEitgXWUKUg5UTbyeF/wUNDkzeFXX7nVVrD0mU+sYLd7S17zaS2bDjS7meWMis9lhJNK
ToOlolmjTLyalMh0yMl/TKKl9m4dwW93p2Gkg41Ac6NQodTwXeCL4/g8Otk27wcQeC/wW0XM0TZ3
I9zSPOSD78MBQx9/rIld+lJQoeh1KXsk9UE/LSDbG/SFBoI4wegAuH+npwaEeXvqFmHBfDxWomh/
a6LJyusX6IhT4/LJ+LpeqoiN82b4FbDWG7SBasFZ45u57iEIgA8acjRr4//tnpf0c4piHmQWGFGy
5q+GD4had//Y0cZp1ql1QO56YmSwHQYX6l31TVA/wy5pJF50jYJ0/uB+toF/z/id45riNaDyICIV
VItAYbH5qeiNLl20yNe3JW9gu1uUK1ScCacMLsKp34ynkJe+xyciq5NfeBrwUF+5gfUkgFD7V9Qj
4v3Z5TjtLz3bHBVDUCrMLu0yKXlqUNTr9HA1chzfD0/k8CBQzHpVYRuvOFHwY0vXBqA9UNTJEXyO
S1g1UMyGI3+Fl8auT1rKtetBlYjr1q6JHuAGZ/jgJ0vSFt0Qq5ejx+3BttGwU9ubpDdGonMrfrY9
bCJ09tbZ00vcAGKUMN+m/tIidgCtrgj+qMcPBE6R1lwhbvjktlB8zqqjqLsq2nVBtpvV6Ye5fgNY
flFQdaPbgFOyPRgyduwvzl/UtOdLg8Wyukz3FbG0xaDK4CtxLHnj6ZX22/yRSO+sxXPsww6j8X79
KWHVYjpdvM2H6jCyPM0JSNpU4FWygO3/KSSVE2icYM+iA/GP6msyKUshso2Sj+q5eshoqo2GVIl3
r412s4cFSlceDQKnkZCB+xxNfPtDRiK4onCJWQlBmscPLq0yojxy7pKXvFiRZ9I7evngy2Xq1Mj7
n+tUBcUtrfF8NCpDeCOeWqHJXQy1iRuUusljxLlJ2VOGAF85eKg8sCDPj/ETijsE6jwq++i6IJmh
5bP11F0GUlcoks1R2Bm2bCPd+0kfIkc1ilnHlfSnI6KitgCKCH029ZkQo4+V5BI9zV9LFARjeBLA
qFn2l0jvErVXxGNBA1wK6qa5XOhNwe8TwySh6+Pqgw4OnaNP65Yg6KwXeMotQyHxcC9p0WlGZ+qp
CIKt+5dRkvixdgpWRovr7CxX/hsEnOXU/Nl0NyzeGcKPorlCyszOSKsA3gD+nurE9LCdwptOn7Wj
i/EoDivPa6b2U3BGp8J/qb2zYoRFVPH2n5V1j3KCgZTMPArnBHCWZXPPiwGlBGSeXbgKWgOUiLwY
CSRrRdkiCpDkAVQaTYqnvOZ7PxfaaDCqzN0IFwU+daKozWSXPcllO+ZVYkWTcGgjFIRjuDIL44AK
sXXDjEA3uVFDGEurrsExdGpAWUlcZOOITooDuOvtFhnGs5KCu/JS/yWwY1XHQAOxMH/lEc5vYCPW
7neVsFTGt2VRzZZh+TH49tAI9GaBdYkJxHb0Tn3A+m121/ebb8szhaT0EPNfqrajUNbBDdS9G8ve
3aLUdgfCvINoo/HM2RPQl6b9StcloRYHlUUAK+t7QCXbemU/yDRMc0mrbfhnSTFfRFn8wpsXP12R
Lv74jdghJA7ROl1KupDy8JzY7HpBaw6ZpNznQkVhmZTYzCmMzwxFnYsDFGp7rxb6HyvsNgzL1PuY
ZrMH9JnQIVkL4udFRShPQnljDeKkH62fM6ugViKh1nsqm6ZMs+XLRqPu8ahr8vL77VHWWwHu6wwi
vHKLF0sS1tSQ6AZkb+jGQCkhNpyAosK5lPXFrhPp9dA3l+fOht84vc8aQKqwA9S0jThF8CEuZR1L
1JsHT5GiQjqPDBWtCfNBiQKVVAYiuFjM480qy/6D1Vcj7JoSQcAz6cktDJHSH4gguabWz1oQ9Gd2
aOvod7iqBugk6G1D6OMKLTyBxa4rR0+ZhTCjCr6XaQxFPpy8K6SG90mRByezTylaRExiHO4eq5re
x2J4qkSAOju8xlLSXa4JoDYvIIrf0Fb62m4iEV84XnoNcCBFpPQi1ZOPLKEB6NQrYCnJ22hjOdGY
9pFVhtMm3iz7TwxlOxuOTIy/uRDjyBteeqnjLFM3fMM2OOOPb40rm0k8XJ6hxkSvMkjZmuEv95fU
EkLn5vQwqTXOMiLmyg64ftynH+SHyB5SlUsbM+tdf1E4eTbJRt6JHM6rihIK7suVe9TdapNLjeFB
QDV6FJxEmrslLGsrP2/aeSuWSpL2KHWMY8YWk0bAGC+LgW8lEuj7EntSXwu0dYoFkiqMyzJs1jL4
lEjhuJvEVxYXnSeS/1Wp5L6DWbO1LLDkpSAoD0YJlpRF/8qJVoASXj4aBq4Uu8QsxTMJnwpzC2Wb
XgNsVfHn3xW0huXSRRq2NwEz+C/T2/OMcx20/ZuqroKxzazgWoMw4vsp9G5DWBVo/dyfDsE/O1g6
0k51LjsQqaPVw75R7lmW2kCzzzvPLdJYN9KyN1rgf5mG7l4oPEh4b/eUNCVVbK4FvWlmGFoTxL/q
84aO8MoFsGEOieRdGf1wMdTI3zY+SLf6c5NGqEUYhMCZJ8rdnMuYtVHarcT2UAVWwOfnEjdPuz4G
3I18vhOpTJ+Yp6bju3h8YwKbvCXStwGatbt6Jqb1Jgb8/xXPebVvOGD+JqlfjTHbAoG6QO55iB7g
AKObm7brX6zg3hAY8Gb96QPDLpm6aodI9DrJ2Sg8WTRlSNtm8yWWvP3hsn4X+SO+UCgIc/zxqV92
cfLWVf0J5cgeQ06U+ZA82qEBBT9U3m8TodI0iw7YV72NR74nTtd0B7aPhO4G7Px3RJSUYcXMPk4Q
tt4GsKya6n3dii5c48tDQ8oR9nwZYmeg6q1+qPqOH2GY+6EBr1q1V92GRo3FM5xfadhx9SiLvuTz
sFYBL0TdZ2o9HRqfPXgAWy8KLt0DVA8mX3aF0PfgToQqAsVVYwh+FF2UX3Y9dTYXtTei8mNA6m4s
pe5gdjVtz0QBVwK63bmQvYv9XOL8JtCjRC5z3onhxZsEt40PatxRaD+ltIU/E+vmMWQ8AuDfcfPo
rXGP4BFcIfG0e8LuaRJbKGzCX7SOcxXJAspGHjNFnXZEjuZcaPACPh+eFD3Amrm5wgZ/TPgLsRR8
+rX2LnTiYl/mGLTYWD07pREiJgd8JyNOywPFSN8LEFwQOvfUmZ5bIovQGAIgoOqRr4hUm4CZoa8F
CHIJwRGll80452w4A+C5TogqpDOAguAUD3lxdfe+2HMJMEIHr0uDfH3zGWdUPMkd8ytnh30r44+z
64VMafk2gc9tAB5SILkN6BfNu8rLpFQ5hRDl/kioBDc8IDpxxdjAv3C2csa0JM1oOhjqLj1ABeor
od5KAOXcBpLsEpHGBmzUYIMU92Z/7c9QnDx+U1ZTZy0UjEYz2XbncA1g+vt5Ulk+Sv+Q41vYCBIu
Ezjlx382167hOEqtu3M07lMq0Xyzs4L6Hh1SpBRODVLXtqar53wPjG7wU0xOLMPXbG4QKYeBj7xz
IsfCLivOnHq/GEV6+7apwOBGaH5ULl3K3YP/fgI+puWEV/q6drbT4KGkEmwibluJcRg04w2Wlhae
FpI9MAs+Y4HssICGmZh4esi32wuc2LatwN5Ixl130BgJBpS5uObtZSPQiQvw4LINJrV03ORKuUa6
S8WcWh4C4LvKC5PJLm8ToCeXP9LlobuaUhoUonP24PUoz+gREsKPbgSu3PwYULMP8swEwNR/faqv
0+YkINnSrazcEhQ7xKZfW8+CUpe8keNXtMcpwQYNOLlovZUmwCDEPX078fvMRFtqhy5bRy8mxC4M
Xmjzf89gzuOmanS7xE86AilYJhtRNDDBeidmFITUMLOoZon9C1nE6BeQbM4uQFiW7wyp4T2t1yin
xbTXwGFR1K5nD0SugTBVNuRQgsySGswiyQfmoRc8D2FMLqaK100Ik9dzpviuqCTKdAgMktIzS0nX
kYRHcaxd6dTPatOIPrQyzg2kviM3jJ5J+QMYPgLQkISDlY1EwmFrRU0NdO0z+Hog4P97G85nr+IX
IyspeKVk7tg6XCNYP/TSUANF01PQHO52wtxUOkc994sAZu8U2glWoK/HkZk0m9VLLakCPCsZ94Tx
6M1IFGvSwMHH4cF43jHHa1E306nYZy/Wo0HNXdHPcYZeCKG+AyGXHJ6D9wQN+jTJAJ2f+1c7+0AG
NNlmQHTN5nYjucnQMaQ/Ded/zsmpMYfoy7ytLG9yUzRsG4AwdcU0cjNQgywkMXVEzbHodrAgo+sz
8AwIN3odhBOpJH2lbG0PeqeyyrgSShrN3qd4Lk55jGDnghrbX9Kz8BdYn1nTzb99mhzMOUJcMrIk
bYw/m74A9pxyWIfz5RFNhcDt7uqjeaf3/p70LF0i7yYVhT7Cd3z4fVCQjl6C2J8dYCxYe0mDsEz5
HABVIxf9dH9dtLWo3KY+9HF8kZVU8E82jeZRAL5MXIUCKNmqrp+nKQKY/K3jrJXpYMou77cZyKgT
qnsmKHKsscH40P90MAKNoLPW0akdSJuglVrNSgOlPEj+/2Pw48ZSYJBWlTdFZkUbz4s5u0YwgNQX
rkiuFIMXVowTed+xItKSywUsyXtUFamnAAqqATyLOVm0JPyVv15py9+T4qeklMky4Bxs0auFiniX
eWWTbLJdKWB14YPRy1RKfiWAtDOwZ+ayObkkS+wKb4hUjs3A2eWbDiJEq7914PFaiXsAGKLGU9IF
1F6oclqRelrp7cMKz9+V3DNy4NHfIKDuhQ/RC9i032jFq+PZZm4x7u78rix686TonKj7sU8ZrDj7
IKwJIjLPFwB3PafMYjZb56aixz8twxg8NygrppoSGsmy43rtyfEGL1QWq74ZbnDPIaPEk7Mx8xfB
t2FVnSrX0q5wFcf3Lt5ds0aPVVnkAWEK3FrrudIOmA2Kr7J+z2MipVjDPXhLCM2KHDjsVpfc+T1T
F9gtoeuSb3/Tmop/2CHN6/FXencKw0WPMNp3kuF+iMqX7MwJ5JNfTWsKnlCZDAYDVp3+RXcCL5sL
jRXz4k0ytCgYh/Kg610BIBYY/iqiUTWwTVj48EBvLcdWl4HPlxykVyR9ekrxwzASO8fsrvcUWFEJ
2BrSBXxwSsBXGzKbkqr2MaOqiGeg1WhvsU32nKompVdxjq4ome+BIJ/tBHba3CffmERKLdByxWas
MxgIq3qXhHKbNvpvKiUriNLqwifAe2xzcz9OJL6d6KeXN+n6dxsCrPREjjdpA1g/2iAIyHZlbkhT
B42CQDhve18G3QL5o8sXSaw1KzMbTmKxpEiygZZy5ISrRQZIDCCMz7Vpf2wLNBohnj/3o30b6JtS
z+CKK8gHCB6lGRnpzt07OBif/Eu9jl7eiWDqZ7YbdZSW1AOKe0wOqIfHJI34qIFpg0uOjxf/82GW
x4XCEoSXhq2PDObDcxovRXpTUmXsAPAvqP5gvSPlhBg9UvhA1mvHf4SDzadqEoLV0WxCLXu1vZqT
/0wvExPByZ83RYlZPrgWcraQWHTS1QkHwRH/D8LakoF9TPjFeSCn+4c1QKoSlU98OinhysfIL7Wr
CqFib6p+cIrfhVAxLc5Nibb94/hyJkFiL0+Iq7gpq152VtXIoEzgNjrbozPbnA+AeJrDeOJIHQhc
WmwbzOBtctqu7aDIz69sC+QvtlaxPKm/8rMnlS3cKmNP1TeYZTVb9lomdv+2kTksXEzO/OPn20so
ttoSZl9HK3BmimizXF7M/PUtZ8I9cV32nPfhTCpi7QSjOzyJKzpiGbfm+xReTgrs9w/832M4VA9m
fcWZv/ItjxYMufQGDU/xy2qQ3yi8TWXYyclaKXL9DG/Ktn67JUq6uiFMIuUe0DiaOXZJBnlq9dqh
UoMOBHxpwZLjrp7/lKmSA0U4LbUzM0hHNJeFrRENrUaW0v7rIBjnZxSMBq04S3sRSepmnCtFfq3s
kW8Kp9rYx3gTeVsu0zE0L/D08fI0Ppj6q4SocY+bbYnduMB2jvkGAiWwDDHjiyrGuLSiC6I0djxm
VeJA6S1mzaRxW4IO7R/tnYBKAWwAzhSGH4FSUt5HKfJPAGbCcKd3vKKAYcQxrQU+owP+K+a/YPa7
1eCMH2tJ+cvT/3bZ8JcNmjp4iA1SeYLWUR3n75zyVs274DN4f9nOmq4mCUR8nQX9klkTdeVjs7Bm
0YZXHuG7iNDKHph4PPe2WUZ61jJWAthsnwbp8SsCwpTmgKcmaSqEATCj9JGNM43cs9vt3JmG4CrJ
ejhuyM1AWAwLzLsFScBltY+eFZhrxfNSGRpH+TmHLyswxo8DImW+Uyu/LbYv+cSv1xy98iO3dP0D
VgpKtj8Akdm0O4yTvYIf3C+cZTcYrKvmYK2ywsECnyPCVs6hTJZDseThhTwawV072nMFQQ7BFNWq
zqE5IAovwtdOLoir2D5rJgtIpn8RqHFa6BoRYSvrChnXUVGpnJiCwnfHO2Lft4UBC4ijNW6xKh/c
lB1cspesF3I2RuLnjk0VTNX1e1eVYTb4NRN71ZLMQm3OcDOVebmfNQ4gZBwH5EvPAY7KzE/FjVJv
syjHWA1dp2oO6pFUOmEw3+SnxY+Fn/ET5363xwR8r3YhcytSSAkenk1bF6fW2hnEFnnog6Sn1Pyh
giv5VSyP0vxdFkDEKFODRBfuPqGIcSm9oGS6yyUWYAhVK0031q/vyOzfyB/IlLqr3U2lUWTGmgKS
cp1YhjYo7AI8BoimVp4yO09QqXbuttiVbbAaAuti8Ao9sw4UVJULerl+FbbqXnFnZk4XG9AwbN1k
eEoxA6jW4O9+XoX3XpcB8U+fc7eORmlRGMYZH/2n54oDUfFIz7P/bM+3iLU0h8XoZJbb2HZFBbr9
dFP+Wfk43l3zQyFREItsDiOt6u4OYE7ad4K+/xJv1qqAKMPLQalwsyUjZic8gaaEY7IlLnAuOnWU
5i+rCJofjNJVimaFA9rQMjQqa8CVVhiWBBScANU9Q8hK16DP1At0NCbrdQvZXmU6OJxdjhEc1HpR
0yel+ovp2q/Lwqrc67yqkDoMfm+Yl3ap3oM9C//pTkJ9BGK2o/2sERjhA7IQZjZS6tQIJcdKZdQM
dGI3z8rOKUX+ueMXroOEJKv2m7teyY4OI2DqAi3uLEmZ9mfTz8rEY8kbmFu4z7ap4QM77FPDee5q
R8g/VFF/BKnO5ZWmMUAFvr5MUJQ0gSBCwdMyDduX0e8PuTYRK3e/ECztLwm6smpHdAV/v94mevKy
8SJYRkHOG4jngGn42Tm8/SSKAhIzbvVkth/3f4GkJQr9BF3GRHPIAYLeBCLiHsjpfH2CZ8ALdV3N
NS8rlvNHSTt31JZnsrMWIIvc/EvsfXtvLnx6OB1IZIQjgZulliP0CY+DR30tWZ95+drYLuXr4Vvd
3Hl9VxIXXouXnUOL+02FfgZyXMFcHLLVOtEZQxWwCFFrjUi1g/OUaPiX1z08o4v/AyXUtHP6mSlZ
O1rTIPqDO5IaHhDzYpPJqac8X4v5P9HTYD6txnE3Do6vQeeB8QqhaG7VorkAU8ZzsX0kZHoCEMDd
+vkpvKq8Qg11AIhWjwAn9QRAcO/RPOomD1tmM4HtcGMSxND2eJ7BfXwuRNfxD5K4sTcJ6YfWrhQA
bDiUl3jUMGEEenohx4w0Z5nHLjTbJSh3upRIFfdPR0x7w1jWoCDhMVKIPFE41SRW2x54O5fBUqXr
SOpHb8+P8DDgJd17vz0ZKbDj+QtCxqbVeEdP0qGlEpazQywe9ParXkohWzZLlk1eeT+yhxvDKJYX
whdy2G68rO1gn/hDECnbAhkUQZInYIF1MIxOOjjiMUvqs+NepKxWsoe2uiqbCOZsMl4PBNR4IHao
2/I2Bekd8rK2DNrFLNd8jgCJSEDsE18kthSUwN0GK8xJTHSwJGTil1iHNUnqqYzydpKjyH2+clha
EisnQc3cBIMOwJ4pgv60PHUJBMoYgPincYvi99BQ92D02Stseznne5DYcXsKtRenudF+e3EBlRYD
M5T5rdIDkt38Putwc49hSZzW3h8eGitLlcuqiRNxWW6tXVT/S+s8XeaQ+xkzseuXV0aA4izfmMm9
9zCeq1kxkybMqvWtPfRO1GoonkIG2aChaCHinK6Z/Rt9H7oHvN/etqtDCZqt1wmqfZlL+evRXIHb
t6v4IRof8UTJsB8Ok9W9tLyrViCEIxhsAT323njYtaPGT9SDBtarxKDI0CedXQdHWxaoc6h2Y/gC
Lgb8LauyI24I+iFF+UtojSSF+T52uBVEK+kJvYhDJKf8SC0iqseTExGXLPLSPOU0fMOwhOC+mOqU
gXvYKH2SfDUA5YzDtWHk03XUyaYpGfocDECEOOWP412kowQqvHGcVXH1Oh547q+/xC+SMLeEQ4Vk
BzcErgIyUf+AA4tSBHSa4RJH9lemOxOv/WmkJn/Mke6y/T3Vq1M2C9lQYva7HToNxLx2G/fJZJDS
KE8iOoDSuuUiC8FXdwWVSqgZDDflXLR3JnJO32SHnVzNMJz4l9K9Ka7GLvhd+oMxvw/r3MWnMeCP
XEcJiS+GuPR2aNg9Lao1GFtvpoO6swttGeYJzHUirqMZ7OP424obppEeI3q2VIYDOyIf3Z8V938D
UjkFSDWc3Hw5nZ2OVMAKs9F8xMd+1y5po6x7VuPTMv5TpKWm+FSZwK7J8S1UrCAnM1EK1QU9c5dV
1tg+AeTcIGpkqz+gOBV/nOS65W4sdDuHewN+dMiclKEne+S2aNI3t5A7YcGDi+IzuEGo2QjCmXGy
WYQjHgfw80yaEvAnuW8qepEBLKKbG4p4u9Pxyp1jRNltbIgLbAxwahYoDcz9jN1sTtJ2rRZj0S5x
Cm+oW3PZtIlLV639Ggp6fV6e4xTMg2OXFg15d6sT5u9LTjWxqdH7+CdKzo6XpiWDhNgxKVZJt+L7
uL/PiRYcPZBznGDvoqx6o8hmFjG/OWtXjuzPQpM10KHexq1l0Ivb1gho/PjE5f7h3beMj2zNjQ9u
ALXrQuhjXHAUxA87FUYGf5owpcq7jseb8cN2phD8nWySc21MgTbUe2dxmfpl+XiYxtxpHO8ZA450
SKR+Jr45INADSpY+z2ncWmUXVeijAzny1kHQYpR+wCLUWiAUxKyzR44sNHlcaz4bMwhNmAGNnpas
IAkFqJxwNxXElD4yGMjHkMtTZXh97jT5yYsK3rnw7Lo833z5Bxuy0ZOIlKISxxng6yADNplEVlIg
1r0yKK4+eL20l2CT1uvZRYp6qym9eJ8VracyNDlI2jORmT7sSFDd/7ulbVbw2h5W4NGpAtyiPpUG
VXFUog2w7UtM3hvuzPG6I6FxEXr10tCFsh4TNxmtVUg6mh5/O0XV+cqXqTM+PqEIBCIdiJHWg/dA
VND4A6H5l8we4aueJ/Zbm8mPi/la2sYZoC0k8kxxIGDLrIMyXSfMQNm4EAO/dpQuhl4iQKG3ShUg
3C+yry4lhy9xsHYuz63dJ/zbHfEpcn7FeLuBDy8vDGAAg/xGAtaLNrWp+0WZLfE3ii/HyNlKSl3w
XvCcs9ZfVc6P2WsYw6rgZoO1vHqnYLkGp1T/d/qbd3G90iAtElxqGN52ZNqWw3ONTsvoZYSZMKTF
/sgIPEAZSpxIrr2QvVbvadXTuz9qiB8rtvsHNIrVnfX3o9/ef6m9u/j6dXGCLl+1t1qPz3gGnFow
6e1XXhoKNPu0p58wVqBpe5zavzfViaLYMLypjCFjjsA9IBJjWu/cr1Ys093h44hWPrfbxgdyI6+1
MAooplULkUFuKmNR48dPGQWifCCAh9TIRFVQHDcAc1JKTD366de8Q7UscjRRSonizf7fjPcToxDz
xEoMB6YofFkaiQupVpDH1x9aKh6PcFDOf7KCXYDS04HIJBppyZdS1sjeVeTTL62VXnbCFQBHg1G2
/+Z5X1TwGTHUZwyggWb+OSzPgL6CDDID1t7dLKQ8dqDc6dt+UxhRcGQRZQJgdSA9xTd2gYVQykeN
RamJ03V3WWpq2k/RcAPOnPfVZtA7exVDWRA7QoR4+uQMhufGRuC5tgw8Guy0uKR8ynllL6xBfvSD
/cTyND+VGCFX2cOhK6Xb5tbzbdubE/YjA5nMCjBDwh98713IG85S0tIyiwS2k2IbUSzxscecLlFK
oGd8mlAOkTjdaX0DqCAgHvNMC+beiQLSufpMPamlRen50SWf9LWDFjpHflmQcLtZAzH9F0GDFeFw
4WH2syiGavrpEFV+zaHJcKxxU9260iNSzFQOMcaTOAHAMWwRovve6LdsfsvqBFPwm0J+IwcHMkBG
lke2hDXMvwUtQWWY041AUh/sLfYhFISle28RESkZf5UDQxlyEBCeEL3xa5jF0m+xVK4hB/ehGEDM
zDg6fUZ2n9+eo7JhV3Ja0Ey63AyTnYBJoy6KanVU9vRn6EKVKCUambiKuKplyctqFKiL3ICrv4QQ
/n6IlqGiYdxoQ3usiPxYc4OycCTGhclX7krhk0XxopO/HUUS79zEriQClAzL98RDEHkmWh2kAGyE
zahHKGlB4lUnsrmOYk30iYsK85zV2fO1vnMaVjnHf92vEt5yr6Ky7tK5eNqgx7uG8DMq03CXaU9e
VU2GXcsmYQswkl7vHWyvG0Jnu3Ag2CeQ+B3WOmh1crBWvmwgS+B2tbzTBGKmcJqM/vAChQnV/CIU
gLFDU6d9jcSO6v59UOCCwQkFvhshrHh5JSM36gfa+rDj4dFV3zGV/B1mlBfltWUshh2q7DPR7JDG
FcVKoXuz84QlY3ZoaRZGnkGJRoYnzSJQ5wlCQm185jVU0PJlVzOxx1ynxBiQwklRWpN7xnWkHQX7
wwSs77IIBIWT7QUY9g3OWGPim6OO7Afa/5rJFPslIt6mnbQmT4zgz4NM+4X4yPiVSh/UznzCjcsT
YUZoa/itR2w+aztw7Xdl1tB0BzCGwOA+IzuXgYTLlet1XX2+gWOHJXWWQ+AtSjh1qG9r+uMAeXl0
+Fx/Y8+U/6gNXUbsjq9W9j5ar1/u6MK//zhEcstiCF/iBufSnrv46nysoyoNLfiumwDXsh+QzIR9
FNK14p0Xr3CtZmVmRQgDwmQqvnAPbDdPZ6p5pFc0W0j9P1Oli3GgfmcTNkE91XK0QO5XM12xHBVN
gNvnykwcjtXeGV1Amk2mmRBbGnDgLwdaDh7m5WjiIYo8pfBPhkwW7kZ7oRVlYs284fsnv1DZhb3Z
uVy7CgHEYm0AApsMDDSaAkTHCUWDeYdjOxiXlOFW0uvAlw6dR3kL5gwVXvnrDJ5iVeZEAZDtOT2p
7HTBaP9IgtBS4sD8EJOfklot5pHRU1Ew/t0l4QFCUivRrBUMp4oHwxFjBP17G9TlB0zWj8Tmv9hX
MjXQID62DCao3cfaLMv/qwbFutHstfmI3ipQ5QmF5ydo+Cq28jOf7abIdXI6jcOrq5grpdH0CSvN
55ebUKlpK2bTSXVWUWRH7UMvQcblhZ0JXszdaf2y8+q0WYKBPGYjgHag5/IIGYSXnhFzuT2q3d13
eZ2qovPQpiWSFZ4qL6LZVkBlG49YJjA9dKZfzneooDysnt3bVEXF1w8K5vlcyRltJ5SD5R1jyCGc
hZ+GLRxOdnwRRG2nrmz+36pWQcz9vlD9NVVNxs3cZYuA1fJ6cjSo53Ec+hoHYS55y2Q0l8ex76+b
A+GbZspK8iDI1T0E1Ma3sb78w6OplE4820x5KslxHPFHXUnIaR/+rms1VZuxQM5BTiNEL2+XVgEM
7Sq5vmZtFSNy1AfYn6IYlWT1EA40DAPppWhPrMx667Vgmf2ome2T5zj+WQFF3KFGO/pRbjOMO/mn
IPgqb1LxcD4pk2UhbrBGOeCMvhY+yIiihd9JjSKni2u9H1wSrNa+JBhwOgYscZ7rRhYZizasBSdA
dquq1YCnzuwCKvpukXs4aq5yBmxZXHrJvJ9dF1CBSJ1XTJ2ItJwPCjWRxl3LzEV5khQT03AWRIbV
9GLRJixN2wFa3WNOOTsK1q2oxlNMhTiIQ/tYBAI8LkDIfbhPDLaD6RngCFRfFj9t0S9tEpHc6Mlh
IZIJYYrgFl6Hb+MBvsKT6ixb1lxQ/aasiRVeCB0ig5wKWUAHNDodWsQeLF9lGzoj2x5EquMpLZIR
WuXhxy79fqY/jyqIrNFgMIDetbVLOC12E6o5lFgiVGw0rZbNPiTTOumHKUVZ2JOmIkfN+E5873vm
+YRCrcWCYOgtJUyfEnnx1SHKswWNCK4tN/7I768PDK5amUqFUkJLPq5ja1VFzmeoVi7dmRwPpKSo
DCipiaVLs1I2E3aJb7xpqHnjy2QChL+K+CqDxiO8G/qFcahjPShUAWIrH8gtfH4m96a1euYtpd0f
64w4NclHgQXw1JIgYdoFFYOHDn7Dn1BxxiVDGYmPU3KYJjdnzE3RDD0/HbJBHPjCna5EyKjj7aZA
ec6t/2Cc8pN/IX5os2/LeMWmIxcuVQZ2f+kpXzdB+yxcEiAYGpc3szKUKMyw4ArINGb8egUist+P
WC5IBSz0wSsNpn3MAw30yhgpKOu9xFIlmjT/IOCfBD3ilODJTYd07kPvH3jpBlFO4j5hhQ30+K8T
4BevR/BQfDE9cdW9bKS2hejp4OFxSvqWUCwiQfLz8OvMf09atzLdxbaGpn1SvnZEJvy9ip6doQGt
B/buN4X5XE3GzHJTrB/NcU05JcRPao/9XSdVG6A+LAnWB6uNFV30EW9NLAJ3EHbfOehThqWWmAPV
GXKVSRe5CnGomnkM3mdPxH2bcLnGbcQ2Z1wJKWEekD30I4HlJmebfYCXljXkZTMK6WXvIFNXZptH
iSolO7DWKM1/g0MunxhYuk1DxYhAxn8RdWEaj7mSgUAr+cbERkHySFU95D0kuVZznRPGW1Tn5+Yb
jrDaOjBqiC/N8PzyWzszOHMLsZUvsE8QR8hPD2eNxrCWA0ai9PHg1zULG8bmE2yXZLeqYQOcrWg6
6YMuB53TmDgwiVxH4K7sXdX324XL1tb01UqnVgbyVaKZ1TtM2h4Wh00Hqwvv7Ok51zw0OIEJZEFV
+rrsfes0cSDwWOEaTCHnJfWvVxS4yGkmiU6dLfSSZSkfXWB8Wmcy7lrK3xlgw+pPW7WVWWdgDiWO
jRFh7j60tZ2MVw3ZGQCwGC0Yu6ZklCoEMFwDQ2NkfRsfEEG8IJ2DY+JBEru4ahrCVDWzsItaf5bz
dszAnGpRbydUp2fJRlX5d7q1NbLOGt53xBS7hXndohB/qmgy83NqUSG1W+vRLNKIaW/8G1ZZ2i5X
rLtfCACHyW/FA2+uypDjhLiKKoOAM3RBbXmn1kblrzHybqFq11DfMyQ7CbM4Cpggr4vEAVUjddMK
96s11makRWGQMy0FZ4jx6EnobWDA9idJRXo9brVMq1yi9ypE3+ErtWrzL8kRob7qySbiq2x9FPIK
AVUsXydljUpC2lTiG84z2JWdiPNjS4aEci228hFOUXcrkTU+qZg1BDkZ20BpAqjs6sy98jgEpvQr
eaAouo3ei17JLwm+g8WI1H5XayxUizwkFGPxbxUQu6aQ2vM8iSoIWlnBqbsXOg3g+klv3hljMahr
LfNbzFOArcuJU57RFAyXa4fCPeB0g2Q+IuYBoiiFtS+k8w2R9qpw+j1d36sREuNojHxifSTaxUrM
WpmyfttxSkU0hcWPsWHQwdwqd/ej+MVVUq2SsXvFt/WVZMpj9o2b5sXrTOhirxNz6Fi3S4qkkaAy
vGXno7n+9m7+ONkvziiwNOxDMryRvzWb1YA0EO/0De9YSjIuBi3kLJNjcJsb79T5/Qm0YafXUUdI
6G35SMvzPwyX6I7hnWBMdLpfwsJ9VTY2QebTgXDYRzRfW2S3q8fcHxz6g5MtjfyezAsN+fH+much
RENomvgwFL2suhyfRfIb27PSYN3EGIO1G0W1HKgevrdWD3qYBCbw0yEXHwyf0c479XCYQ3Ov5Sy1
k77LSYlbpor4W7RWhEGdO4ThycFL5TqaPSHjMQyf0gzg36dj1dox00PjfoLyrPw3UX0BAXwMU7pR
uJOf9Ksh1mNTIlsi6aq9+ywgOjYUQ8j5sNmRfHOPqp752zjCYmVRzvgxDSpAMRuS23mzhgbf5DZ/
UlgqedTaraQZHcI6u0Xwz+Rq44ytIOZaXFaMKVmjpOPE42UJLLfgmM44JAiRmXKtRIKrbtMfuOj7
+B7mUzIdKCU4EfMg8i9RVhK3Et91m5ZjwtVO1Z1GiQ4LulLFukUMarCmM6W4LjAyyCGUerz3sU0T
1rMnwPM2nc1WhRdF+yhg6j8QYPoT4aOAtdmzXNQY1xuHFbhM9y6XP7zrbk0JighJ2VMB23WA9uUP
lFqmQDZ+7k4VPCER1Upo1aSbVc0NZnnokrOteI+HpSXRf2QcAaqIJJZ6lbye17XyzzYI6UC8dsf9
cIFacF1unOHWy3Kv8SPS3b07Pzfz7sOk0H38kwo6i0IFaiIsy/WV52e2Yy8FHdQ2Q6igu6oZXgaA
QunKwMKI4p6oC3lezaD/DY4fnufFID6AA/0cxe/2PdX393fFDoyV0jWmzePzfe2LyRZZgaDPwi5H
RU2BJzLq63MH61AM8CHmiZAXlIeYIIBPJzJyBH8pNJKatifasufgo6pIVloMOmcE31gANndvfKLk
+P2KJYcUQleTpQ80pHaMMYMTm4ZdA0FsxZ65we2WtrrLjFK5gTkrzxifZ+4+yHsi9PdzqhdADvlE
/nxEWhjgsSqJxL/nzZoyNGD3phoDK9vHf+g5ShFFaVZYVY9eDI+EgTbamHa0I3/AB8gHH17ygFo9
rv2yZ/JXYBbBKVgCE/nfy2Iu8VR7hHQsV+piEDQuOigEHRY4yJ8aFWyVXrDm2cXdetyYyLhF2UiW
NLzxlEqSaijsWARUEqH6yt89dQ6IRzq2LIWH6YjuWk6yNSVoZ5e3dZrExV616047JBieL9lluTOv
Rs0pLVjs1dkCkzyQuA8C7uGb0UO/lmsBWJNKdLImN31rtR3kWzHQNuaWje3m8LwvHc/Nsvq76ABo
W4FBRQYoQING6Xh3dYbsr1zdtlwr55pzpW6UlNm3i4WbRm7GmxKT8dCiEizxcV+HxrICdG5Yn/12
OBoWplX6DKQKWd7+5sngs3E6a7F10uN5ckAamptoo8FFK9Ya5ghCtJoHv6kozI2GDCYkbzKU9rkR
DOl0oLYarjSNbfiLCmVEK9R9zumcRGfsGDLrgIPzFL5+8MV0L2YLDkRsf46p7CPn+5Te8Z9JAv4l
Hf5ogCtKwSAse5rfVUzvvII8ZEnjaG+ZgDgJFWl2IhHZIbkLyaRQ/CdSBA6k0FGjqJxbgk/7d+Dw
/yQJf26MOjU/ij4wYhMLx6S5wyEbpv0uwY8KIgCgtRFxuyQK8vvFd91Ih841NQZxkqZHxjkraOmS
D8P/lTipFe0kAzz6icc4BP1JHAujXF5b8uZDikUP7qkHXr7pFRlZl0w8TTKtiJjd2j3fdK1BIheT
wFu6qqOtfWpYQ4rFhH1iIbLCdd9bvdKxdM4+vH+zb1a82nukimTGlaOVoyn0OvvZj/pZ/NnBAoNd
hIbvIzWuFF7nPSnT1SyDHKK656EoOXDAbKOapzc+vWzYs6tkbsCxH1qjIuyeydKxYniRQGXMF0xs
PEOQavrDVv0zTyCvPvKfD3cfku0LL705TIZs4eYDCvE3nwd+AQ659xc4q679trOlUZVYp5GVbYMQ
e8o7d6qZOiJD8iUNA+qwWX9egFm+btKZrchY5RZaH+qNakv4KWAd9zXiqxTtDQetEp80mCYuGX1l
Z7zxnRZ6M3tbSlJze0AddLvZ+Xr7Y8F6lhH2pqFvCiBeKB3rzcok++73Ww+qcsweyUhkpKHMeAI9
imPD+0kkfDiv0/wkSfLvVNw3K0HSh2y0yVmewjTcWDkmF5WxicFs7EwfkLYVGY0yMftDmZG8AOO0
QhenPmi1WfF+pDf8JIoHQukQjPayJjW1xgZ/VjkvvoYhvf4aqzsjTPWoqg9d5dsPOOxXaDRHObUl
Z1Bc9FZld7iNssD8r7gtY1caA77Ds8u8Qr6DyQpLmBoriZaMjTWhGAaFUndpEEYPCXVfxGwnH9jl
0d9gKPp3Fpn+dwcvFhvBcXXuMAMOCFFvryWHH4uuSWvsowWb6fZIhUQIoOeFDoTFrvcx6mIGu864
UYgzZllAF+IAX6qL3HtORnShBfv6MsdEXU3sGJva192DVXpohNuO64hVwYjR4932eWU1oiPdmieR
RrxNiCcieEJ4Lj1yZj2oWS3iuYnOOQKSTw2QJ1ci6reGZq8fcjggDBFv4Y8EAewcAStMzUYhsdU8
kVAKMucWttC9sxRiWinSHTLVR1jjXRauLErVNwSxfoVJw3ofaZmSyVRlwLS9JThLXtqk+uVQXUSe
TuwtwDiV5JUSUKg56VjcfIRM4aWCoh7A8a9w8PCOfwPdF0etjMiUZuuYACiiEewEx0YrYkB25c7G
krRmmoYPYZBSB9Nk+Bwo8UBaUUe5DYuJoHxMBy8IIISFOEa1ynkf+L51doRKbxEoW6yPgHzas0hL
v1r1Z4YZkJaycFZz7GgZYIoI0yxKZp/orQVlaQk2tSLt6YdwWhIiu0OBBijAHRPSq2V0507QPzBv
Vq6XcCrNAyNDikjCnwVk6Rnba/m3v0Fho+1Pfz1mu9y+r22V0UgwOWYXd+OZVH4Hj8Wgna/EcI5l
Bx/i5nDouBF+OeJPQHqHQ4tMnQRGL79qBY4lt+0Efq/G69s3yDGaKhBaP6al2n2UZGg4sbjvheFj
b5W3odn/XhvRAW0HF3ZPqyyJsb8oc6dOTWjTOg4WJkQWrtFv78FJZ3ahyD3yEWwHuiKLe/2+3mOI
F6fpKA7rRUHHPGxRiKwLXfV405vNCVwEJNti/9FEHnB4QIdJ46F8f1tkCPy0Yx7W+ZO1HPJJAhip
FpabDqudY/tYCN88+3QqlRzaAUngImWhU2++pDhmxW+VS2bWWihpizR/O71HiXq6KqTyIcJE+Sxy
rPuKxkrge99d9xmQcGuIIP6DmEbzvtg/oLe94XHcZ2n5eGrpLRWGDZawiaY/BsIhQzkc41+LtcaB
o/joxeJeKfifvZvydMokw3LJzCH66t+wNY9pbK0YcMXI18lWobKE+h/q/T4KlyZJoZnnq0s3kf4A
+eTkW6ZGsgwq04zpeZsspce0LW8l80XLVGd3SBO4N1v2gXVOVgweL0l47ycVr/1m0LQwBoHx2kAW
+7KE9/EKC/L7bIZY2Vx/3OPMyexdH5P0WWwfbx+M1yZhS9XtMeN8AKT07z4UrQdV/WueykAQjcju
v8UJDN4AbcTrG1QhdHdGx8IRQR8yK2t09IRB+P4nJCT3erPv7yd6zo7Gwc8EGCLfHz0RG0+pThnw
mRglSvbmQJw9lyANkSM1jkF+NGNyOqeGptqJgKMHVbWOLeO9zEcNRkS8wdg3qkqLd2X3piz3Cf6/
a3/YOFAi5ArI/6czTeLQt0OWtb/RPgSELVDuLKZRAm/RkNERI0+YkIMxuxDP9MsbPsOuYBsQTbCs
sEkQ0vjopVzByauD0vUbZezt0OyUssvPS3e+JFn0MZn0p22DLfcoIqbVo7rGGh1PtoZWQVUs24VZ
CFDb47WKk4txQ64q+ezzCyUMVaWoWHdQRqubjth1bkkiuiZzooEMsS6AUogQnfil5LVVk0sT9Ajc
KiXeWzsv+Yc3BBRL/9vBPJGZlEHZFsIdA1PudPCuucjFFPM4WY35244cM5lzvqnCSCup5iC+YITs
1LWJO7eck++CYIHjbTZx89TjyRfRStd3relXAiICsqDz7yN8Z6/4L1G8/s6VaXgiyWrO6Yyhlxsp
jdt64OEvIQq9xzUn4TsDyGdFk4Es528W4wjIQa9+tL9X2BgyYddqin9+BvvnBE6ytKG63fVBf7kk
NPbt5y8Me79p5kAarPFwgQ0XitUdZK4vvu4bVYYSlOS/qNy5bIRBA3vLJEXIPvrBDwLMgLqW3IY6
5JdXt+ucrq3M3RtY4zDwI1obuks5VsgircLBtWHrY6/JsMb4njPhQaOfPX11lkFpjOLm/UPpWE0G
p8fU+wQ005G8MOMZNhmeTKjniot+tvAR0Q5t0olGiVKMKKdiBBGiU85Xyw9EhQfzHU2fEwb8L7x+
5Xhcx/cCudfy+J3bWqkEZ4uaWL/FlDc25lGxxzuXEjwj04EOvq882qO/W7UTFQZUk/piBjUlEqjC
CBzqm6+Uq3IcG8xxBzwkrNvMQVgby2qQnsTKR2C/vTxvSaHYqAVuYW2ZGry9qvgKBK7a3YDcLChv
Nl/iYF44RHiRjnabPMHFs/ZSLoqPGVH7e1MzGWvJ8ERvFGzd1DJ6fBtrjlqutGjB+0G0Qkb4wyT2
ZaenIoOVWdNyDRYgerGEF+NnPJmffJl8400ptIKoKUQQ/MdEri0yzI9QLTLLSOPhqkjvVkrW/rlB
cpVrQnNMe3P8ed/bn0aWi3fZRNxDItQTR6Bzw0UTsmWeM8oIH6BurL1Ph3hVzkIcbGJy6A1knxvU
AX9c4A/nMtd7Z+9yd1jOE7T2Gw7qo/2JEVp7T9DKDSBj3zsp/kUOHLmK/MQjdSrmUU7jekObsSlR
4GzBFrFbBKZApgSKprFjQ9XDHS+lrwltFTMY5H0o0vA1Geft9LYcELJx5bvivKoca9EUTIfLrVhJ
tV8N59r2sqlcod4YohH3gQB+tUIEOMqfxPEqLzYDt+DbpS4ieYPI+LmTj0on9f2eARhlDGIL4Z8h
Yee3nOHCwO3H7V9JGuiyZ3P8CNGUW4fb6JWoIxbkTEP5hfgApvULcLYuC5TtSshy+uZj7mE7mF9f
0EACtXMue6cQYJLXAceQRCWr7nSoPwUi3L2dI3MoIYYLgPfb/h/HOeRw8Bzv80A2vPnmdkHiPKzL
pK07KOoKzZniMZPxIi2JuPnhgbtPhn1+zGqtb11BLPY4a9x6LcLZwNRWiGRbea/Wv1v+muAzVoDT
9GOwotnP96wMuQBXnNTetW5+olC4SVjsHc2uM1rGXo59YMWr3eey0Ew2fATcGuhsGYSVd6NrLp4q
uLx9slA7n23OHI7Uw33BHdX/c4GsBPaR2EDp/ox8vh1XfHC3nRdGebdsPG+dU9xUI3JRPdHb3L/d
K1O+vBExThYvj8euRXyYUewfTVOZTo0pdsxh+1qA/RiC4YdYPWQvCEqJavYjWZ0N1QVGd/naA0si
/G0FVXmDpEdy25DQbGWNd7BYCQauah195jRSpVMx7IoBaebPaxnmn0KG1H78ntBQseZNXoaAGaLo
G5VwH1f5+5NDIo/VdGgWkNoZOHdq9DGhJcWJ7bEViiy44fPHkzaoSJUh2MfrRrdT3HBMzNe2SpU4
IxOQ4p+h9Z4P978hAOzDceZb6DcYKIN/qxCnm92hKCL5BpKMOlsncw8plL80DCuOKVnDxdw6wH4d
kW/g/nAMfLf9TDF+zjvTjUAPdcE4OW8dqNbLnLNWfP0lizuYjPrdBCx04kUw2NPKr/OULQxapUzG
kPxVabYgbIpY0WL3OQMTxYk4PxnRsoMOAPiBni32Usa4iXDC+5CUNdGGwO1xPbBs32Etp51GKvHi
k+MULAdPduX2rN+8Uk9cGk/LVsAIjNX0ug9AR8M3nEfz2HNRWZu91/kr6VtSwhF0N7/aL5u8+7rc
bxHTmEY6Cwu7j2JkBj6nurEzvr9q5r6cGhIq/ZKwXFI7dlaz1eRuvuAX7/b6eLlfpJeo8ADMjTbx
Gtb7rI1iVyB6pOrPdDeUmD4r+MhBTo1sAf/A5I8NqilcKbtRMi3Z2enLcLG6eCJ9IEN9xwxg03aH
AH+RpsVOuBMqo+RQE79Hmja0LyZCmSt8x+3A/ZAZL+XtTEx2BRB6roGKJC60b07evohL6eVJCUZm
q0XMwLq77zjHNPJgizz34AwZPsCvw//OlEQOUVIS/UDPEdn0rtFZ6Lo+2H0XLeBx5mxumm3ckF0u
0nW0ZS7yJapzw0IO+KITAIr0Z7vjHz30F9IG/6+9NBi2LvOD9hDEvrydU9TkWuqsx3WZtYx1CxNC
UarQI/xfW2pf2fgVGLO9pm9A/XQqrxE2Iz9B5/JZIznhw/rjKF3QUdM4J9CHvXNMG9Xo+3TIYRdi
Af1GkrqxOxnVPo5xzIZQ4PtjRwsWgHLimvDSHT4cKKxxq2hDegAbrE1iUS4YHGavo35bhKEZ9Weu
rBFfF/Z2UN4JriTI30hxtVDmjelO4kXjC+INmgguksXVjvJXSEu7eBgXDhMTV6tIvgJxMmRGm/S0
pvo13Jn4+aoqQwNtQchKx4LWbZy0b4MZV88W9weT2Yut7cvvWVmRI6vhB+pmEI9YFYGUe5DX6N82
zZUtBww2+8vAgU0RcehImflaMaIYEPu6Xx7PVt6s2wIvTJeyJwxAHB1v0bf9SGa9e0O7qqoI/gCO
ugG96coMuzfhVqiu6bBa1XFwgmxm7+04GecH0lKSzrDkwAtIAWPXv9DlwPXYdrr8v5x4vcJKsy6c
ueuuouiZRNG5/VBIb4TiKuRFhqZ3Q8m477+NBDEHrDgG/VKRd+U5cH8n4f3HVs4oR/rj6APPefZY
2LT4LN+A5H0PQ0ZmibsjrWG4SLFWKFFNqAXbrUP3dR/x5aSFcWso/+N+XXOlqoH4+xhyZrW31cZP
UxnNIfPB9xz8MHgtVF+m7dIWfK8wtYhYpL9/1NfXJAvvmantGC7ONQxIjiYn9xY3k0F4gHEF6o2Z
S3Q5AMZdE8lb+j8NoZdCtdMuz1+NT+DTSN1ctiggOQawByRrglat4NUzV4TnTLMpAsjeGSxWxDlQ
uYowqr2FlCmhnS7ac3p2diWW9ARoR91X5OL/0NC1JjPxmrv+xCNm1ZxEhxNLtMczTrJ+Mbj/Tzjv
iJ3tHFr2G7XbScoEt1H7S/8tMSA/8ZkH0AvM/yCk5VkapisuvXqMqIc5EK86yWYsuJBP8qtNzQwQ
yb0b4O59Ag8xII10kWWq27euC35j3AoKW4raDFdTzIiBC3Ajqrr9FVLpBECXyn10dMKHUUPrTdOK
5AUIdrsldKQUgyXcHVYx68nI3Jm5mI02ZIp55NvPyBhC6F4k0saFcaE0LKpr3vX4QoqMUSQk4tCB
7mnJRsCMBlVD9Or9BzaN7INBYqtm03fmIKwoDE5HKdTjkjbYARTsobr0qC2aW96bSMazo3+3WZ/s
abnmU9tSfDiWNlJ4DAPN8i7lfJxX7woLz52Fj2rRMb41d14l90p/szQQE51MhrzhTKzgvT1tM0Qr
tc0VI+7P+D0zl+9+W+KwU4UcmghgcuzJd2z+HrUSObuhkX3Vvy9R32UF9EYXSjk4U+BdVSQsDtIA
DfrBhi+kw13zNuM8W5ZvNnstnsFUC/PVRpEBYgUEBonee3f/g+g2ijH//K3M/Z625XORQ56ZY9t4
ZoCmBMCkD2IfPI8jOGvQO8mQlJylEG83kOt5RpzIhM0K7LIpK9LgAcw72lbblkhWwxuBBJm9nF6Y
Vx0axLEVOM4kvGNaHFwR9u60wfyG/X8cRVdO8QuWnFRG1QMWjOPw5wDOl2A1pNPqfOL25KEnMDfz
eC+zgKcFiTss5Q2UD/bM3Xf3OXuVUaduIkE7cmxenhK6eKeCa0opUQlVfuuJp98evF6Up2hcDTf0
Z3A1denCQaxKYJZ63nF0NU4hbSaXXmKC97idFSLfRlFXBY7oIBkmTTzyvqAg4vTTmlnnadUcnnMU
uRFF1cRQwNgVqO+/sIehup5GVVq4Z1TqV351dlqQUdnAGGdmNsd8CPAK74mbTPT/hjJ5GMaFfD7h
8obT80b0BTIo6za+BwNTZ2pUL2hQufJfw5bM0uxRk/zSDPcAF2AUM5w9aK3jRbTNmhD/Cfe+qVZ2
UZYUTwAEkb0W9ytXiNHldbmU/FGF7U2Deahk3i+b4pXf0f6OrzqeGi6m6ox2WTbzVa43ox1BYiSE
RDHZXL1Miekkbr7hGtLYF+vD7JsvHVYFmr0/Y79nI4GMG+56QYGrVsaLfgbVnkm+6Rks8+vI/Zkn
Zg6nPeYHziLQ8Pk4HgFKldggQTFmZGpM9AMZ0bIWm6TZBCDEqeLS3DL8hF9Ju8zofJ+cOeN7ug33
d9r/9Ct5D+PHRFmrW5mXpjWy7+9JLpmqPGzW13/6Ud7+zbEJrV9oiJg+ftRJt3uKZPOnpOfgtJ5x
RGB0ufLgNNDh3/It7PYs95xj1hovz2wVqb4ss7mpn00PEvIdpOJhwDbSnihDg6Eo1nb1B19gvpcz
NJs1EDyBulhJwNfcdNmMrjPLrry/G3T3XKZc5XxhlvDhNTAwt0GZDQ9ymrEME/wnv30V5tZAHivm
rOyKPuGl722SCajVL2MievxxYfjknGelliRXi8VGDM0T5yr4N2ChAPORkHj+6JkMmvVRXzTbRokV
7uklXx7wfmu7C31BIWS8rnMl++SxNRc6SgamoFiYnswR29PBo2dQluOAFzuAsy+3Jml8JlPydnTl
/zH5VlAlE5zUI/RCtRPYSQtUmoe2BIliVlKCmjjcsZatlzfBDPLqrHkGGp+2B0P20spZU79azpNy
lwPIA946MafvjNUMatvMe909qvCppmxBrJZVK1ijAc5qyrVHMAO738JCXVjhcZLSjjtjkCxbPvzQ
RACywuxESZhCEh0sWTeBEXOO3yLESmXGJxbNrCg8e91MwlL6OgwWfaB7WbUO2zPrghQq+v1bQJcP
PDiVpE2e7CVbKOZx0O55hRPDIOTtN17jtLYWtW4/SRVI2dHZ+gr0Sn4bREvnHzDS7GaPr05buBBB
ydZEnjrEhMcxZKZLKw1tp6yO3UQ1aZn55wxGnoGSe05uPJ8phuUeTTUAS9AjvGWaA91/MNDJVOZR
48R0TzSN8QiDolQWoyNSyHzqFwdfBPZTUgt+GAF8msjQ9cqlUHOICUHyYKA5UAtsU1QndOejz/x1
gVKuTor+iFO+349smPjjhlEuQYdvmZjo2Rq6hYX+he06MfSLHgIFhTiIacWN1IrSIGInDb8dXgTd
QuTzRrRTXl/wiBoN2MFyEF9ZQKAgoCGqsLxc+9OukAkjosTDCPpXy0xgYoNMPQ5Cs8QgiFOwBml7
tVulZSdK/+yPQxB/klFyhIojt0wRg2KRCjmpljRJ5CyMI5HxZMDJQ6Ms7vljEw7Uno+W6KNNYRUK
tMGFrVN00QTe4OX7U32ctA8K3suknKlGD4s6CJVy3yvfxdfixqOOzMVp9v0grFytGF2UfNErYHhE
ywP/GtMct+JB1ZSysweeIn3QFChtJOoyo0+dp/1RF3SD86b9R2mUW5B3t7VHzjPnUV4d1rGotS/+
v4TkWwwaxaVJ9J26t4powsUXvo3ghiq25BRq+yHVGQzhS20RkkACCU5zYQrovP1InJ1nAl6aQQ9d
+3VXMfWMhm6pMFbHUbLt5sKqBZ1ACrLGWQNKsbWwUS8P4YlvxITe0LKo1jbY9rn4qg1cyJnZr1xk
fMxMoKGHPMUxYQg8d9Sp5vavPG/Dbwfbi+6DI9i7eVOGj/rZ9TKwpAt7I4wNj4HPRYEzAWbKM8KH
wCoGC5WIfEfWXe4ZcGflXhuBiYAq8onPOuDXEa8pm37gdROIUZPCmcVOJpDYkPm/MnQNxGCsy4cM
ifgFzzBHdAEKIiKebExWxH//2kFau6QA1sa9oNvJzyMKXVMTV9aHiDbbEoCcWh7BhFTIXcmQmXHW
fa9marWFrzfYOW29/rx1YXLUT81hgoyBRllKOij/k0Q0J6RhLqAyrjNmFi0KUe+FidEwFcnTEd1r
bBEcBJzMHeZR2fYSwpsQpS3WXaxM8247TdsA6OU0bHHwdCN8/xLU7sF171CAPhRHBxXYs84kFS24
6C9kJ3B4B2Qh6/DbsUb9REDWN3BM8+C6RYopeClOTOfikpoFlsdq3Hw5yNhoOTKCxYV30ajfDkLQ
3dH+Jqr6rMwUzk34BjFlsZIgSU80UU7+xL61mJJI8NGAHYxqkbomJsuFSpj6uAkHgj+uafDBEwoS
jvHpI03I4wC/nBhQ3OBYR9rQnNwpeetGLRWRtHbxzHx66ZhvPPSrO/YhEc7vs3VnYSbjoxTUCkO4
ByO7AD06AT4OdStBNycqOEuSgCe9cGEHFeZg0iXTH0ou/lz6LocHUrspKQsOj0D9Uo9FfxQtcMD7
HmMdQBTIiNoswEFSEURV4SNPmSUB8AzXzStc8BxWT5lTdpuwQIl7wrwtHQXoJNsldw7inCU+EN4f
6TkgB2eA5ySZ/SpdF3Rb99VcCWO1B3byTVQJYbcmNw3R6YSPD9/Uk0ovN3IgkPevs63mzi3o+lz3
OIAbgFoTqsEcmFWsHgnWwvg5a/QtFkSl80UkP+739WVpbSU2f6e71IzZbUhoaluqnU9Dbvul7SQb
JiH8WV9WTIgRYP/2+1y04jHz/1Px808p3GFbE2Flv3BpHYQP13+Ylco5kn3NT3dGsKUxO030tmEV
R5dtnRApmooFjizzTZOw83D1hhO2w8Q4eVqAzEtRXRx9moJIpdf8tAUuTWq8ecytydIzEhfLP8Ud
tstyeypnjsM/xjgZLAcDtpKxwlaYLqC5bcLpnwQbFUfPfEzIMA5tbxIaLB+TcJywNerTJM19whAE
3tpD+o0g3XRWmiorXtQmBMm30fEMwGRVY9uJFSNRi31ZccTEZO96SklidIs18dA3KDo6X2S7r5D/
zr3ratwjcgX1NsLF6AryHRFwLRyRhHCzAQvsX3d5j/WgNXcSPqphse0yrf0QPYEKDovKhLsNSLRt
N3YNDCxY9fnmOIMgaR5Isu70gaTaSzCAWdfOXfH4ZR+LosLQX94OFMcBGZYaCcX9yqw0E4qixvdD
3GV25STHiRBKhT1a098jP+GyQIXI0ZN1ccrvrC6yrtguxHbQH8vsy6qNLaLZSiWkp2+GR+YkbjOr
WI8xWjX1x/CspLjgAMJ82KWk3ZELjpUhha6PV3cMTG5V+jOWyiV9tPlt40fF8pEVhxwvFBc/OkbP
ggyu5U/hNNkEvkXSTQHTWEinFRNs6PD3JzFTE8X5QZhw1NMmQ2AFQ/korw8u5SKh0xlmILxM5Sz5
RXp9tvcKZsZfobRvFyPwt7WFhLCWoniAtHUakX+cAe02debbfTYx1EBuru4ChrCxlQjJLkCdqDw4
Cexb0e7llHVpxj6vPVXSPECkDzO71WmCWiVX+LcYmd6LKl4b+g1lVBuaLIMdXXSEPxjnBvVt5BlJ
41veR5fPIB11ngHHg2L8gc+k9emKP1Btrwsyj+T9ZEzM3wsqOe09NGiFn0CsU750599fJ2sL3lXb
0YzGhAi5S9oOLOTifYUqZIkpkNvJQP8umGDalxLFhonRozNst61as/ULrvuc3jceZkdPktgXfFV3
aaKth1X1+upnpisU9Yp0noZ+VEewZEaNUAeoZLiB2srCNbQGOZJUiOr0AH/98aHYHt8OxXb+OSnh
vH2CzvjHNyuHS9sK+zrDkyCYrGKCXlqFAx2Iton1oj8V1+KQIh65GcNz1uwRoGGmJQCykAPdgAhE
tL7efog5kX5FJpM9XZwWPTWr8Vj1HHi0yodInVIDhw3VKV9ZOn2X0qKwPZdlS/0UcrrdHsN/0fLw
VluN8Wp37gde023p//GSCY0geS7tU0YS/pivrvF1vt6nk8oWbLLn7cJvodpnweeE+wJOwmXHowMm
LJ9/Ck1XtCe69iHFomjfW++5UdR/dwKadjw+gVFmFGq32plD9MHCa99dDRdVvSeD9A+yus+SzxoA
/84xQ/jxi7SlOed1oejyCvlmS9EIdmgPNleVy+xffzhPg0AtuHTCfDKHuRC2unpxa3R4/kQu4Vf3
16j3P4cF6GPvT3VQgKlj9R64P1+Ea6f2/I5iXnAoF5tDQsQHAWxcMY0prw0hCrApW1dAy/0igz+7
++qWX+IpIwvgxRiuG7/BJzPhgkNfPBOHVYILxtcDYdsXYhS/ok4XsR0eEmWOYa0ngxu8H2tvk/KG
LzyxI4bFzOf4OXmTV0gigz7L4utnXyiD+szdajKu0w41ul6hJjDOEOIv9c6NoXqZ/MSHBEa007Sq
8YgfP82OSGADzJyelHhD7Xnzk1wcdM7XYnQGynIZEG/IXNxu2oX1Qr5zZKGoOApFyjOzEz/6QKUk
XsP6bmlTcJrYyC9ajy6S1TRj/TLQdMPETugZIuo1RK2SbCH/rrh5YF+O/OfXVCnvY82LfL3u2YBh
mvgvtAIrXyTFK06kXAIdKQRBBxeadqN9ZdqdYraIZKlox2WqVdBrZ+16qvxgVKun1m6v2WVGq718
w9aRhy3sv1Ty3kWNoJWATJrof4xWqerRdO2Xe5lVE72DJLb3pKhBqhbGdTIb/9+MzGYfg2rs2dQ6
t6Tcpm57d86kNkDmH4WV8s1xRdQo6wgN4UA2oDfBPZYOGwHo/NISHk1yAqmsBmQdO1FT721s2Qty
CJJ6rCPLWgG5eO6UKdumipHvJyOBDDSEM5VXSdDMgi8qutT221WR3/EmIavSTxQVk4n1vp7V+esF
ohjplY0JIE36zK17YgbKGzNxSeGO7tGJyVB7Nht4Rm/UoP9xBXArEKQmXGkHx5J95DInAxlyyb7Q
+WdbLw7MTA1fWXUjTFn40YtHr7RPVg2ttGwJsh1sh4nf4oe8MVtDN8zLWCGfF0ZsgAUOKFdguR2w
hRxAKQamVruVuAkH2GHPqPtDgT3VtImJBWl8zHwfGQowgk8+EgK05l7miRx7gcXnHIhH+H8nV+Lx
IJzyuyN75idjVvQd4kzQHzmi/s+69aplAnyF91o4GEesgyaPFqQ25cH5BSMJnx22BP46zOoWpKDJ
67B+9y+IiyDG0cK2pDebGsoFgjDCgZHLUZrzpL3SY+FcpYeXgaJoiK0nr61i4mOQ+SUkguPp32T9
JY0bvvagqOgun7gqAJF9GRaGRGJBF52wF92J0NpICKgAlC6Q3fC351lSImKHqrwuZ+x/gi9Tq6jG
efxAa6IhnL0hNGSmkpYP9G93p6JMXaphzo1wWoN130AVcfmWUBmHSHtRhcF8RXKp1ASlZvB/tMbh
2jDrOzgMIkWcELzVLL64e3DnMdfg87aUSbJMqyJ+WoCjrbpVFdggeEMqRgVf5vfKusydgwkx9XTE
MB7RkQTr2DaWOvFEEeDCBYRylCbHo+Y1RejypqneZhXAMOWE4Z5BFrFkTxcdQSpR/28gS9zzp9j4
RuzAfP2kQsQQEwWQAL8HzpB+ODYrSFCW6RJba7uFTKkGEhNim+/veMtek3vugamWF0p84LdlbPmS
IdkJiQyjdJClFMCwFB8Gjiu1mqmIQyOCnB6CE1Fh7GeznMskNo0L088/wytp0KVHNOA0ktrOYF2y
8MqQKM00WQGd6NvyPCdqRZHkR/MEXH/UmcsXMN9RnZJ7X9nmkhX6KEbX2R3ERVHkE4755MQCiqJJ
2b1++Sr9h0U1BjMRv9gxiDRpE/j9h5A/SY0SGn0+hcLZq5X+NFLvI+kzkBoal7XfN5Db8cNjsevi
rYIfShxO2qG7CBv2GmruKg0S+Ca5yqOUraicU7ij3nlAoIGa2Ekt8XFk2yIKBlf6pA7snmwmNxmt
6NVvGQmQBXd9L4sCIcE9M4Bt8iw7tFDXwIaAUBbBUyIYGHy5DfJgoM+LzpEUcAwr74tuGRXj4RnN
04jko5udJhAgbfZjtH/5d9IBqT3pt8yn65WZaJi/j10DZDRrQ/+asAskmEjsPedycIhGgCxcXipf
7Rhu2kczHK8pcHwvmoHcvUnYLdQoC8qOv4m/s4AIL11FGU3cuX3FAIxMqkDcxKpay/bwnEkTqJ8b
CAHpdSbE7btMFd7i2UIMfHrLbog8ccol13bCoaH5yKU7pnXKH8AMXLKlp8goEP9fnVrs9o+bCDp5
N/tVgfcPgN/eqwgIIFh6pEhplKxBo0sZeJBuoGatd3CDelbHN/kPO/q6fwW5iityHMbX9gc7PynQ
kBXTMwGKcLrTzBtojgXq4Ms0wygyG/pDWjjn4O9tkiIUP0kZYjLqrRSPwuFQ6PT9uSsYReOJ5mUe
QJ/UdKa2rUITUaZVhizl9ekEqXV7R8qZpuSCaTUZ0Vi9HGXp0ZHht7SV4byppTaWllKhUglet7Or
0ZFUC/ueK3rmkgSoJEcTspeJDC/WNgZG8MXaIIn6Y5zNFl09jbIjt1K3s3SFhSyYwk+EBXhSfLJQ
9LcTa34vlE1Kt5Rcr8CXB5eGDRhsrfF2HqoCZJ5f77FUzFm7lNT2DfR4yUa2/X6clrgPBmBFEwlI
f56tbTXIrK8GthAV29tHza1DmG8I1ia3rxRxzJXW6TZSbW97jVxtfapCI9DsOBAip66Ztxs6m9Fb
+dHGbilTwf3FMWoQfRL6kAEXV1pRw8NElTNJNWcjkrOXlGto1RPrdzB+rbELA9+3upo5PRORNtIw
MwAVD5Q3kyq6j2chNsS34uxHWZtOhveLiEJepromg6I/CtcA2bq1jH8EjzlBeRAASjatg7Hnz3BA
gSqAquT+nRB92Qv3FksNtO2vm9JdyfrIekOWGmAopIaB20GBtfMm9rBy/Ya2ommVT193P9ZdJz+m
YRcP5YNd5WI4DmQZzqr/AHk+IF93sFPi+X42ypt/9Aw9Pnpv7EW+yGjxa6USpy714oz4O9kYdCV7
qD9DLyoh7K+N+CYAtKu87HbHdcxO8tzLXpV8p481qz0/41UOvOpqYWcFVVQYX3wmn5YFM2ygRJKH
k90aIjMIyv59tGGK+gIiNL8H6kk1F/yLb+FsAE951UuLWTkeVs/dcO4OFBNQHU6rWr2VpqfPIU85
iNHJHPWsFQfg+apE9sNeHSotMY7klKgBus5KGJSCPQSTryhUJgVjTdxWpBl2xwzuBft0pSUBgRiv
OTVwT7Rp5DeezsPq3G468WqY1dS9PQmrYCT9jNVvEWSPs6Tc22dNADfGEDwVi/X5PdbLoW3b3WHG
7p9LrhOUd3GAqb9L08lSva7x40HnAwV7fiEo64FNW5Q2ql/yFU1/coohzk1lkEjAka4IJpJyQS+Q
VkgvF9TXN/YepZD7oSkR4qIjlaK5sz9YLWipwPqspZbOUM6HHYI1oCWM45349D2gtuvawnX1FO0s
5PwOL0A4HEY0rassyKLkUGcnkd8PW9H+boMhAbUdtCXIxJS5HQieq6nOKJvFEgWPMVoN1n7JBy9q
kBKbKTT6t54eGGF94chHQncaakQI+Y0p23jEBCCg9LTDSZrG4SlfDoK+akAFoHW03B1dr0IiA2N7
9qEkjK5IXfAVkJI/qnart3wcEjUUI94TOnAXxlNCNaqe+4+EIC5s97S/8OgsS4X14Sztuw96PveN
Rc8elLqJ0buqNKwAIiDyfd0UKcNP8u6JvblPPnREourot4DuV23Vn5r26BDnLrIJry961/adQTmI
GSl+uBZkAzL2Rsxjbx7qvFcA1c+ca1dIs/kmS/YhQhwPHtokXjx87ldBfQTDGXtFFX6gSpYdEezX
sk6RI225kga93WNay0vU6rI9iD+iT+cBOcjtuB6Yfh/1tH2+q4lhcaRn5McrTMAEzjbeQuSZv+Ov
rx6elBrJyldid1QZKCw0qxRwJ1zT9D9ufjjMOXTLEIOSIxvntvmtDCeec/taZim4uPL7/FiWesLI
HdEKi6S7y2eD4FtLULhsoA1a8cpTXmnSIo8ZQSUs4FyElyq7XsilgygoVFUcPyEZgO0CyQfYn37+
/jmUDsx2aOX3fIsXTcyQkYRtYI3pdtq+WJANswyw2/DKW17yZA9ReOVNP8lhnhXJFi5DX3NDroDh
tCMtv9nwmh+Z4JIFKwpgs7VQP9HgL+9MY3Nt66XXErpdrBjlt4y4kJ3xQsbwKGTOCw5JEGkQrvVo
461vKMevOiyy3JC9yr5OQPwRtZ2vjVjpBHlLxUuQHbtN0C3uPZDwV4IJOKIz8jehSIgr+yvuSxqw
XII0eUkUhze90R9oB9y1eiTOSjhzfKb+XE31vFAp+GUBdOSAlU6FlnqlKr4QoTlT8G+EDn0k2q3w
i83pn64Hsup+IF5pkwxdFCpQ4FWHVai0CiwP032Z0x8Ywj3dTxJWhyCrhgfIknoSR9uoB/huk9ke
aAv7EYwCi5Knx1J5FVHa9x4ydipTuiD+vEaH5dL9RaSAkEg6lLshwTrZ/J5zAgL1+Fl2SSACs7CV
r7+yZsu2AewfBfJiI6LFEowoA7CMwZ5Rgp7ufWFM8djEVz5puruLsSUAoIqJfMdG1oy9noftO+v/
coVivhRBWhkcxc6D8LdemxTExNGYl9c10q2Ff28X6fWzaD4DM8/bPsW/FtyRL6cponnrhMAlFX8z
NsvCfMUHD7nwb0Vk+mjz8iBY8Mc3kbIltZ10qZq+aw9hYzOlB4XnRBA7IAWs90+/QmcfC661UkJC
yKUh6uwXjnijJiOakvYQ3EWF7FS2T6gqpEKxgDuVhO6AIOntLx48EnI+b3lzxbq0h/JK3M7oTE17
1cC7XOaU114DVRuXW73Lbk2P3E3dGKvcKjBON1mwfG16JIirKHABehvvsj/7F0mFHG3yPQnvnAsl
pGtzrET1YKYTF1kex0Env8LY/pJ7UI34/YMKBExkbik/ttyxY/x8O29IXFAPx/EWogYCY38aMkKz
MH1GYKvLsoIO6vNw0UaId4romIeVVT7HuVNVO/+CUNy+XRf+7R1bByREdcl2vwUGKwPmPTS1EBZA
RRge77RlryN7qnFqDR/vXcXM3cL2oKUg8I4Q7ReeGnEdD69Kp7pC5gQrFxQeLE2XQB1C1xU0jR6a
cExXAacz9Yhbn8JHDpLXo+tf1QNeL9wtSa44cdqX1nZTazyFUofwgxdw9SjUSyd2HC5b6qtNJuM+
gzxV4NZ4jllzxEpR001AwQ/BWoNLPs4Kwcz5emQNQS+MrqLVov1tNnieHVM4QHYZDy3CY/pYFlno
/rbsBf/FnV1yIBQ5DCBBO9BNM9lf42HSk5ulhz4kyYz2qEIY/mzZK74d+elU4rMuh9N+R5l4nASB
Fj0S2ijFbySmwKeR5aLi0F+xWY9CcN9bzkwSMln9uIy5aO2sKmRxkLUXK7KkWPP9gdXFekN4HHEk
z88W6wTx1BBMdL75a1EL4+JnmB21p3FnPnlVRH40EzuE3JQWfgLaPxKp1kQNLQaYXf5FQL38s5PK
B3T2CZHlwnKjxJk9Km0Yea4piPV7LQ/UemMT9mB7slRfUGlRxwnZ2iN9oCcIVsGMJqAgqxTRXAf5
d6vG/XST1rE7sqvGRaBdxlnme1oBpJ2Iv0Rpk0QjznL2//sv2g8nZYD1P1a6LPici5HvuTnySHJr
ogMv+tncS/uw4ulP99qygNxvvtBPgwBJcOlE7uUSFCpxEXthtbjKNwzXRYi66ff7fEaCkjZAALET
BXOdtQYRth3ARjQ2kEUYMZz5JNfjpaRtcf6TiCxfsB45tJNDHwbvvXjflyameLFXD85AoHg+ESJI
sBky6pGwx4G/BwysnieBlBenEtf7j63QqhXtWPkEfBY9a7Fd9DWpbc95qzlSgkxJ3LoNsM61zbpF
erIU1F3uoIDO8y6J93fs5djsXcLDUU2mD8IUNOCBCFP0uvCAyqpUqIyWHUq22zwrs25XLYhcA2Ec
C2uW7ZQE2H3v9IRShhC7LFpEmRNrkYs+E3XFibwZEh70LLQAqQzTWlV43P+jKT7gY3dyRbX1RvpT
o3reXsiwE4dsddvd8iJvUX2aYuMtSWcSYMxKptQU8BYsmdH2KSmUpw8IOhdu6YoIKvGz7QEq9m0V
tdMZOGLPnPf2OEV8FtQR0ZDMB30UydEXa3UhE0Tw6hNEtIOhTAKs1RvVv3JmRgnMNh0V2KpR9aCZ
f25l4zuRooOCCL7Nl11E4G+o486bNrnq4I5Vbqsi+2PExCctIE7co2lLjeOfFGizZWz2uzFOPLv7
GoucIcJR1FcycaxT8MGS2whT1HbIuk1UfXkVcM1KKdwSTBEsLkiktW3AVx0oeUkNpK7m9/pPqWeJ
ZcLUqQgjDIWM+l8o5Nh+LQvyANvW9vUL3JbfK175AXxcqvRQ4P9O5qnrmnRpoOaf2iiknqIMjD/C
BeizIwKezslli5E6o9MfEfAXliurTV0NLqtwSKVdSRaPYbMJuOZ//OK7FC92t7XBM9JG3FIrwp/0
UegAr+WukD3f+yTZ6VruVVvDocpRelJzMp6xAe6cQiB+0K8mjl1EQ3y3Pv/zPGctgdCBRT0yOSOW
461jMdoynn9kpN9whTOJjZOQYmderlj8o2Hj3b1y7UxZBo1U1hRqSPp6fZN0kNjefb222VWyr+Sy
aIRObRmqcUM9xY2LbkaK4jWh63f+1VowPdDqb7WWxs0Z3d0EPYnVKTZ96xa6djcuEYRoe/vChrku
VZ0rBDvKfj353qb7as4MpwWYduGmxkV6eOt2XO5xpOGBcGwmu/rda1bWaxDs/7elYwHyL/5LPvLa
GOghO8Ux5bFEdy8mBxQLGZA60aMjKx/AOOZOp+yooXwFrf70faIyMwVB2dGdx7KvMF6IgyTDoX6T
SLZbuIljJDTOadPvxOVCtWdlzLtvuQVUMLWAa67UZK9SNEijZaCUwm7AKbl1x/vWt2d/Wg5movSv
CsjC5LR7bnyTsFGZM8EO7qcD7VTAaeL2SrVZwK9N3ixMjr6GJqZk62pM+e84yYj6YsAE+/Hx43SP
Ig97m1otBSbq//fh+CF7Mp6RO4AREjbCkmTQE1YKMfceYa1Vuybumgf+Him7t5kF9oJrazKP30Jc
wfME6FzNAzcW7ngqNlQuCFAoR+eJzPkhb+TpLW8zYVR2bPnwwUJDzkeGhFI/jAm0WKFXRiCT6Mqt
WCzG8COPPDVy6mDVQghVTEIg0kP5bECfFDKknqEtuPAZEd9nl31/T/uhz1a0raTyAJZ8F8fJJX89
VK1/3hWYCuTxrB4K39tcCQdfPtv2e2uPltPOmbNJnaa4YHAM+4uw1ApdL/FdK60JJSj8uBoXFb1q
u5T2IglavZjUIE3YvyAYDhXQbiF3Vl77ccL7ysDF6xv444eFYldpoHv6pbBHmhJMcA28tYCUylF6
PYfj6XFmvgLUJiHo6sjEdLxagRcTLx2aAAZhvQO4yU4CxwIcH/ONFIeqbzMbfWYVmkle+sEpYEk4
nmmbUq55FK9d9+4TqZTih97vkWbyMjcu+4/p/GB7srF2BCGaLYp2s92n/VxmYu8RnsF6/v3uJjdm
VvwcgII7yNtHyNAkUIpzezmbBGvlfXLSJKZt8n5ZmalygKD1PCwHA0kAzz2+CSRSMAaGuFNMBR+I
6Ux6eNmsYBVUXVWn9AnLl76Kl1kFj41287b9AJTWlY93KSQe4oJMefBw9PGJ/qOOm5kJUwsHdEQF
JZDRA3R558DTX2h4FYvihQhkEBUyfolZduLNjg2saLlTmWYaiVdxHt7mmvbHwy9LhRz847xP5eKh
EFrfhebp1/77vaopHfRUhiVDNXQFZMT+jFyixwF1CGDOV6H4Zo0++nzCke0wJxMZAprcUHdotOIa
nFYjRfbVs+A7Ip9XbvBP0mRfFlpwEugOLRqsqhjOcqfme4/ti12HEjHjz4Ci3uSuKSn1oohYwiZ9
wlh9Uoi+XacixewGMbEJuRIZUxmqq0kGeLXJSS9f+cTYU3l2YpBPBs12zxiQzYaHAx5qjYDm9dEl
KadGvxUuq945my80KNLfcNKwYmI8Vyncm72gZaHfmPVpcBe5g221Tk65puYvbStUonR5kBEH65JM
D3G0D1M6PafnP6UtWMXmo2f9HsjoCjZz9IL0sN/RSWEmANQIh739E72KeOZ3hlt6hzdBtVTnxCjF
O9oKR8B1GEBIYyRzugBTlgrEqPpMb+vVbutqqzwFJSkWU+v/p8pTvrL80bVzrfWdDvln/3A0BVWo
mIcEAOBqprkfL8TqHmcEf+rgu+WgunV/qLv77QEXd5YURvtGx3qmOfNobvpZQwqTeiH/hjNwflik
hKsg3SBn7G3iqBbvnEfJ8bisbS+4Y9Vuh75AFQ6W2xilm2qZD3tBqvOHvMg8orW5sPqIvQVOk5Ph
mrhaLs/Iwsos6zT7Vd8S3Nm57/xhAnrTwhWHFzIXI50m4QyreLU+616V6oGSL70zO1eVaNmjjXb2
WFnsEuzSU/qeGq5Z3GpFwV5fYZVmrUaTq5lAyqkdeTEIIB7vo8ofX2GYhmb1yr7i3cwR447H0JoP
hUYIA31G+LSWbClAEpPlNc+v19kyMgd0CTN6Ppk9m7W3O2C/RAOB63oHTEd5aO+0ttS5eMt9L5IC
NRK+8gcf76w5EH+aGhKDsNK0xGtYToW3qPqd2l4We6/gh/y4VytPlq/xtfWuIDTt7KbqaW4z3TP0
nCViemrN0ALyae40za30+AHu+Mm+ABhgalzAIKywbpqeXuH8wIvgvnqBDOEBPC7Y07msHon019BL
gqcmM8zTLRrO0XGCSjVgjgm0aDTRf6LPqwXBWjSpz6dyW3iSPIMuIdnBKFgGmYCn91vGug6sf8lH
MMvSdYQP7GiPjodwTEcrEpkM9ggaZW2uLJM3C2oq5VLIrqfF53XVCx8MJGETAhSp0cp/vCx2x3av
F8chPFQgmI8fVzxBdXCerOiaQ5qREqSV3u74nliEsMK5WBUSborFwYYkFNHWV75+fGQTwKFz5Fni
WDne4AdG7I9T5x7c8hkey6LS815mjFmJwyPG+AY9kP9uVT6fXyIbVuVvnQTSSZADjIOPUvq9+Xs7
FQ7B87GSEGfmMMl/NrXNvyJ70Tt/Ymz5PsIxkvvQVgOSVLTg5ca6u5ZEUoOqL653G4M1vFufedKm
k2eLIe8c8QO6DFe44e4fMRHRnRkWlf3oLTrDKdkvn+ROxDDeAj6PjCAtTtK8xSuI6+xySaSSFXvB
DVw5bWz4cr3zqXVXJROPqpLDP9WH7CWADHmhy28hgZOrRq6SY8Svd/fC7doqK/M3MB5FDviSA9FD
tdXO0Mvmj5vgbCjI1jDkxsmO1eIbjJDURgn1JUIGwn0K7tORvz2LUK4CUbWpcSeqFEwrTJ37F1KY
dQOaUcCf86iJxu99FhReR5fooGL/sKqIDNhGFw5qCq26CU2m10MQQgEIjHjqXEANbGWpBe9CCD4m
D0eDnrsnku0kLSxQy7Hz7H7Y/tL0Jwkp7UVek97+0F9EsP/fEjcsOCRAx7+Fe+pbFB1ejxvd7aUi
+/U8urxl74gRPNVuHckYr6R12syJv/v7RJ3WMvMwzFUIaMrhuxYihINPQW2EruANnyYPTxSjQK9y
x4xmJvFYdGUMQBoWv77LBjePKFO2BvYiAxvk6fo1mFMIYRKcpoBl3eg+rkv6tljAGnGlz+fGKMsS
OX0UH5b+Nf3ztv1NASKuFU8YGUKnAZDdUaPtZvfho/kHapeI8TbSsmKVen8t24KXgum8SLyroGuo
R3Tt90LomQNwo9JSTv0X6pfqH4WlV51DdQ0zRdsXOX45hUCSeFH12s49nrceZ7XjtsksduvvOMCU
GpMAvkLLKUuKiFBc0Ru0GEhWtzqU1rv3CfUBgk3qMO4B/at5R3K0HYw8ZDCb9bp53hyna8IASGuh
jsbUCahLA0EE5s1oE1OqPlF6HELdFjum1HuxGn/jTQ0laZqScVIgB6zjnJv2cd6mWeo7AsxzqIZn
SxbLgyKgPk3VcCF4cSEtTs/zP5OGidBwW47/lN74wWScVCyfn3ceVyawSWaG+HIjETHb7WOgA27q
XSxStsI/3RYTFPsSRSqE3t1PKe3eUV32uu3qf8Dc5tDJ9t7zDxIYuR592OWkVmjFTiEwADKxvbh/
YRlCSL4xayZuNXFDGDsVkPshTiqcaPoOGebz75hKqgu2sMrSb8xT9G0VJCj2fXDVRszs2whdpTCq
N3ikYAZIQcPOoPQrpLPmyS8HpZ/bylW0P5oHVjfiLC/EeCYjsXrj+CPCN7wHFllrYe7Aa39wQrpI
wFrxU+HiswW5NiO0nR1QhcnJmZF0cFePO3LYx/LI3br0bduTWVhIagNRcHhRsMf8o4aJ0MXN+Hw7
IYhqoOdcrgExldh6Hh1CP7yWq8193KoMDF4RlHw+Cg2Xrw5Aobn/GkQ7LFlUzLizN72RCErJn0Y1
HRu534Ulsm4MsRqDVXR+r/6EivQvjMurObnB91JrR/uQ991gdmTrHs3xQMKFTjPmchD0SKRjxjB5
+1/4VPv2KidVNumaCZp/TsfYRbgN92WUCtC6xbZWSTKSh1mkuNIXzTKjVyBnNg1MOBwcEpfdqkBl
V2tEhxIsKaXdOla7s+lAXwUecmr9sxPlAiOf4PwQauKJDoXkilTU6Q1AWdaEarDDziHR3gsplQ1J
KmlgdSVwo6ej3085sGWThPznHd92pNWdX1wGBo5yLCar24x6vxhua+saKakf2ZHDGCWwdkg6rHQY
SXVosNkNlvmoo2diJ8+Abwm3wfpSNLuFJQtXQudY7ut9wQk+aDrCYqmnO1K1TeZsmLl9r+u7XGrz
D7yGYp/Ea8xPsRt4BDI0Cv0/u6JbQr8aCdzE3CxsuUujoN01YK772nSvSzMSA7eEeWJgRVPEFvba
EGxNuebQSRryVp5TvdhxGOQw891D1GgPO1JnI80b0erxA44jU/4X6YhNshWy6mkConN73xg0ChPM
e2tDv2U0aT7mA5IHckVrMRwmJz6VtVBzAHeCVEs20UQrKH32BBfs9/nI+BfM+damQE23KaZfGkXm
PEakciXx+RVqCiq4ggkhFttmldTKj05VWnBamDO8jNv9cigXcsv0x8yxgH1a0OH9aSSO+fejMTcz
eSynNsAmVwrwdC914L33NS4PC+sDFIWcr/kwOB5pjtgvjEdAOoBxyzTBjxI+8B8/Edziy51I92Kq
Gem7V5j3GG4pjHKJkzVvBCx4XqO+nx0iD++KduoSZhKE1CGaYP8Z1r+MOFQezYPZ7b407pCwWM3T
D0KDyMpWV/AInSt30DvXvsTnLe+L4efnVAOqp2oeLTj+WvBFUwO1gD1Pt2FMWSUX3n0U3ZTnhkuB
NrK9Pyx3fMlLd2W0sHbL52pukvXeDO4PM2L1SJwL4EKwxQGxYpaWXBYqka51idtI2f2/UOklmGno
6ZgV1NW3bBhysjVgC4yY2xEs1DVb1vg565VZVkB8KyKC0E3AqjPgvCU4N6D4Ise4UahGTQoIxPx9
sZIp66jC639IgGEXOAI+IThDjO881m6fPbAh3gqvv6nMdOY8QYLyUYTQXTYiqf2AJydeqR22haJI
cbN3TeD3KmYr4pbdEPr3kw8oYpvrGllQexnBNrjiUXC8YVWFssVqmsEsVLr4srjZUaf4iQ3cPddj
Z1oOi15NMJowpmyd6IlLw3kZWW35OsfV7LwKb2CnxdhIGQtqo5btBu5vQB80UsPbwnETK+3TwPoo
KxAAxn0G80fxdGFs1Zzj0y+Qy3tJ9vzorKEkwIC8aCmHflXMcEJ6pWyKPJoMj/xHSuCg6BR+by9a
CuSQF1SU65ruTbqZhlSNROO+9jxEWBjSf+tMKzkOnBQYG32NvE5Fu1RociIwkG2CbFtRAvvop5ha
22YO6f8yanpyszoegx7P5rxRmOqeulAtEa7KBFwj5oetEjg4eUyQHv58jYgJFePKIqr9tH2U3TS4
Ni9utp9p6Qg+LdMc/cLgEclHXQUHh/aaw40EVVeN6wg27ORn3BF+S+pUZJw0ZpGZGQa4PdZrgzVp
skuG+biDQUGs5q+WNqdh0bHeaMI/efhwIa/DI5o7a9T4QWBct2E+3bqvextlGp4NjG5xjW92yPuX
iQ5xcbmrrIiYBTvzDSU3AReFk9BbLjHLSyV/XIM4xKWKu1QUfIU4iYSMKn16dBbGvUzxBwW1QERE
9vgjGQKvx80jsQYhE6KTb6h96V9l+MvAxi7akRbvgubJ+7buEHnu/wCYxtSBe/wiseTnGjGDjntP
QKmy1LIaEGISIUCjUTMSJddhM5FyJs9jnxjWOoFSRxf8TSWODU4gPdVHLVfwds1OjGicARkvfY0r
QhSYPHfnUBo/RCYqKFOqhsjQL4XT0gEUr7MRhUEkkXqz14ncljafO1Mz0SR2SqNSEiPsCEIFGFPA
sUlKnNwTpvHrRQS4CORDssUB2C5vyix0Z/jkh9S4cDmfSkqHq23clXZTQtRQ96hv+GKM/7TFKCFc
zCEm7wYoxbBsSWIYFIAYLyo0bLpesEvQk6TdIQgZ2LBfYzMdRv9So/kih2pJ37KAB3XahZLiFofV
8xzpzQIe6/iXlnLMz2pELglM155CStJuUhN9AWsWwo0OknkFh6Y93SLGHO6UuAUait03f3HQ0rld
kabmfUa4ZjwwED+eeByf9+5wxhYkLjRN7R1NP7YpsRP4lCx57PHivlGPDdQgXlXU9qMGn5Ll9Noc
56bH8xUlLvIluMcQAsl3RnT/bz2VOxCskZfch4tMsp+SRs4mKNj/hkDqYbCzUoLeShrVUqtYb0xL
gsBLgKH40MpXcyPWdl3/jUGUKTfv8KKroTe7R/+x4TXm47tEWNuyvLp41yUc2GaxaJynnbfVMnyP
Osp8ntFBxVv88zlSP+Wu3Ahg1mCOWEuAFZROoQ9S+pjc1fW62rGDSCE1tHE4dc6svuHLvOlebCIM
eeT+g57hZQQIcrFTW8fsaQEdRwYxNvfammFMw8pIrKdSfWEveMh5AaRWNXOrf1N65MiDUpEmjiqb
tY78DMmkUwY9ixgJk6nL6bEJtNCW3DJ2uQyPIosgN8hCqNhO7T9AaR79jJOTNHnWqghtTi4+XT8u
VFNfBYSlhRm6UGJpTL31j+HjFgtsPVZ70Tmi4tCE5kHKr9vc8aauwWzgk3r5ooUaDayL9+MC3hNj
DzIEZpbUNxakriY1MLwUaJIKa6dSM9MW1xYctbjIdplkSagHzOLlqiR+4xi7KD7VM4+sw+1HuDqZ
bECjw2WXT2UCmel9tCBLYJn+/25OTcuxuwUKNvKNWFGGgM1XkhhWIGx68xFU54fU1M7k4LHcz/+W
noxdk/dC42+jTzdyoKF6rS7MRHt4lxkCChRywzhtG025IU7zpzwGm5EYXhgQ1CnBeF2NqIuq0NGp
36OHBnTteF+yOnMagAjfH1fYF+y6/RJYsLNIKJTpMnVLgE6POTkTkvFwVzCMs94+qcVZJRmjomE8
UjtNEcu+r+Dlwb4BtO6mV8cMzd1QFRz0cOPdXCMm4KRycVSwYLG9T+3xlwcn+8oDYxIRYnoOCZMm
X/aVa+yiWESolvLMTPbg/yETBazSawOkWt0FvTcUiO27dUHBwzIjtkVS5FoyJwkWQ2uRNljVfyC7
Q2n2g7y9G+dEl5yNQ+ZAqQ+Np4Q5UZGpa3H2gSWd/+MAq2cLQFbTL85nE0h/O6AoXsHbu3Wuw8AE
X46X4p0SrUD8tomFI//HhfFqZF/Z2mMS1naTaReddPmyOi90OL+WAY9yJJlyVK9wo2K7qK336TOS
tbGnXmRNxqQ5juoAXvlRrC0uO/MipdV8k51ND4L0ExoM6sbihFnNhvV0ebmERyNNx6/RzSqTDihr
l1mchCzciyyM8HP1CMfXBAT0RM7ZxIj+9/mvdjdQnrQOjOuaRTUiYvGx2EY7CdFuZOelDuq6aqM1
JWrjTkf0uVcu0aZEJ+9tlDMYfrl5Ri7Z7gdSbmcK9CIBbiyYt8E6d7cmRAQTcQ4SnpkPW2rCBQw5
lIB1f47WHzfud04VvbexDyz6V6rGcO1nMX7ujtj2Sk4s0ua17Hz55K46WxPljRo60dHgCVVFIXul
JT+8E6CEP/u3qaTqphnGjeBKwpIsjqve55F9KSdP5cdzEv7ah8H/tjbyKYlthjASB64+rdI7Xv3s
ffheOll0zDaVupUi1xRh79pR4Mn+a2IAU/upxXk1mv/jrxk3oRQUjwfgIQjJeXL6AaPd9LBXYALA
TJuBq20oPmLJBjUx5MXCjNDEV8x0vUX0EDW4Tv0CHI/HEXo6YMtvgudOvDQTfpjg1Li6ztl9nf1l
aB/AAY3niUZ0jHIXTFhEHFbUcnPzJ1qyeUSCmdl98I+jnryg5pAH6A4vjGu6WwgRFEEPA5U6NMWv
mhhbcbX4lCyVFhI6kOgopn+AZamldPu8SZA5KTs9P54el7BepAnri9suJVkgJYTxGugQQZlkplyS
ZztbU1+qrl+dRxtTy3j7slD+rfH/qXDYKi/h6t1mvBsIgUv+2wwm78x3i0UOivP52cwidYZ+DXIG
4iXWZr9UNV68oeVi754rk7Ya9e8+S2LvHvJDKGCNawF8Hk4pXLT3VMpIlN3LhdFjNjjgThE4nI83
PACjm5CZzPpJbmvqLqLc7kZ8jzexAD8mc7X6s7S7zEiOhVxLqAA7wthU1EwOacp91LVUgEGJlbKj
m9UG1WmndT/ZCXXR1xsYoiSDElv4xAd79qY6gSV6ukwfAMFF6Xz8fwN8JVm7kYu7csCN1xTCHJWK
noPPx0LbW7Nw9LKVXDPsWQmUP+OsdkZpdvGKc0fL27BqoAymvZYvH2q0lkh1qxdO+QLqDz0W830j
+tJkqTykt+CXGot88kXkTt/1iuP8JhYdMLgNAU3EmPxkmuBNAsVG8s7huelzXk1a9hcyHLiGudq2
K2UR8XY7DtroME9lkM9zBKalw/kSBwEPfTh6kdWp+rSb2TcDY7NOQsdWVWsZ3qnCB+U87kHdm4wV
DahEWNb7zvJBbXu2AJY+28qxE4T4m12N7bRhJgH0cHKQSKCay/H7iefOHrIyvDEkQhZQYyLnUiqk
6EknZKqX7qbVUdJ9bBuATaB8ugNDlldcDSJXvPKBaPccPBZGMg+ID0XsaUzWBHwr7uVgSDaUuGqK
nwe1YfWOEG68NqtSsehWQAL/T5zeCBTSC1kos1pj5WiHgmyzeDcMXJ1iS0r8RtnT7+K/X4uuGA1L
6lctBX16ECCCPEhiZ8CJC675mpmAr2KPOrKVpooPM8HA2YRhA4l34VB4JC9njVJOke3xHZTkE+Id
VRS/SANTDYsaSQQbNs5a9SdMCRTrf+5Eb6THKo9lUp3T/1jIcnQQunq0ouk+M+QUlaFq4v/xRrHo
ku41dd2+6WE6b2QKTHW4EjV4RkJ7zgB4ohC4yOEGCBe6m3rn9WYjNKiaWP9X219YAZnO5vSUt+Pt
SDZC5H9Lliz6TaTN5TPf3SuHBvQwCJes2kAM1zBexMt6/+KLibOvqGzy88XW2BbRg9za5BAHryGf
vUPhwPtqDaNShiLCLD57AqLQEnx4oFQovTMFazPLySnJvH9dNN/mMx4UUuCVT2quXIoEUHkKw4P+
ZQfYMtOlCPoTRJ3GuFtPKzlm1/pexbeZy0L94OAjhnOpvyMzckNbjUCbZGcsjiW+267KyJiT77aZ
thtJ1ec52O+mi/hAep2vGAd6bqVsrPZGJdJHva5j/w83cWb3eooAQLOkGoL3apY4XaoC3VXrseGN
uikyJjsL3SauAXWXpbSDP2F9xavMtSHXPkHVe+LnrEajvXPJtfkUVjeVD6/GK5pSVSv7OHc1Kd4Y
SFj8xP2uzD/8DfxTVEl49a3Ip+8RySZSsxcA00Ef1UHy2L+RyUAVrMvk5kdqFMf54ZTPxem7Q9UQ
CoCjoDitG8zgd/xs/gRH8jLCgoaXvcAorITEt58gWEAqEL+5UapWS4pxjvj8piI84s4eQwbK0NqW
8evzzfkLkkVYW5Hu6b1g3eE8da/bSe7U9fF3HKriVghu9C0F6+rJ45ZDl882wfO4uBmud3ERdR0f
HhRZQ0mkcspuyhSVF9jEIBUD1+hW/k11TsxR6XrUlFEB4HlnSwCSanM7/qa38IamUNFzVELcQNxN
MpccxLh80bqJMD4KJADl9zLEUa/Ghvsafh8insYuZNxFe28u+E19VqoBeGZJ3lhYNduCPbWIOh7O
I48dKDHlF3++yFimobYTixxvCv/h3REpj0NXP7MrRxKeHEX5yO83SRaHb04M1Bpjv/TA/WRVkvN5
eIXpgaCyKzG6Ygs5eTWEQp2KsxePRnFPnJsnWjdDDaoU96Mx5XVAkQyUEkA+DRvewhWFxsgMFQbM
6U5N7ceTc1jBfeZjN2I+Sz2ISqoKd/oaTIh2asqMMOnOPXtc1jrc6Idfdo1sLy7ZqXIIR1ZLiMVe
m6bKvIoOLLSlnYMRY6hHsM4tBpclispJ0fRe/iDALJdPSRSV5WSRZvSHOL+nrcK8ockHGOjz1vlw
tPKq8kzDANiw4QLJi3HE1c8YPFMtKVY0nq7DzJHaDZhrhRVshmBPipSUcj/e2prvc8lGdI0u9CZ0
nbfaG1SoL8KeiieXcD/BtEC13RZ9ipj87HoRVnRu4K+44YWY4cTkq8YQavZvDVIImD+I4m/JZ19J
4nA/S4FK4JzTVwZiFQKGhHggAFvUnE4AUiCjoiVjvNhD29F+vPkzV7OuNQiDepVKiwO8WWKJuDh+
6HI+aqjsiHNGbjbgdwAD/OEwEY8ETJcrGcZ7ZcU3q7r8gp+RE2ZU9rEu/XLGo+nEH+CQTPJ0ETW7
yG0dz+4pT+XTxPycC7XSsQBLU/u/gu6dRYB982C4AHgxLWw6D7j4G7hQZlPVK1UKi9pXMUK6kTSA
DtWmnIQ0D7rokD85f0BFXwR8uRFzWH3ZbCgLxoRYOTPYSUBDFLFnXzb2lPNmLe39CgeZ1Wmlw1FU
1sHUqNEh0LACqeexI0IlqYqJBhe0r2jz5NzuFVPN4p/t51/MUujn11pL1uBdw+QEJisIX4CqsGsA
SeuI3TMWPOIEf25UqjXuZXL8hyEkUuzF62saLd3uv8RkDOY2PrgFPaX8qI6+yO9gcFObBx0vAGzw
S7JGu+xqTEsF6xDt+klILyQyoupzHk7zN3blQPk+hnNKKygdcYPVKMb3WdpW9WKeIf4u8sO1+r6D
Lp00jW3Puev7HVUOBzlN7ZUggkyqGLujL3AI7KD2iUVHmOj+G2GcVmlBgBYXlO8DF44olPELJkpL
ph5pp+74AL7+hD2Uo4GnXpk8YP+50AFHFzuAtT3xpkPLmGaPLy8y4FKQVyqFwU3T8munZ647OUZ1
VnlfAWikR5VuHjdj0gh8hkYjzIbV7jUlUA+vJIySB5AKi0aiRXTCUyOxlkLjs3aqKmrxV3ZHYyG2
rc1jof3s572PTQ/CwBNoHf9PHa+rHTxhIMgAhZoJJWXHAtaCQR2QB1PcWUBM88KvT6/QaLCtSa5m
U0Yjvca6Top4ysQVdiXoBeXQlF23nzyQQ0kdbbjUYWJP5kzRVit/2tNzOgLSVJ1DCoKZkYC3WJF9
6TjQxkGyA/R9UM+iUNokfMvvC0FtT6DwCsFS3vHT9/76dQnVzb8OjdD7Zxu8Z9du2ullez6TJ91/
6nTynbqNWznUhlfba6xsfQQUwxyOGYgg/vQ/43VPjqm9C//Ef0uJu0Cy/juL736nnTPe+Gh3c6/v
R9JIPiKfG/uPKAQmtKJlj7nVNZ5oNHfWIdZNodvp9wHxuARxigZkaz78A6Ta2resJ7u9eAnp1kpB
ritAPjZjnBJI2ouqZ92YLXwvvQVtdd1YR4aMbPFqO2yUWY+qK2bU9Eb+CBbbjRoRoBaRvszSsOyZ
6hME44jYU1Wdifry8KlZthXMpTb2OszYulAAZbqH2cpt69FwoFo5Gw3oXANnhPodgTZdaG6Q2hQE
FB98yXjqmFfDI8fFNUXT9NgVO2UkvSwvGBnnatucFkJG/PWQoBMiK/0AOiDeZcjIvvtizK0rjQk/
th7EBusymS3jWD6vePZJKwCOerZ3eu7oxsRA/IqNwxJIQ67LlpmJObvA4c/OZmHs/wQVt/dhxOX2
9z16TyRqQnQH7RV6CMUb/ZW1bP+hwjsApq/IMavA/hflxuAp1FvQXeVo/VTilMKAQGn5Z1UGKGTX
hfgLmXgauZdvyAjQKhw6qxAvi3Euq3QW+rIuls/j+ywsHhDXkqa33Wxl9KpMW8SWixi+gMq8Jixn
FeGuHMldPKDYOtksDQPvHmYJcRgI1zSBeZXrOveEU07i6HrcX+J313OFtlkkuWmUMI3Lu7SaLg7F
FTG2/7RltIr0SnpErE8LwFP6CcoS/LY7fW8NU7XbXzgarUiP0ZCb8dHm8vYHG/oGOzuEiipBx7TZ
rabs+kQixYBEcir/CrlJoNI8Cfco/JyA/hNoUb1+1btNZl6oKXXHaDI6LsM26Ik/zQ6mlQl1FGPx
fKllFzLoelTbFdgBj1Bqzp7nUP71Tm8ga99GpmSUYOZjFd3HPbu/F+FqPl6cgMEGwnzNXmf1X/Ax
96AkNoH/p2Cj/dbAHed9Jby7ZDxQZU5IwIBjWRh+EJ3bBNcdDaTeYf9YtCH3KPKIb3zmrpvgSf+y
JE/npBzzKQ3icZSg9hDw/UCja+mCE2O59wq9Y/SelJHs2kpB8pO3io5WhHOm71Pd+RL7nU+6IXOY
KlTwu2RUsOTeSOX08dx+9+aWNs+iXflY9k7JNo/f5kD9gKIeDLQt+s7kNmzSRiqniLljlkC9zO+d
Hsmau84teQn3d7rFAT+6xoaBfEYnMdvplIhDUZCMhkp1xxHxPil17T8HJcSlDTxG+gEFuCRnOXB7
wz+BHcdDbVxyjq9bQECl/kS0po8nCgJrxrGd0/gTgggnqvJL/Z5YlpbUQHb/F4LjgB6SvbM+QXT+
xFEYlMRWHEtv0R8oTiDpHpmCjfFqC4BNdmXLwoHV+SG8/5bBcyZ8NikPrNJXkyIia+ABCLGmh56L
x2wN0M4oYCZCLWzNKPH42y3CMxfSMdoVFnYnbWMeevxMenVqCq+W12sE7Fqv2wdYAOCHzu64Znpp
yi970Hc430R1vU446CsWf1QjKiDOWZCuMUVOuvgy7kJqDe7BGVuXUE9ElW1th9kRIFA1rhmHpXrx
7fqtLRYiAk09FU54LZeRmZpzOjXBVfNDt2SbYEaoNSaaFt9e7hNOIcoLfilrhhCdzRd+bw7o66WD
7ff7v0lPATH0HSUjZ0OPnSYoEGGb7Rj/l8mw0QWw0Ucey41wJQ5EFj7HZD/PIOsLcZ9l5wGbMtfr
JvgvrFUPJxk+lTLRwVIpSrxGqyoD0l5uGx7BsufoQNWH3+Fpp3FDKkw6EBZK66tF9F0RMS11fm/q
TLlQypyD2ch0eVadJ3zsbV2P7cQVIAbtgRV4pwgezSRt8LK6OWbNwc3lXuG7ttC8L2kOr8AZKQ3Q
gCU51qK7f1Pheyz0wBqxi7XR/Mhf0GWS3KSfAa0mZOhwXeyRglq4ehHIuWtUuh5ElD93Ljt6612W
eFh+Onb0XWEIXoZuQyIQiqabZlYC8Vw4VY2AvwCkvSDrnoBlXVJhem/4QZa6qc/gp/JPY4FPMwC7
wvINT72Ng1eIniwWr3384S5gcpCmwsJ2togEfPqR2psAjO/Q/jyQrORg1xLdEnx9YdbNypSwmAqR
5q6g2PV+s6zTjRmu5H/SpcmbwMTbsX0WgSBzzitGPdqnbFZL4B1A+ySYYvh2OLSyu+fGM21ucHQ8
VyZX825ZSwFBo/fWn8/+w6FVb+dDKQ1XbcN7ZkDbn2Ygv40SfMZ4HXOR+BSDCz+XU46w4eVEwP5y
OEkZJRFYhdZT/QoJXAYRmysS2886kJcZ4DsayrzjmbRM9pDrLlDreAy6lNZ/Ytt1dvFgUIroPWJy
gRN8a/3f/UJtUBwOowuGaSa30ptbeeg++UanUprokNkPbOkAC5IIArqCBD9a+U504uTOBziJ8yNh
gcdSnPFXZhsdQWCguR/L0J/hqwem3s9OXdFnlayRPLt7qWW6kq1U0EsHQJdcbiPpHTrJ3sgdPigx
+IJPqeh2BBC9YO+2LCjuznWJRMRzhYG7VH2jwmCY7f8Gl20nFedA/tUTx/cuWSEt9Y5GfGcGnawD
yP7f/N4Y/mGpM4n58cuQG86Kkl6POWQNWLPOMDCgKsVWXAJKuNlT5HQjSTQriiEiLW2A9fkN1hCE
zi8ujNBic55lJjqEf0Y7lNH90bg62kZFElBDZ/xanTxMM/KFO1DpL9fvgBBdk0V2cMmyu1nf9mv+
J2wU4Zy+BIx2g8NZzLtmtYTlJWclXqAG7SDj0KGq0XPXNiEFHGJ0lRiKxCzxjdLV89x+Cq+wnyq8
D6H7cOUTT3nPXQqHWjrKT+gOE8cc8VAfUhcy1gVxkG9yHJ/uNMukybXQiZ7e78WmmE06wx9a1eue
i75izxsGVlP9+fSgKhCjuWoTckK2+2mXpYzic9KHWQjpt+mtkOkXCUtE2o3EDaT001WAF4uTuAU9
//f9bNkbhR4ZX9W5YK+JmoAibnVlYVHDZj0sDRZee5CNCReyOhOiFHEPA/Ggm0UrxlN0y3bODMvT
EVGm1NDReCI8VZ5dYK8MQIctV415JkhdO4clWieWWCQpLaDT3hQ6892x6e2+3t6G8EG81v5FoUfL
SS3E0F+/Os9Y8ioj6ueUtFYwVE687GXTDf+pHy8iQBGI7y9ZF8BX7u2IP2T4x0CiYO02zVZ5uTBA
2ozyWJYk9+kFR8K7MdtcPj+4FTY8p954oV23if49cDiLxZcWX3sXrOC63gbjUR/+0y2JWuJyysWl
qGZ6novRQk85WEIlhPTqvgAvurcghCHjLZot/wW6JYHzkRZberwqyTLf0Z00FN/mZPly5urUkl5u
xxUbPgdJLQtzKsCmMPg1ToR8a1QrSnuTc8n3lhejgJGVbk8rPl4zdEYXYmaTlMGwfFEfEFhMquhr
R/SdCSvWZ/Kagm/XQ3E7wlTPvW2werHg4eUxesetwb+GdnVxQS+ls11ORIdEzh1W17Jc1jnySFgT
c3iMPGqBT8s2ETkzk7EvfnVMEriE43F2YVEOsymG7sfb46FslP3Bl0so/m4o+eymRkxMG/jYxa+y
YweWEEn+dDIhk0U/CRHJznmQ+zUt+kZGt6uwkGKDIsY5vQwDCXk2H3kUe4rlarJxiaXo7hlnWI5u
F5Q9ToakJxbPV+nvkgiBi6c25jQG8zwumds806sckLeNDE/H7yAxdAUDJ0gIa0uBFYGL/oBgyqWR
RDaPQSvKz5BzarxZ8qdzBqUQH42Ip/+dFFLdwXDw4TSDnUwcNOZUZDuBX1lB9gX1r1fK4zXFhGSF
l7jGWyS1c3RjhWZdIW4Okha0SpAJRH0UVkHaA/lYqczAyWKT1i2iMGDy77guHJfrRKBuoQXPYTPM
Ev2pVd/YHg7cKxNV3XFpTygeBNYqaqfzxkrgmO+K5JQhA62ZxTP3VQV1ruYhvHr7tKHRUW6fiieV
NDfWqZAo02El1g1PyOlEczaVvA0/JU9js8LYWx53kTc0Z0NVNGO5TNFOtfVVMkabUsuZuxTT35pg
pI+hgh2gx0Dj0zUPIbMjHvmQX+AE5OCkdYz8oWHjIGbnP9G7CxP2ucgbp8X8QH9tKGWykUuyS7E+
6kBTYMoiuJZcdzQ534V2QwtfsrsWnLxXN/3M0DknVCvExac2p+XhzRKxx5IrDUDR4u3qO+VzalAe
LyTStbYQpFIx4oPpi+kuGh7dHxVpeUuKbt1jgfiwuvyzSHpT/Bd/eoV15QV8XcNV61eF3XOMdCUb
3KTGKJh5TNICCarGBNSaDNc5gJj+PW9+2qQnn/HYt0nS75d1G5NUz5LrDoZf5uZarlL4m/F2F+lK
Z5YP89j76lfv4G0zi1Lu0m6UDtgF7kPc3pgVZnat64Myif9AwFfPr9CFfPO+B6m3wU8fmV2DAQnA
aB2raNKbd/7eSJAOHY0KNjYIqyj2ZrQ8CBMsKd2drKS4JbB2J/LVzm+FVPaHo5e9l2z3kOjB/qO8
0yzfx59d/OnApEyFlC4JxWoe3v+ADMDV+HsuB4di9V/bWxT3hKWfQioEHjVomPI4Cntd0OGm4XKq
SXlIBVJe8m1HQBFYgTaVK1buGmCFnXDlSAj8u8ezipGgizwTZgJZrRqjfjcTFWDLZz4Cp80S9egv
ntWXOeIqonqBg+ioJd0mBibth5o3ouLOXLVnpREsNL0hyNn3rK56vC7qwj1Roh/BkCrGEEkyONc6
/rMxDQI4Kavz+SRhpZSvERX0u7O3vJVzDnKKB+iU7dGYbyXbfABx6EDn6OLl5GYbBhBQzhlUyqNw
6UZ1eh8Sf2ZrEAaf7IUU3y3PKhKTjMdngpNZJHjg2NlzO7YRvgC64F/dfnkTcUehOLD1H0CM7QYl
ttl4GwxjM0/peRdFMTF41JpHjyze1qrKCfWLnA2YhVtioH2rS9hqZl67bDdhoTSo3SwR7wfSPF4b
wSBEFPBFK24rawsAv6aUB4uM9gTjyjFFSTVk1SP84kILx83AyPipXpv3NOlRMHR7/JKFK3CcH8qa
R52humHq3pHXNUvUl6Ne9qmYn/Gh9s6DMevcxx8WBH3L2Q79ELwcVZqKooOLYCcv8p89FvUOH+Bj
aOOE3lXhoQredQdQsMTO7SxMNuWDF4H1l5HnmVXBDkj7LMncqNRgUH6ThRu0zZ4zZ2rS2Gc7SOQJ
0PnWxULPbSTy05YLd29hpdzblFt4/8BEX7S+eqM5DFVXBbyzKvaWi4RNDJf7VmbhdUPHvFuLX52t
U4lbCgd4y9jUdcALbLimBJM2GZUroBi79LAc5VVG/VWY0qXMHvw9r/uiWZgk/EWpikBZQ388JD/t
lOvDv5VYghoqfrfZ9wJEqitTz6FsCAJVTvDx9N7KrKpWnVl7jj7+bfGX8XqRcDHuyFW7Vq6wZyYY
CW19w3nHcui5ljHSxsAM50rHNo1XMxHiziFd0b2w3BLwqPnY9BIVtiCGUVHwUouCcXkMYFoh9inw
B+ywxO7w0rLMfmTMrc74lyzT/xxpjVtSWN9E+51i68ZWO1XLn6V0HJtiIYXQykRFVcBCZtlpt+09
EnG35Aa9YEu+jrIvQCLyh78X48+Uf1iaOMew3bndLep0+XJ+dVTBZN/VMs+YqN/8WoS10k5t/4zh
x//ruJJ8H4YN4/kQ0AWbohelSh4ticdurz6veiQgOrBoBvlhWlyKHYAgd0Md7CcIYQ3UUsJ264Kr
ZlU0v8LoUDKSeRYn/1kERzpVZJ8g8cCmpv620ZGdwEJZbe8Q1pYuoiyj+BG6fP9wAy7fyMCWo80s
0doKn2g6pHvPto0WWAor56TYbzUFSQJsDlzz1LMXvqxqiM9QtRGneYGL7UcaaPiRyJpazEp7c0ew
HG9gwFYaP7tyuYHff2WB2Kauge3zqCVNpYKd2G7p6CiOP4pDMQDl/jCyU7bK4EkESIr2F32bY8fn
whT8L6up9MVCFPCknsHYfr3UPZxY3MZRrluSApnGCLpx1I2qCOeQ+WTWTv+0Bd0ERN9ZimNPJqyW
lvTQKkU/fj6Rl+liua77wd+myauSrbQtECtYQhXM6rfiNarJnfqXeULXh86U+JTfGPGnLFY27EFU
o4LO4GP1dcz1qlhKTrCzuUOmwMQblezH/38KnitRSryWN1H9wh6ayKP2JCkfz1e82n2Jp95v5qns
yraP+V9+r4NRVFJ3lJYT0t8+3EyJ6JEifiLRVYv0JKr2+C7w0No+2+itPNzFsg5ZjQvyGsU4pDIi
XyjDgSLsXqjY0FWRq6U1mKyNT1KxmbJnoyoqM1av9+LpWd8kGrfOOlQsN9kEoyU4NpZ5MiVh6rk0
7RDWTBSidKAPSMQtsHD9tRMCXezLvuSVQJeYGN2z7oiC/84mOHOSQ/tKCV+HTJjl/ge6XhWwFoGc
uBTcIgvCsTvkP+qjO27Fpe804dPTsyCc0xg6VGH4FGJVhsbnr5f+DTNVfwBbvRb14U93sBRcXmRU
rXoWb5a0ITQZrFBsd5EaC0G10HPEFjRgtFkUoFktWdxZd4ytXAyTLxeZLIaFsTP2lnlw+VbFEUtp
FhUfXc7MrAkfLi3B3MK+9eprH4yN+tTm+RQOteyyupPkpeHYN660c0G2C6SabjCKYL9vbfWmSyQo
yIAtqhxlDCGtVkPk4CV5y9orVbiCoJt604OwkjtFPFqm/84aZwFxpZ0eAgjYVd6kNuz47Z0ETULC
nV8d1E+xdEX+dvGwdegZxZYwlzRPYgSFqcv2+fCi7ZMZDcJ/OsfY6izt9iaBjZa0oqv6I7VAjHgI
u2jSaG7cVALDQWd6/OZQFtsOynxF5iKPMoXeLXkd0R1lMx5Cj/a9q/zyrmNefOb4CuYYI3b7HpAG
40uN7qBtATANQfVX5y9gEDGll0G7bpAi1WETG6yvg4vCPTnBOo5S3/CB8EAEk2qcq7ueutVfw6Po
25BuJPRnhBj+ebAc7hO6IeIzSafRwvQTJQZrntvhpZeAaz9a5I/dzoDQF/yNHdOdUxpwKUERIu6w
HbXcocf4F9VumJU/chUzx1xVlbkgkCKUs9UmQc0aG4nwdLTe1P0O6GTO+YDATntEZJYHIj8BVQV1
eDIUjalctwqLzMmKpzC7iLRKMVGUm4qO6OQMsWcFVSdfdiPVHXCz7LDB2lJyQ3BuFMJ3YjpiV85a
K4uMSUid3evaZHIEkurkR9V+pWXcr16p51RvA7lTSmN5I2HYGYeFe0RBh4pMWLLS3UMq0n/1HkjX
yQzU0207AAKugQmLLGYWRV2SUgSj/nGb9+yhsHEEKKefOnwFBDn3SrQMO7jac7kbKe7HRsPxjTnV
NFcaIrSVc+roMpsrG1t/weY1C+HBhB5UQX1d5XgcnTSe73tHf3yJZAPaBzhkTwDO81C72MyJ7YpJ
Kop6AMIYjvKACwKAof0f502lBsHiemPLtgTmC+fNhYZsZ4pK42e8LXw//BrpPEMGRQHJsm09iwii
uKj0fEFKLjth/9vCihRVUcjd/752dlDedcvtS0RV8JZDfexpxr3hdizi8o2X3dqiIILxwivrPC5w
AKNxLyDsFHZtmouyS36LP0VS2RRAvF8iXSzyRdJZv1g4gvLkpEL3jIB7G4rccXcV1HKVD+4bjUy2
15Lm18RLAu+3KSZwYuyeaAl29SMGa9Ll50rds6MZb5q9jtJNjFnbLEaGDhqOxPze9F92AywV8zGT
nYEpHpFROCAgjOQ5PQ1kT5A3czSiB/qU4AH6s0JjoQ3x2kzRI0KQlXhd20KeOtgVHikd9l5uznHb
LoJYV+9KWAaAgf2PI5DIMayFoV483H589F7aUbKjuRw+RjfPY2p55/BfPtT/bcLCSd0GfvWhK5iP
Bs+clyvoJAjrTYDIaKb+8TL4Ikj3fIIcvoZEOZN8AzvRl/I+O3Apf6WQcsdCojoGskKsyYbAire6
1f1azkdu5AQxqr8wixhE1SJ696h7HJy9UJR8N9UrfqTlGFC2vgckq/THfHkBiMWKXgakxqEAtck7
HnC7SWb8QyCjHbIqRd7fZFip84wa3VLfckOBnqtdut3e6IFPemV2j0FsY6lggwojIeqrirUtiyfi
sTO7ThURedIXSPJ+3sPmEE9FcCWkQg1hvsFb82OG4U+HBL3iizdF38bbz+wcXEJELZG1uX2rUD93
xoo0AJ1vUcxe2TXkcZwqe4zAMtg9A7P/pb0bk39ClLgO7dw74n2202EBEo9cqoWh26hd7cabEf4A
9XgmGaZK0V6ohfW963lBPWYiiu0eFj2hzpRN0HJ7p2L3bvgIWvC3YumGZfx71E8MRDYiazbCvUDM
A7AcEFyD79+THIXig3tjsnx54JK2UNmhJzaEOLlDeZRpitqiwCldpjgMvbiG6U7a9GyouwgIzhKF
8F3Xv4+yRMVbdtPbn0RVnPF6jejl2TCdX4+xucVrNtikoWc8QJ0FcDKYF5QrkavpTQ5Cg6BE3FG/
/8NNV++974IJ4ifDkgH3jhT/29kPM+uA6v5KzRZEKNOiLxC9IDKTh4mMt9g3CyZynpyedkmn11cm
5O4TzLnbyeUbKTIqTD3ms93FizR39bOpDo4NmvKcp9TQWAVT8r8vvDfiNDKBjE1CWzesu+bjz/VM
C655Uwna3qi9ehb3WUmxLLFX4HdRVBLUrI1dTNiA4jZVRuMSvJpTO3Mkbnfffrt5E+WOl+t0N1w/
9++T2ug7c1xLAGEFTjpkhjhihdEnpAPRqk0WXUgZKxo2rdCeHcZoZs/9HpUdNr6K21IdL2tKKqfq
paNsY/dNW3o/WehJ+OjyW8n3an60YfhA/agm2++4hwu3iTfgrYQTEAuzSgiRkZ21Koad6kYjY4u7
aRnUtw85eZApRjeSl4hyDT8dUyAtfMBuKcBIBa+h1123ECznkAAOg+zhT6zCPChHqX1OKlhPB9eP
o8ca1tv2nFDL4PWBVUBBdD6DDeJ6dRWgfJe/Zm3RPYIfRIoq/mwLCJz9oVcYXcGf6W3XVN4CbbWB
FiwaNFdSfBeemWp0Gn1CvpXViDmAd7oP4B4xbRIgUnOYRRLoHcVvs8aV0tYWwESVpC/vCkwsL57J
TYVBzQQTHPcQEK1H6tIO0XMuKRjF6xVbKu9ZbhTKbtY1M+1z3QmJEI7qrFEwLjR6FOkKK28VzZ+r
zY29AiFv35ju3F/MT0x+Mu7xsKaYt2BmglXBAnyyTkY2MYH62+jB5CrChDJY9ggwkBeWISnTbBlQ
HhRZGi41TR3UWBz5H47nRNDsuE4TmfPDjT5YbVxZrnkso6fHqfC6x0XSUzQ5iVR2ESbE73nscLQ9
F1R81uDVlrKDwUKTtH0hg+Z8AFkxtPxNwfASewkEAvZt0C96Sm+PFgmY1HnKNxE9oXqKMkhckCJ+
w8rh3JBy8mzxJoP6ThZ/LuIzOCLQdVPTDsJtogg2D0ZE/wqpSNlmf4A17kH3+b61xxDuwCG9XZCI
VnWBvqoI05J67ZOYrlHoS19ejpPNCO8bj0GOnglFPYRFYOQPcuHVcfHl+XkF7LqXByGJxeudm+FE
Cm0HOuIVYBa1xDTjv14LvuvVi0Y2NiJ+bGZ2kiolD8hEXhTr2m2cXBpvvq8yh4O5SLa0nenKNoD7
d9n+GY0e+2PcMCCR2UYOA7S24xRXuRtqtyVqPc4DCIzpECCDR3qLmrwPNFPRzclN+m4a6nu6pC4d
agTGWfTVTQy3c7V0RHizhpUiBpKtCI/obztRUyzqQuCHsV6vDfgr6VsN51XjjQRzG/0iPCnax+Rd
DQuLtr+lnJRxRnByFgqnLSrUBaNRafSajvgzbVe+3ZgO8uiHbRFSGHECR20J8vhVjHpClRx9c3wZ
TKxcpe50dsoAHDhRzgEOR8LFthatXRycdMisDIHNyGjbh8ldLsmwqsZS5Q72QxCFP8rs40TXx/Km
oziAe65KEUJZK6hdScl/0JAtAeJIr+H22l+CYNXbXa1VPoEWdd3BNKo4+yKvCHUQp6lTt+SWCIR5
TW8eB2EzZKtsh+7aqyTGPxKBdmXLw167jGbfCeb3CIuD4tYfE5gTEiuc9rbVAF6BFWxuD/7fEhza
ZbN0oeDimqswko5hk7/kIunYAXYPOqmF8/yRPRyVQHdp8nbh54nIF4lCikFaR1UembBZqbUKy+Hu
Tv9FjimQzryeSn1XNAwDD06ZdajycfRLVQVicL5HI7JOR2aHOeL36vqEaO3aFTTemI9qG2EtlLlq
JC7g9KPmNU6VAMGCIFhnm6DyAFCc9IyrRwAE96iGU0OavepFC3Tqc0FMiL1HBAWg7o2vMkZ7F+YU
/RBR2OgxpO76H7xCwBv/dDnRXsNGib8I5eY0/BxRD2dtNsEfdnOVIoKMZS2Tlxv1nddkGKEELD65
blpiY5l9nJBSaoe2pG5sy0WsH3kQbxUPxKwbl4pvC/zajkPjADrKwXxgsGDQjBM5RILQ0DBy9OqA
qPm4phaf4XGuE30J0bc8Q1wUFFl9g+bpktTcnhIlqhaELP+zuzvYr9TdNZMsX1VCZXutGFC6OoMM
uG3LIf1exRhgvYKssbxML6btwTgq3xWr+EKQar02/ZU63cmS0RIwAfl9qKu/ZDPO1Zat2Fz4QkIf
ruyKOMobxQfBfsIXJaaufGZTq2MDzYjjV86TdVg9ef8r4YVuyFdUNnuQtCH3QdhWCjam3uw0bf7E
DK2vK3mDewhqDF5pC9yTIMK2eJal6G8aH7jcB6VdRu7p8DRQW2/UjHbsw7Bld2smMP0J/+wKwajp
/aQz3dxPeE4MK+6711x4T+i+SQ1X1j5xCis3Jq8UuuNM+Jh/z8lb7lLVazJnzfnPppHlo4Sa6TlW
7jyp8xW5EK0YTKblYdUVNvnfDiZ79h8leVtEQ3BRCss7JOPP7v6l7cEqgUZ6rNHm4RUNeXyo/hGZ
JJ31cMFk+7793KoW8PW7+Ij4qlo2fOy9RhUS3mVgs0RTQj0/JmNXwu61HbLeRcE9qvxbthsiMeTF
utEntoCTVjr+L489m0iE9un5a/MlALKp1uAdgxXZ8ToCOXpLmvxFOXxrevVCGblAa7LY81jxcYO4
v0AA/xHIIrAVTWlfeCRWbaCiYDB67K07cFznKDVODx062cli4LwaTHLPl61Ft4wSKWXpHHLNz070
a8OkOQ/sZ4mF8l9RDMwBxGRMG40sMGgVQCNYHnqI9QweyldzajkGylG30K087Z6oF1tpb1kCEufo
JXLneA9Og+zuQiek/huWkl5NEcrEzxvpOfnqwG8+Ht72OgfDgQkmbK0mJgpNQe3GpUtXFATd95Tg
A6KLgW1w6LNoz+fiNd+dljqyKfMJwONsINktNPAqCyBsuJCX0IHlkrKmPju39no178ynSN7ECxOy
ONXV6mWrhvA5oT+TMhbgVTMNhBNbMfIzu6bkIjYJws8QqaEa+I2LYAJfsoAAawulKhwjtpeMJvhK
9/aMlElrvELcsFX5tx/RV3f9iTCrOK+fdSHH/YZFgBrIBT/EeHjMckcWNmWh7GZ8f3U4w/qFIkEL
yux+FC0iauhjUFpsX3/Oh+oFqygYMV3ZuGD8WLsA47REqpwxCa01aadb1i0kFaG3K9kJEnyBUyLr
Hbf1LyWC2T65VlVwafACcouY7WxKK7UoF7VQ9FKddVmo0sbeqirWUKj+KyVhF7R/NAlPq/wDQ56u
KiVayOzH7Ct2BTi/3XgRPebTvFSTeHdjkxkbnyveRk1lbQNa4o8fzTZM8b7QGKgWBXRE0FbZL4pt
0fu4QRU8TnkrInMhNLxuEgztmkiwACoxveDvkpRcwBxjl+LuBH5Qt2bo9PBmbFiqN4zVtR59TZaq
/uzV/ePd33MhHhfYm2uDDhksE2klnQE8Jsylw4phpQEqaFqKGUqcSIzPnRX1TTHpmqwMMUpWJTny
GbdvpyLAoyvlO45JPn8F2v89fszbRhF75eG4JAjNbKhLh8wP8kokSzKwsXadKQgYCFrVxcpu+Quf
LJBRR8A//qHAmIAb3BTThpqaBjFfFohr8IU8GMZ+s6q0n1YcFn0gFo/bkIt+irehOIwKdXzpGMhI
dbG5xBzH7QJXAguiU7MZUEzl4XmCG2tvhbeANHIjjPowF4D5ExUknPGw1sbgef1gzHmurQ1x/F1L
nuEdbEGobkAUOF+jGhHePElTOXzBokLZxBJrdjeTxDbj5oVLbcgkuW0CAjTMIdG+XBjKRzscv5Tx
BPvfJKYduyHNRPjAIRYBXS2Ln5gLZC1nGaY7o1Xl7tzRhFmy0dwS6HEjMeos1Hhnh2PaS+mJprYg
E+2jZpDyOou2Yy6bQJ2o+FPT+/VzOjzXAwZ1a0lwhKo+zKUiE+r/gL+2XJA0CXM7TtJSIzmVME6d
ZG+bGeZpv5Oe30kbN7wJvWFx0fAJdaPd8eVaBXvo1jFvJU7tQ/HR2LH4OpM95Ns+y80UvcI0u9KR
t93+O5ZFm6pg1xRmf/niVb4GuFwCCR/it3wwUxu2V/rRG4D2UwaxY0rNzc7MPNkiQMvHBvrC0+wL
fuupDL60JvubL1Lu5qHq48bE5DK7fzz/A31QNKHvL6SNu1072TWthm8Iiu8MS6zPx3dmajOtXNkn
zwmIY5hKLQNmA8fGfL6XRRyfxX08a87HdAhDyHk60C5AokQP9wtjB81tBJlaxfwZddtXPcZCP2zP
BLaXKnLv++XZCA4TU7PNeWGFHdYmBNfSqhVcDlWj7IeRjG/+yRD9Oc4udlTVA+GiNl0hZkDI9VAT
CWswirMpPnUjl4AaIKKvKPotPnNvnZU4B9JXRCvjymyMJ+FEgIhwXfjhq+O6aXTu1sOm4XX8vKn7
Rdw+Vw9+JZfofaFiBSbjPTLbZ0yKo9Q9S9QZX5Ae6JLdOiXBuTIFR/AU87AooexcvZ5H1xdz72Ok
btF+xG8qLMf3RSd5tvwiOMpTO5f6d1AsuckOiRqS1i8wA6LuhYs5NYys/DLZ2j1tIimIFfPsbnYC
o/CVwGO4yFvOrqUNuUomRQx2JWmLEp3yFLJUjvONLAKYapyP5fEa/mDcpiN1CD4Xi8XgxnxTQzoB
nj/V9jcVYQuFTpFf1Y782fHR1LmRFIl8zNuorqbbdSIxRrA7aGRIvW7a+Qw1J8nnijSfmvCEZhFD
kzqt3beQLsGQpqzRx/8MCj3e1GPh23udfd3M0wOZT0Fj2Srw21xTDUdgOjJ5ZGOBQjoVu4ono72h
Ff5KXD4vganFYRe397s0EchSaf+kDVvBI11sSut38mhZfFVGcrqvK8Q0nLpNph9EoMEDpwKGXKan
oTlcs7Y8lF5z5NoW/Ki0+XRuYbY4vEl6EMmFR6P+ptmF5xGVln5pAO+k+6Ofp4smtEIThW1gacN+
OE2M62MN9L1+oGceNNrNkVlzrJw9vTt53G2L6dPQGY0J2VIvNira0w47sje+jwuyDjLV5oWA5739
yAwrZlCG6GwmjMDVpChCf/77oUHDVeAjXHzmvmXwL8WIQpaGUp299Hai6EHkJkDlUy8Pt3hfX1be
9cJEbSMdLTD8PkaYKIQnS3KmR72b7SB/3EDiSupLBX2JWDyBgktN+9WQw2rJJbPiYgheIKG1gbpH
kt01N8WKQGtuzT7JVyGr9OXjSfZe3+LdQjyU3gJBeO7tjE7Yg/t7lHuYEBAvww/QtnLF0HwXpylL
HxtEKIpwoxIDPfFZkdcfDtJrETb3KLOhwxIgk+mkJ4QwtJLuVdIQDbjo52LSbG62HplMhclkb3ij
DZ9zj3gv/E76NSFF/riuCOrsrCwYztU1Ho6eodkfmdzHD436kpQr5uZM3xbmkKb/yIoaT3+z9RaT
D5jahVtSPs4VehUavzqLeBg1dhOMpIwXmPCmrm5YGn1EUq4i6ifruORpcVX03PYYS08BSXqh03qS
Vtdekz7zv/uXyu4afzbSHgpNY71NJ5l5ZOKibskyEm+4oQJlphn/2cIl+61PJ6gldcenIzP9pSED
+5YIK71XHSyj/IlMHYYgRDUilBZT7GyAVTEBTv29MoqHY44UVzErzm9jVLcjbu2Ru1lcgoZJo1d+
wNx1GpTHIvazTHEyoQrnnDQXXoHiZSk0yLWa7LSAwg0xPt8FdCzudNPTiCz9WkFbUIsMxekddBUf
5X4k6P0H+qUwcMW3c0umY0/suhInsnBhC5KI+P71X6W+SZ9ihx7MuLb+hVbsEC05PNcE73a7Fvzj
j6BHoznHwCoE/OaCUIsXXwIe5QC6GsYr8PX+zcjZE2Zjq0ogOB6DYeec1LKfxPbVc8calU7iDuX7
hgd/B9f4JuPjYtU+Sr7KSjUtjAU3vzqGICF5HWOV9HG45C/F0X/BizmLwkqt+muLOahgagREM6cC
1ygSPHL51NrYshnuoAOFXKmQqKSTQm8vMNnTfZQDYtBblwnfz4k4UaOLDOxcFjh7/tYXnuPlAY/m
pDEsW0NZz+VKBOqkp9owIzMr24De21VJd6hwgcWBwEdICH6RlaUjzjo3pqD38DUYhQa5OD+sGkkl
KS0FG1i1w1LGMh3+5D5Hu0y2cZfZk/FuTpfTs8p0WjUim/4PDWvjTnUyB2xrGXRbQIWkEMSWOE69
/wnP9Dojqdc5xOIst8X96sKH11nV/aFEASHunIxorPG9haMfgv7LeunHVY4f2uu/Bg4kHczBfALD
413+r5hhPbmpE+GTk//KNqoBBwZCfOVk9GZFn23KRoiGKXjEB44Q8q1hi8f6felysWqWpEl5pCYP
ocLZYH8WfCQ2Jw9LjwAgkh/aF40KpDYM4LXQdJObMdF8i0bOmuIn9GHf4DFZyqsbz3qEad7v0vaF
K/JxB1ZFsZxeoiwACnwYw2CTJKV7fsSmKJ8sSgLS/OYGYX+aKnFsrS8L/sh2e6w09sjqSzrGfuci
nw4U0b+4v/bOk+RP/H+oyxjvqdT2/iwS0Eb4cANihbARYUCbT4wQaBrQ5hsw5SeIdMAcwuDCkH+k
ECWuD3zvs6Sr3ode9q8zYFvFYfgtH+Rjf7XIHPJeOwo5cjypns8JTTpIfCUOmkEIi74Cii8663pP
uJLwh52a/3PdiFKIHCwtrhOA9gK9+HhwGswUxnBcE1KeZkwAGw8ngCzDb/DddKA7ejlMe2Y6Fk7a
EsMAI0xT7z6/F+7qwJ2Zc0ydm77LixnDyacmLAvUeM6AGrbL2AWUixkIl7sttT98nh5XqFukXyjC
WVTmDuu6wqgAJovesUVJfLMn+LAQKiOVj8CJALVJWvQ820fJqcY4CpQO28SwrdhTgaqvTpQ1crSo
7Ud97NjggH1Axnvj/6wj9guaP8034bblqD13p2jwNvHUvpb2wVOPYkXWecziTigu+1c/cpVGyZlY
LON5HApkJOacdUVNRu2H8oYcIO5J4OcPsLu4SQQOU8wmI3NbYy5sAUfKHbTSbG1YYp/+fC0UvcVX
/dOU3NobWljg/T3uTCnaL3C7taT8/mMFmDU9y/FeN14H+UTgdDOV1HzEdJeu3A/GIB1MrEt5sGcX
sAQJRQTEPVXUZjRctbjIj+Ru+kj7GpOXq76QYL3ItBgXVhMv5TLDvX4YTbe8339OyhBjrMzyPO7F
5ZiICryQmEBhGzekXEv6s21w9PnOpSTkjdCWbXMy0mGLwcBbkurUVXa3Vi6Q1oGWzLYMSmRNc8/F
osk94OiaR4eKmVZZerafNYpRfq757W/GJ4WlVqt3/G8+Kvc0UwU1hKf8NwYT6UZW+59eiLQTNr0T
kef4pWiKaS/htziyM8jCDvTewOS2xRW703crxh597vjzomtRkSaFU418u52W5j+mnIcJEcMJAH0I
CHQq+u5akXAmAIt1JKF8oBkRvD8Hc11NujTGsMqZgPiQZH8W9EG1U8yrdxL4Zpos3wKXISqpXQd4
WCdXFVKCwHouSVjsl0nABt/L+TsevMgqQXy+n6aEQGiDpHRUVtxWaXGbmvW9Y/8o5TkYYJKUYvJF
sZ2WdKMjwAYxFHsd+X11L0dc5qOTNZeGfviITP69pY0C28ql1SxjMWxALT067FewIdhe/pzjKol1
cRQjuiSENHqZShHA1096hXD21sa8rvml8bOr04QZhGMiJDt9QV6tonUcFaX8GjwJrC38VuTTmHwR
B5FqWw6NKD5by6nYSYQSqjgGNybZMD/N0sAm9qDYEi2Wte7Hz4K8Ja92oDGtpE9c8J68BlniLCzl
wF09yFgppIwOLAhOvfsTY869WfrCsjN1Bhh6OO5s4rey7uIA0w5Ebn/+A/RsJFSYnZXV2XLrikf1
lwpsyvOH0CFxj31+yBCoWe3RVUl7z6hTHHntDF9zrTFRQJQ6MXSgD5U8dnylcGcL1WqCs3KTs8UY
6p9EZJhPyab5z5Qvs5QAzcf2XDhvNNu+Ob4FlrLhvOa7+3rEa1aV7ixx8eT8mhcAQeGFq0HT6LSY
fXVir5FDqbyQXUP6WDCwoKjwxLbRbfqR4aBbcg2BSrJiK/4r3RcqJWkuZarquXMA10wgsCw6R1YY
ghitxScJZrSlZ5QlTXMBNM6l/pzo9Y5Q8BYG+MSZh865HCXXjC0S/uEpmkQsdflJYiJvjCQi8qmn
KeBXsrpKDA3IwHHPVt+gDTaTY1RbteKkH3ZqLUubHzbUrdbTjGuxfvwpNClOp231L8N6pkhj46G1
hOfUU/4OHS+8EL2xCG063ps1g5n3e06XHGg8Fgzn/8zR8V82B0SQnBCziLq/ukKlllV6B413mpGY
WfekEXNfO8mz2m6VAc54reZS40SqR7fh3MGG0/WHdRRLiPPIYccYFiNHTnkS3pI+I0bY2IDo4FpC
ROJ3HfOy9/08g9FNbeUFvjugTkSBqoYrhneKxyFdAy9iWA2MI4SbPphn6n1ei2X9lMo2qeoFM4m4
jvUg+azr8MuYk8WYhlsPO7Ihuzo9/jLiWQf0nWq4+LWtYR3jNtpYx/Qqa1GkocAMybiiXF6/B5t3
8t4/jBUWR2Uq5hK9oH9uuPAn3Ofnkvw92Q6Rvt6evYS2pWy+5Eo1MfyF156aStSBnlRQEhyTP3NQ
2Srlu49YB19PP/EtxEDFZapXklWssarZxbJe5r0R/fBmdCiJeLzgkADoMuF+oYl8KDopcMlVxmF5
mN2Knx+EBCSRig3JYsfFNMCWiIrBaM9YbYbMQ0qKUMbbckH43n8DflsquR8oc7gS1SqoQk9+uFcy
X6J7b40wvuByJ65mffly0wufU0Ei3qVEvTcYDiEFhWK52bfw6W7w+imsUl6QSpQX7nUQJssFms1m
RbzdqqPaVPeHE3PU3Cl3G2rfuhhmyBFa8Pcf+JRARNSEGQbeCN1u0+OGxNqUioQL6kXczRvF6VAP
EPkMtHi16wwjYQrrytdZyqXzHPSoSB1ia6nOtXXGBxGpei1I1VtQ1aJQvy9D7/xyqEhIWKMaP1ek
UaxEhYSegy6DcUPzVCvhaoVn2QD/lwUj4FdQEQUJgM6el1VPoyo64qmC1NX/6Pbhc+j7QHQFx2r7
dLzKPgQbgO0t7zYftN6Gq+kVvTcidhl/KtTWzdokGGK0/zzUwHLAVmu+BNKmf3PD+MCKD0V65iAg
k34aQRvv3xfrbdl1JilY0epvbLmXvJ6HB9UhPomBJ+hEvshx9umN61RkRZvO2Uvz4mF8BlS1UYeH
3J0EwD6iB+EqUKG6VdRNp5zAbjpKRaqJwU89yj8HQtln1r0BrO2DMvV5NEwbjMC9bRM64rkPEw6v
e0lUKUlrWSHBupAiHXLrioP253nbkuNUrVBainUaYsniaegj37ba25JKyQVPVuXsXbQY97XTqRjG
1bXdKe0DF6YCLuafmxONhuPk5XkYlvg9De/WDi2GYfoZBTEWO+OFRv5CCJLRC60Y6ZTjK3eeddIt
3Hh9IUcpsz0JsfhI4XwAUD6wcqHJZyqNyF+T/AE6mxBbAh/8Z6BhnPo6S4X2NSIsJWLVOzjHbnyb
+qcHzAeJvm5+6oYjhhYgwri45/I6k0d7eEPFgok5gaigPn0YpSfFidubMNF7BEIvD+7OlAZpoB7i
dDNC3kVnsRT8GRM5afujQW6GluMp85RFWd4rvvtaJNz6zNq6THiu8JOLSFEnQPNqZLiJZfyf27sY
xiRST1g2nJnPS/hzImKjzNVbbMJ9d01GBAO5AVf9m92NVvp30H8tu3t/8hpDNjndVQwRfuglAeQb
6f3daUOBzuQIYjIwLJVBUQYQ+H/NO++uidL3kiCKh/afZCtcgmNsAYmRrMQm62TvBOl/O1czNBzj
jii8CpDvWwzXqolV548Eigta3DQM9/ff+3fba3Z0Z2fPkCvx5csVmP39C3+Wlt8UvZSPyL3D9jQn
SWh7bh9Z41l1NKkppx8DnwLDlg8qtsvpb0NdDRpzf0aixdZuPoi8rccbTQ9Y8icLRE04HUu2y9a2
QqFeXduxV/oZ6iXQYcPBzvXqP52hppq2MYcvtS4CvGmHRFwC9dC1oPNKCSaT27iPTeY4V3Jtga0n
H0qLHhJOab8xmTrnfQDCtUz43DAVky+pPBZzEg3RgV9+bzVxY2nBDAi1x8OWxnCDHPUsd87GdrT3
1oirKT0a526UOmYDXA4UXZpogLl6v16cvq5UWTk2BWIbZM+3kKzsMysd8DGjeZVAz0Or5UDOcr2L
LUMpr7t4ewKDQPRkk/beKGSpabpNLInGBqagfQ2D9T1wiF4Yc9bYm6idSmKHfK1w64AxMeyxVsPy
qI/kZjyShgjvgwQwlIUWh1vi6o5XVXDC44VfjMUz7M6ACG1O6h2m4GS8WCFJyCiNmwISf9fan+NJ
giRuPW9sNiuUP8M/Vr4Uj+voudxnNLiVlSooCfjAmXFauvbO19eYizsHagtoP9yxyKyH+NRGKIeY
2UXg21NtgJcTzi24dwDa4/jErr3kL6TawT4ZagHkR9Xx9IbOwLe9+BUeP6LtMz9OgNJfJxh9XgIw
Oe0pRv3FtkBaRUF+NhnD7ef8cpHtBmbvItig1rHZUHKcaUrNPcVAEbmOqh/10m5c4y/mjq0gPQzY
vivJPRDhAHQUcwJVB3aJmCboR4I1c08a0PUaPl/kutql2ThLgLMjUozJvPU53zWkFoQDHV8dIwxr
kGG+0eccqJDwiXM3T8IvpCsJjrEKdM+8CXHS9hBWWACqhsla3F5ojriLYJOGls58S+Uu3t57+b5t
zHnwQvjebxYuwYIbdjBO/RUZ7Af30alWJ0WueqgqddFfnL8j2gMmmNQoCWURm4HktTClglqAhVcn
slHkjtANUo6EJSltsCWHSF2z5qv/222664Z05NGJhw4x1inUJWzjzIb5dq8lEp+B0v8mjkmHMy18
Q6+86IOkJ7PTAWEybG61H98+O/HGlna+0KRQ5z841LphqjchIQ95QzW7xsybtpdUOoJiLcN3u0nt
KNxAgC2xtscEnXntH63CWhFWM4jF9wvpO8dTH8lv3f9WAXEoSnc1gh/V4IFhHwA6WF/4xFL0lONB
cDQrJbwPc6YpxmZ03+1tXj0b59LX2yxwn78RhHAzOptA2CzmJYDYsx0/knFN3DjBS0nd6qD231F7
9pd73k3Oy0H9MOfjsj9pysJKOGZcc6DgtZoByEdfOPgDfPwXzySGZis4y/6tzKCWNBvepp6n7WIU
+QbVjPoGdwHIh4uHwDd0z8wI9POSb4wa8MUTf95bJsaxuYIppsExZJV96x2ZUy0rmTKdx8F4AmXG
HuO4Pqjq9E8LQ4pr9yqqnUMellwpLFsuk/tIQkOZp3MPdSLeQ7hd15TU3h4mVjhjni/7YrFJR6Sr
jMrL5JxzhNy+xSpD4fW64HUht0ysAhABOkT9DjuFnx5dPSZvg/PmK2/GzAfARjPt59UBPT8yoXuH
dXFenBdhzLGOu/tsWzJq3dIQc/ozIp/Hm3XghND8sXAqYcxYCa+os5PR+mFBv4eH1TAXoe2ryswr
qCU9mZZraaTiEXOd/+obyyPnPcekck6+bgD9V6eJ6BB4EGKBsUWm6JEPA+3Ekw4Bv29lMIChLa1S
cyX1QQQjsA9icDzMw8zSjKt5Ty6os/bghVW5PkTeLmJrH1+ZtKQK7gFFcjD/Vye4aFZaJOWB0RmB
Nu7cz9/xRyhAlOtSX/okRAs36qPTOjalK1RG/9ut4ohOimqHRVqprw5/yUzVTInLXFxCn9PCWfjV
sYtFJ6snQQeJbEWzS3ollsEgpGPhM90gkKOtKfIsJMXOTwvTpWlBkComC232d9jq5nPsu9SsW57T
fWLAxG9lBW0KXHUZ+MVES5BjqoO8ViG7hMkj0kzaaAa1RA6A+10p+2z2gEqYv8J4PL+b7c46zDs2
DUyok8l82VYymazmWc2gcTuE6TvtdwILJjXf4hPSeZvj+c83YGaKdfxRFeymStzhjif80E1Lhzlu
41WQSnzO2UwjuORfGBPNkWIxa55J3hHM5Lg5uUTKoeSOLcUrxFTgTINoykDjjRE9SxxaYSqS7lcO
TYDPPcu9wfKoWg45SfEiFD9GGXYTVWwM+aaJEqUcrwOKQFVsJD49+k8krm5+6iaCJizfsF6BrAcW
DzzwrEEN8NQ5nr2mUuXyaygt6ZLuccwMrghqsk6EGHw3uevjctYp4qIFQ/EYtRlxWpcad2NUXSWr
2Y91QWfw0hUj9g0J9TYe0i34NhqYQXfGIkDeauE0aB7IOkUiwnTE4pWuYlfxLoplG/sZLt21z3jR
c4fsWya/2MeFsXlmZwn7Hw7iToOoHOsgzwhjvt3op0C3EsGkyl+Zirtn3kNYjL+e4nHvCphn0Xlj
e6Nik53Pm/95mjidbnUhNsoNUXpO+MiNkpAUCd9FaLGr14wsaEJErhDCQQrmB49h7mQvwKHfC5xn
1hBHNPgc3GNXjeDv8srT1wU0gGHsCaPgU7A5x9V8Z0ApAeHtoG2RiQYkG2aSh51dr4y5/EDAXOFU
TB76fQHa976dNHXlPbkAH8KkSMglJur+5sjwPqrDwOAccTA3KOAichoUC/aCrHU27QBhJVSIDyQE
5zPpQIy/SEd0/CaYTMzmDTL/NOOoG6INM0OczBwIk8JkwGuFWa5McwbLMvBfqcIpCVxWIJvOVmbG
LHAPjEWWK1N04El6THLJ1chsFxPenWf8qazPM4/AQxg4QI2CoNmjT7MyNbVWLF/zHyb/oCPjvAvf
f0BP5RALPKnjYyS5SOTJf8YphC0+WwZpoaDyQseCpQi6XK9+OA9Plt2TGNXWUM+ulelWEaM53oat
WrlktcH9mtWMkku4Q62Fy/7EdJtBdyX0d1MBc/yO7qgMqzhoyQAKQjEk8rn/QEOfqosEy+MuUURQ
ThOnaKKtM93GikCYqXOkozpdhMqc99HPGUQYNHaLB1XAktMgj2fZCBBNlZ0PZnhge3bxeoO2FOBY
G4qHupkgRo7Qj8Sh6vP76dk3E5gX99DGo6iO2aOGOFGVHwL1kmq58k0mOSZDcOcFbR2gKLlmxqUQ
+QFDLI+ek9fSRSp0WTMRovypxvJEcHWxOzAOQvqtdyyTCSl5eBBmKzW+3eGmD5cKWwNvvjBRwifb
AZ5EdFJYusn2I0clXL/7pgYRUtGB21SneQAnOXh0hH+H04KshWCFThwAsnCV9C3A0V1pqJf4Ok7v
7Y8VN6xUNbGIoScJSpONLStX1WufWsQtvIRuekHdtUkeD6gw2YBqiMiAQzhzxuc0c/4co3PwBQwu
Ssj+04k84wkb2eB0lMdfHk22LJn1pnWTqrTYL08D16W0p+swo9fCav7IaOqQdycTtgcspwxkvHCQ
Ibpv01u/XuH0vXGr2UDoLh/gyI9440xHHn8vLYniBgFvPAMOMYHGqx1kIaoQerc5GkLJbUNcLtgL
r32ve60RPvmGGVkCf33JycGD22I+41RozozSmkPT8FGHc+YRH+tWbxmlK8eKsiwB9MIrrXUAKzYi
twqdoEvj5V37pJPiK7RQWTHsyZF7Ilck/8ozEaa2YiK7n3qyiOWzTMMh7XG5XbubQzzMIqfMEDC8
8ZxACSR6HuRBfzrsDvQG9iFPsK95XkPaqSWCagytpn9S+DMY4Pnv0gXssy+ClJXj3NCPXq2lMAQS
4JoO8Ue7LLuhe6ch7Sx6AsQKI3pF4Jx9kAv3ymoaM8KxgQ/sQCPD7kutPC77bKmVzRqvuZ7x10Ps
W2Re8xSkCGyvj0tjxgz17W76ud19YXU9qtgs3c6YyXblOkDJ3aZpREdzJV3rtZVovkJYjW0/rRwn
JtWGlAvYTsgX6I+DvhCwq4lHHAOdUm4h2RP6ITejLXhxnzHS2shqz7A/i/kVXNOAOL7eD2m2qApc
PqxPWxcxgTdV0n52Y7XRGmEQcINDwynLpds1RiSoGK1YXwyvePd3toOIeLAoxDk1XPwABTYIGCom
bFUcw+SvQdHhhNx2yZjB/P3HI+eKZSvRFuLnyiM9mtva7nKUX1UCyFRjsYwT2nKPcD6dnkoqHdAA
unP9v6MBNCTf5hBbhnSavAqt4Gtr0OCSLWSJ06aeAIYf5JujSe5K4SVpYZrzEUxal+qjwpPVhGKB
jFW3fSMZ5z7ksOrxmFVXuJvRLEqp2TdAo+9w/WsJSnFkQFPaB/rNPia9XPPPup7wyAsFgGN/Bl1p
v1MwzARMjUdX/hgTOqCUX7m8fBKdeY+PyOoaAa4ekaoNKQYKzdWr6s+jcOQMFmtNv+q+x4ikPFga
8fzIrb3Ck04vQqa7npGNfx74I2bq9zb/HSqQIQt7IWJV1cxnqk7AD4cOSg6XpP1Zt3r7RzKLlu6o
YAQgxBsn0CLOjc4WopYx+UvAg0gUvviQu+7sETMzWXHXdgTcDAhtzI2+9KXsSj0C4JyM8/T8mKnm
XghYtahzmopB5EtXw63p3a4WxZ0V3Lyzp6ISvLXU0kvk/O2nq4+3tJ+IvGdEkmFMc64l9DigLbDb
ijXw568A8Up1zjGIMqHgRcRxMON5jFuyI+u8udfLccDNNwMmc/kl0vkxZJX30Ca0RhqNyQNRCIng
ITk5Le/dbK08zJEl8UFdBJKewRoEWWT9uhjU/309aN9EUiqLjfObzhfc/iofrq0bUrzf8qbO85wc
X5wGNzwFiX5gkBc1BHHHg+DPu1swEw/0VGzZsIR4W09qlqfu6yvI+gb1e4vaesnJzWoJ4/Gi6B+V
M8Ek2FWZysHS7JGUkguSL7CuhdQMiGAgdd2v5t/3vOwvYdYri0TuUZc46StIlBUMxwgR0VMzthtx
yQtEUdBFg7HGB9p4TAY5VdS5rj5QrSvsssq0+Bn8AmegsUxjPkeWKs1LdqYsKeEMqtlvNIZMWV4X
E3gLiFvGXvWUySH51GHzDJwoXIyZCWXqd3TfjcNdbFW4gj0e+yAXInCxJrJU7LWUj5+e3raWhnen
QNHsia82RKGmH9YTB4UHadb1FYXfpvvHbelHaDbeKr7giNxO3UzoFVzND754P6p/H44wzM8N3YjL
B0HqglCmvxMzbOgTlpLOJMb3+nLQgP90GmqPZ28ZUy2DPYPnd8bkE8h7L95X68WrlAAybs4SceYZ
n816z2AoPXVKHgceE6sFJ60XW4nGIEuQiLbg0PzUMcq0CW98mh5jdmBQ0PhCYOYtIvJvrVukXQmq
HveTYJbtvgiOqkFMftzEci/1RXhj9hK7REE/OcyVqDXaE916MUjF+hChVA7YoLyFgqxGRlKMd682
asnkV8aANh3HGB8jxo35DrgGYhhW3oQFf9W5ptPh5CQWSzERvRQ8r9MuvDyz2oC3+7HJ/4a4Guji
XCps/dAzcY6DUWVLtG/lYm3CZhGShCNadeCddU6gkowjI9zSZUUYexkZw1GioaCOWFAE1fDva27f
lvqYOG0UEEp+ChnRMHJxXzuwH/gCwTywE8hmE47geSUS2yC8YxHF/tccEl1y9r/wy3IFAuql6Fzh
UvYcG5cSsWZCSXzAHCM1zkl0r32c5VNuxntNY5g7cUbEgSvUVdybOpuQ08FZNOi93qtTswIjawRW
NrutEM5s7lvDr6YNwc/a4ILvX6TWq49r2Kz9Je2xo8EjK5hQKqKrVGcQCmUOAoWeBCIY22dk0Bmm
oxVJP81u2kfZeS4XoG07cZhTE/X5FoGd/8gX+bK5K045zNyFW/BnwogOaUqDH0c+zuJ3NHJZ8yx7
zAoICfNCfriddMQWijl1fTpqUwbqvS8+uQ8apujwkIBjbFTgVma+WjVwaMZhc9ecxk57jq27VsZ7
+/l7BfF/RJgXZJQ7ZYIzEFdql0zZhSe/4FHFwO+HaKA4oV3jdhj42HaSLPZhStSzPYxQ+08LvyIq
nuTYK3Igt5rGgYjuzHlu4EH0szycocDyIKtXPYpMxg0InY8h8OmDCamsYS8IRK0rcscRsXqvO5IG
kKnkX9+IuYDqVVr/3R3tRB4L3nm512fUMXr/4pWU/tnyszVWeWoXA5sgd6XssclwVLi1fG+zJo+p
Q1W3BwUaDovPV9D9oUt6ZQnVlykMznoiunIr3ZqbGKaBU6zddNxp++jL+y/7WZa3ag+tkGVRA0Tb
C+SOrVMmWBgt1p4y/9+lRAX3sbF9n6OEDDt/33JpF/1Z95op34AzUpIzTl+01Uf02VKKbV9QG7kd
l5vsUO7JFQNwLrlO7OelX2V+p4uet4PXgNPQ4k+KzFTnDz102lxSFye+GTonkLK6O+kcX+sqo5LE
NJ+rcRVYGvhbEMS0GTpzX6oJv+CwjwhiKAK0riOqbbzbdeoirmfKcgdTMExBWveF8dcWNsvzbMCk
21hTjAxOcWK7BLTOF7ApCH6CGN4+0AryLZomh/gWuEpj+3ZFaMSKbyWbQvvkHnVxsM8f4LkU0d3H
5ZrNmDNELHfVshIi0vz1et20Aq/8bs5zSbkNjVxEncoFvNB0yXUPRSL0KrT/k9eBXGd+XiXoByKi
w1gMQvA9+bW3JB5L/5SgwtHNWEJxy2m/krUbRiwgesN/5AG/Rgt+/jav2orIE5L6xTSwMM07w3Dc
Y8GvhS1rm6gD13XOkH0b080l21PVojebCWLwYYjg3a9FDEhtEO8mhIhEcSKvYny0sGkCATEITxnj
1uGu77Ep1f+x8oaRYJOY6e0tYrB7W0YsTgTOFmzwcsDS1tNhy32/S57E+Sev3+kCjiIAfjVmUmzo
P9ojsc0ECJtf7/9oHgQs6hk0sh/8r7cioAv6H9M8AgmaAwIIbXS1JY3XJ0vR18oyfEGhHIN8A+zk
sN+Ty07VBCtDKYKNkhpYzPJCaBdhkXkC1dbM4Cm5/dgY1dfSzrUjgVHGznT7KPyTEWPmp8kAZL3T
+3AHfbAdIiHIe6XCQ5yz54uhf4qcUOK0lub92ryQEDZ7SsUZGeW4b2QNtbve6bYNvw6bbNbZ0wgx
/s90UBg6Ac+LRCKWTVPL+/Hh5D2OObbCdcFliOOpcMz/syKyCqaeEsYlBiooZBNxGvvPzyjOfkGq
siuL24PzKRhPWCXUH/9fzntJxgIQxM9miIINdthSoHQpdXh85uLT7Mm0zPYuynA8dZAebrP0AJ5g
JfZl1Xdhl9AYZSe8SlW3EKWCehBhFfkqEJfY3tQcTsK1L6ScByN9VahWQMfuG33ADVa5tbiIGxtu
1TNSc93CSYXX76sbnYI1gR4lsubBBK/medWo1c7z0nbveL4WigkjJYI6l9oABxQXBfEUYfz6nDIW
uZ/hqm0PexzQJN3oV8ly8S0TAcLxGZI9wS4xeIPMaDGV0w0LNxzvg8scd69Y7aEAcyLi00EwhS8Z
qixT8Te7F07s4NVOJ5bxsAy39Ifzo4J+IfkNv1d3i/SWVawnCVSIat+xgkERepZwwb51+0PJckpi
+x9CHPKc6XhZWNsfiIJ78AxtzJZjR6rrP4I0IzGwIZF5ES6RW4WUOKHwh+Jh0lMhmuwQNuR27tvR
jkXoFrdB6qqEWukigvpuv6F5XIGAZQFwVzq974VtAtnRbPk5vVUFMLP45hvh4jkRJnnNxnMQz3iW
ySbjgsXa0d6DTacmHV/k6jbRfnltj/Angb/joA4/38Br5ZaEgGAYvLNegzPa905Q+KLHTwbtHzwF
bO5kSuSwPHshT/HHsvgSYqA5K1ED0/43rHcyY9WjdrM/ElYpuqAh3G0VxmztFlBFqW5KSDiGhijO
IxdPAYr6yiH3gEoFwi/YMA8hrL5aO1ViAb46Zl4mvQCtzKHweIkqqwH8hZ4wq/YP01CRBqtL5jn9
iC0Ywp8ZVNindscYcxCYjTMgykpXEdhuwluEvJ+Y/uv/K2KEyeen3ulr1UU/+z6+TYbLAl1IJBg6
QuPEd+4yOZOSKZxB3bxE6up3v0CFjXL9kJ6ROYXPlEyS+wkXR9/+XulmR2V9Kiyu3mcwrel+Bsnw
xXRYeiSI34ifOk0neJbr6RA2LiP026BYMiodhFzqwk2rI5bpqtIrjaswXOibaAkC/Z8qP3ii1rZU
Ld1FIIHkHl5aiZT6wGOUNAeSOCNPk2YQwpy5TLzOQZucMtCPRLkhFv9LvZEIN0NKzcb/Wqg78pV0
mwdut8s8ERErZ8MVxft5sq0oI6NrZb2clgS/RiFeK72CAvNA9zcfJr4JCP7XeYorswNbBPVsdmJo
IwdXXQzKiLOWDn5sKxwgDye0pfo2hT4ue+/cYFk0XIvfKaEWbeBuzztXtF2b2M/yoqzfqWaneyyB
gJ6RPeJTjJCFVx0uxStxLmI3dYntKCWtOz9gH8CSFgPCJk8ccznd7xENIdRHQIZEHJNPKD5d/8QQ
pkL2BwkH4mNNMtbNPWtb7DEulK3N+wuDBdlU8r7fqBhhmNfh8pNtDw8qJmpK3Hmx2CPOg8kdF/le
bCDK8UhAI1XElnVQRHo5hYZseWsL78eblgB9MbArb8gA+39ZJAyJCravT4ItBi9exZCZ5C4Gn6vt
e1gF7CkOsIaQFWlQRnWctKGgP6r/ysrNgj2DmyyVQ+cNdGCz3AsRiUxZeR/kf5GlntvvIVQZGq42
12j//IDuBtQ5DGmO2JxNGzXR7Dyzx6TF/usGVU9XzWTp+9km6OcwnHVgCMtcE4V6wB4ucIeCz1W8
fW7NtZoPB3QUzme/7kjkfFvVCXu5pYHGsfcFr4Wd+EFVOZgZEg0982CyR51hd2fx0aXhxExy6fVH
7Vj2/q0TnPGxC5cbu723fbI1eVjy8jMxnAO7aT3eJjQWn3mMzACbSXu8ymT52lQg1yiJqotpbT6N
eoU7pJj14HXf+qXeYV20vX54CO3dPteiCrNUXL72JRq1+E6cWgcPOoVs4LqwhYFO64rMsnuXE7PB
xUyBR01J8QrTQXPh5CYVYrnUU7j3IdSYvnEs0YNU+1SwJh/cvLJqweqqYCDTxLkolI8JdUEYELwn
6EDX1zSN96eyUMcBv3DMe4UzGHKBH3FlZGqNioeQ3X1vH/0C9pmLr0peWzCrlJuXwRkCeRqT15LW
d4vOKfzmlqDGgKobBcDFWir7V/Z1NwiNvIFnIFD8QfWb6ICuqJt60LDM1ry1UYZM3H7D9UVwY0tF
R5H/j1WqW2bSguAJ4tIeLCbxCeTEUg2j/bTwth5m1tePq+rf985k+ZttwRoG5v47FfIWUMjvbHc/
AHnjn67VQRF+NWt8Fe/NtakMv8PDCqG02T9vEPg2QmQHXrK7XYBtXoBFzvfmNwDUlC2LIz+5DRYK
e3jCQQSicqk75W7+k2TsNAvph47Xs0/ylnxU4fiHNaAPslgbgwjKxk3i0Bb0/SDZSqcTUSgmbJ8i
3uVAdBn87VnF7Rseo3Kym9UPsgUucIuzcOFAV4NNXHrAfbO72Wp1ihIUjug7dzNX1BmJBrFqBbBd
kwkKlpGaXJMpmpCWdQxHxIyTnYgJlL6m+3kVc+oaagrVrLj/uVkXgsWpOYlx7JDGUYXM1yWMOGDv
nKxwO1Ur/yEORBv6/xhoJjeGLaXrGc76ncUOHClNZM1DlYVbZRiZN+2L3xLQppgqM5V/UXX9vfFF
Nz9gFEVJ7wd6sE/DAiSipMHBKdFhngfQjtz9sMEVEK8WnqT0bmc8j2OAUE4Zv0UmOW2uYWObXyYq
vAJ4XdTTWopF7W0hSP794TqMwCcH9kt/eWK77w9x76JTfNj+nd89kqs7zxAnj4/bdXWYrjvZve5V
u5zAGsk52FVHU0n0NtBtrCBUsbGSR9i2Cjb2BGjYWyEalwc+8JTImZfc0eITeORThVDgoboGYvwD
o/Wp7Ih0SrAp1uQZbStFVkwkdz3Ys16kldCg1MFTSnqPqqsfJEG+NJf1xy1k9HEMQ60zbQbkxpFu
i7IGZYy49SDLxQ9XerIVQRzhWyh8ruZB7jg3uEcwfMfM0noDVZGqJasK6Kc54sArByIDWIonZVSP
SzjZA7APHE287Zue0Xuhcz5c1HQ0POO0zRwIUE4046GJssAQzYsix714T0Ao4XnfZxVox95QCiKp
p1UtNfCN+pjHc67uXv77Y/GbJUzlfst/cSfPZS0G7g3as0itkEcO0vUXdKR16Hel4S3OwcK0GmZJ
zBNs988SZeLlyht/pYne1Om6l/rrviOiDJBk8i1Km7bhRuZmPxMQUnvg2xuNWn7RZPMITHpmFt1K
IecCEu3N812KkvJsLZkmQiPOlFdWKNVvDI+2S2hx0vxiRC+buWf1gl8T0wyjI0dVCpAezrCrsEOY
/8DoAkoBoFI2/6fpaYK2pOtpJ9vO9XULocpZo1lqlJnEs1/vgI7lOuqz56fVcBMv5V3o7XrcV5Du
PkUn+M65ZYPxpe7lkBWQFy9KFck+np4h1sdCMkTsnvNMC3yKTq1oLh+4qXBFFwLGza0ROhE3BvEG
KhflUiVaPUpZLfmDV1LL8rAUOWnFpgVJuVynbIq0nEWY+EXzdsg8v95HfTCF8xBzDdcbvomcwuE/
Y5+LK6Lp/gXivwDulKbCifaS6NxVtFb93CxUH2TvHESzxC9si5HDxDzovgIQ/WBWrVMOXS39WinA
pyuT/5KXmSzElPc7bueeNLaJXyZNKGjvTs7VijXT4BtqMb5xGIwsLhOpYjwI80iIjiPasMZNzEep
Pcjx0KES1B/vuvEyQfV6dp8Bq3LgQgGO99UQ1jB3HwCPDAfGPt0It9lcFilkR+PVf/ucorss1/ZI
HUPkJeGY3Whnzkga0dexZLpco/4Npf6QbCp+HACiiOv/VJJhIwjRmGFl0eQkDinwcjHgU4XPvBvm
PeyXLuN7FSaji1nJBobYXCMj5EKCHw3fgbEVQvDuuJshHXrRzK5RAZbAAGwW0NBlhigxCqi9hBfT
VHxeKYfWw1pZUmEl1qWwNE7a8ZnNu37LP+FBMHYdfgaJGSqDTkVixMi/BOHprjN9n0SGhV4ryk3Z
dFMeKFpQyzijWog0nhZdZ0emYKRrRRlgXaNdSrcVQZi3+qRWnXwQBa6C14hY/SQiUyjF8oT7SGDm
jGGiGnNBvZVTdppWZqps88zvJYSa5Zwfv2K+1+3iJOoSMTytA/Mq/cA3hAJNOKSGJWGdM16GuHTN
yxmIQ0jjlpsF37MOrHFUMe+Q8Zlptw1jR6JNmxC9epQga/b1JGiDqNrZbU7wm6FuEgP/Y/50z24j
dZqGVW5B9ArWe2DRGCxdLASTAEfr03th6h2r4DTVpo6LGPRmq7vUd2oBX2wkGhBkZrRAC1R1HDnz
3qZUtSCz3YgYC2iqstxEh24rZ97+g0zlhzBDUV1nTTK4tbLDYlbsjbFvb1oKsZ9TGRe3nAJmChqA
a8/F6WKGFd2uhNTi0mH6GhSKH76mOfpLBQL1tGcKZtAEO6PslzMk8g4wzdfqMjmd+LiK/KncjGjO
hoqv5O90zc4ZIle4wlnu1UEurrsxnmx/iYIvlvRhKowlKxlCEJq9GwpgrCDr244q4AFiITPVDpgd
8ie5dj4aaqNJgQfZnAfW2FHt5xQ81VtBcu6Nfkt3Jt5kgGXGekV3J2U5pGicGTLjdSBOpIRwSNw1
/a5S25cgvr+/Wisb/k1iANQaN/lZTA9A9KNo7pY80PbIJ/3eYXZad8PUAuK1JI+Mxhpi2X9/cwYo
diwmyH2wnM8hIjv+2dVikSWHb+lNmGxGFDzuA5e012WR11f48V8XHFUUhOB7z1uwzsiHz2jeXJn1
SA6Rd0dQg7AB4ghhOi9vNSuALzu9LlmxYkV1pZZO3ZuJ3qqOHbfq16e3/6d8luUZG/ZRR9ck3dp9
pTv8DlVic9l4JFMXVq2iyIEovfcSdAn8cLlPRjg23xlUMRp6qI/XCJbFtODV2DJf1MLUIgZ6aiak
QxNFpY2PYYSW1LB5OClLgixCPQ+HmRmuClaNbRhMgSVc0mpJUmYsN59MtnsXUICu6T1gKtA+I+U0
5Q+GJGnm8Ktht96o4G25tqK/mZxaaLJuA5ZE7Mququ9Z8KIbnCQrfeGzkKsQkYz3GDX/Bkc+JRXU
DlhezBcgHy7CBno8Vs2zc4MFYLqvSAadlkueSu1LfnHqgKitqXAFkMtoK/HFNsIhOjXKOB7IhcHc
lMVK7pur9U06D4YJhdeB6yp6QQ0KEK0DXoAmAgv90Fb78ppKvWvpYEBkPe4cEHP3mfCb8upu6l3e
yQmu+Ur//DeDZGkNy1FvfGYC6V5LdzrJXwOd61GTVaaiu4skn0/P00HT7cdoVzSq54Mre3IFK7/H
zcuPrwZm93/qMRfDKIR3FRQeJL2M1gAYMDfD8DRrQz0H1xvYQ0+VfJOLNmSLn0LZgvOl4oW/xcg2
E9MVGv+h4jng9X8sjF1sSBGVWp+efkS5hpY9I9CPXNWUdj4okJjAdVK7zBgb6rdcyvzdp3KEyxBg
4WtHDb6yfBkPVWgQOln0nEULy8PD4fx8+68G9vi30VEyk3hjrgfUqaY6oxLxkUIb3MX9c24tNLln
G16gjGnjcQ/FlfKAQbgm4BI7W0Mwwh41atM0l3YqkVhuVN8oduKppheiYmlnl3g5tAA09vffjD65
+G8coX71qQcy+9ON/xEF8XU3j1IhVHn9k3HIUNRf+65ghTtZlbU9s9LfGL2Yl/Xxy/TJhz2h/4M1
R37QarDCGhBEB0sK3Tb8uOerZDME79Bz55Z1nOZxUaVtapkItdsSHbXbIAeV1YX0zk7BlMzn/lj7
g9vcwCn10vehwj5uqhzGqmUAUUr3C0Qws+XxbIbL3IPQqrH+8iDUWL2ZaDu2AZiisAiaJn0eOO1c
2ta7OLCTsfyqSOSvEYeiUcR41ES0RClL1BXYTZyVl5Vy5Rsp5MRMrR4CDyOt/jOGwEuUFXLVMgit
+sfeCcUAByOvp6tFUDWbrPI72JBHoFCR3YUBtGUCPLkBloWyj9PU6ZtJCY41GzH9h54GVXrFlrPS
x5y3hlrrWONnTWI6AWMAPESFixduIITX/yZFxNugs3eaFZFZt6NtVbC8EiLr3MY/uj72TwqSDkj6
FQLiJJdArgHhNUr++Vy8ETvllrUwXOrF6xMGUCBmr/r+6NOyPFVCR4MRPaQWsLlchYvFqozgn8Tk
NRxx4LkMMNklQOB0De2oyMVCfxKMHsmG9ocyslWmZsueGob54hC4Z+Fgimb+Ar22viUH3atg2NNI
55Wyy3rLhXdFUi8PGxUU6m2mWv+hsvtwXpZvdhWXE4QHq/bBFrE0T0VNCxtTvfz4iCHg4hRIPL+0
CKK2hAOGrh+35my252FhGv/XtHcfs0vhP1voJIS0YxQVoA9bX7MjG4PI8dUhd9k+GuzwEobVcn4o
ExAwhJsJX9Gu50q+p7JjQOzLxDcjmvsl+KGEv2OF3WAKL9ugFdMSWqYJqO4UQqTASk9O9inmDOEs
lwHNp13Td2f6KdsqlR2q07nY9X/s6uL3Vem8ON/5tmbk7/xakm9/wFw3s5UMRclSZ7hs5v++M4r3
obV1B8NbTRl8Abu2m+TaK82tHuacnoKJ7oAYWzg05xzT/hdnBXe9IuC2Hh1gxvr2zsYuo7J26Joj
bMx9J5+YfVTBDB1E+k3033yxT9CHF3iXZzV8PbGrHWeFNjB0TnDQAsnv9+jqOTtyhl690iwzWiZR
pwH8REYlXfUtQ52JGBGn/WudgK1rEY/u6b8hOADxmZbQHnIO82IVlA6bZMYFqGp2/8sAso672I9u
/WTMna0K8iyxhwFQ79HJpDkM0HwFSqjF1ekyrDmCxjlydvW2w0lcWiLZTAlxe46+Qp/sRoPcOMXB
TfrOa8iaABhbYdOiuceTs7MULeWHVQOw0bgE1d7vfro/hyyhSavhXrOADGFsJEtFTBL6zoLv2MiJ
2Hk1ADt/zXjPqttXcb+P+L6PUXb2NdyUP5u2yrEY77DRmGYYybq9j/RBOsoj+yw93baCQjgLusVh
0GTNzWAt+VskSlxnWNsehZ4ipRUmFm3DUz2/qpC91T4u5XFDi7zdwjozr7LDz6tShH7UJa/9gjxq
NSyCKFQLWbw329xoMZ7VdA95x1X42FsJgwzNKmpCy//saRLdJJ8FYsQHmZEezLkSBWOi9FBeFVJA
JioOAqkfyDMtw9gFSl0gg/qL4H6ZPufL6V1ixWFzjoVGa6uVJPo5/V4lOYqMHy98ijHzXF3SzFcA
QJl/G4ErPQYzYni2z2OMTmLBF7uCO2+KJFNzn/dwYqQDJE9qcdR10qZAhVIVgBVw1IM8FEcNCKeL
z2wpOH+Yb9+OeMzFHLakASqOs+M4OQ9myXN1Yb+UnXqIXrweWf76+cp4+lnO7tTgzRfWsI5KBpHI
Dt4OggoR5OTfktyOpHRKPjS8yoc94TOIiB1oMv6laGecqnHSGUDcykWnIQcAxUju+X1rwPdiF6FE
CP5c0NPblohkfdkl1Vv172PVOgeK6zmDECceVuifSvJwySxkpdc5OLIjGSUDBWgwqNQjKg5gd28e
pl+qCr+5S1gW7vjZ2cAs4guiUAi6GlqX+gqtQy7Ord8xKbT7RTeoIyrl8WAJdY+zCIxDzHf0P59O
E8E6XdfGJp0da+/uP3hYdOdB514PZ59YMwiv6e2CVochDlHskmShgP7xueBtGHfXB96Fh+IdN5mk
EeYgmgppNVsNVDE8csazbPcz3jxoW/MIzM4v8M7M2v5BgyHan9YT++eIQKRZ3nR7TxLJnpCdQumE
TrfL4G0GUYSXudJNnoI2OT3rlAqgorIQo1YzklLHFIZK8ep4fWrmKTN+21ga5/aGV7CLW8wfcgj5
pil1JCZ8CB3PLJQKCvRX8ShGBws3zdyE2AFAkH3DoR9HiXrQUiOP/+26rIyFpPrAmvUSypy1ufdq
CW6MhB5duEkImy4z9G6AmRyvEjJJa9JnGdNk1b2jTcXvRdvuaJm9MNU3VK1oOF0Otx4n0mYMoZtm
2Z619XD84n6G5STXirUghiPMLljndap2xu+hjJm4KvYEJbv6CA8DWWzmYoYo4jcX56GUUCVWsZ2r
81C47290kaBz9iPV4CWaRFxZn1ml0pqWdXqUStv3UjVRKPfHTfPicGfG78WPocb4CCenD8xiYjwg
qSk0wAqxQq7uD3SS1FQBHDw6+O1S+L057AdOyxpHhkXnBqT78f83WSC+qSmknUXrnUHZFEbSqa5h
DfHODdqs4SyUcqTisuBLqHZWLgyE5NcaSigpvrBBitRXqnYkaX6TQyd+M5QEKLd8VFd1y9MMf3G3
5eRp3D/agB697bJDNvxPketNLav8TxJgL10YJv5G0fEuiFjl0FXcgaezU1/15j4WLw64q7IqtgB3
KicPSU0iyfVEtCSN3S5Iz5ncI5hLW5hJyQN9vistsCN3N0QXfY3ROQoMW1/bdhPTe6+bmibHz/aN
OZ28iTkksWBa2Xjoqo3nQlDDw5brjvUZk/wNPYtxCu4ph8y/ZhPgDpBXDNoKHxY7kFaN7A1nZl9d
Cn7naDqjJ/FMDxGkmgk8YdvLWpUYDG5vw7eohjpRq2GA35Y8GDqugd2FqyLVPDGE52RheZA0GxXi
OlujiE9OXZz1vGSzJNPB2fFkSGCuYi5VZDB5OMsolOrUsiB6dOFhmh7ekIOSAkmTM9X72px01fNc
YhR6727iXpab67jZg8S4vHRBNnb278uo5Ut9g+O1gV2PZ/k3HEZSCVIXOjd8hxSAieLU1T0BZY2G
8Hw6DCpZHAayaFW21skY5oMBIPN88eQj6C2JVuOn5NKqMsdUuxa5oCCaJN9vAh6OhmsIpxvzEVzt
tklni1x/SEnM8Nke8ApjQ2p3Q5FtLUHP9TmjYdXMtqMoxN/YBquf30Hm2PJdAP9S9qhkw/I0YCD4
Hk205b0qdtAVkU5joHUzQTHpsgOsjD5Gpml3ia2VcsDqw/BU3X3uar+7JtbjGY5dnbWcvtqv/9r9
4W6JLYlJYHYPDvscglCfzMZeF5/nHb5e0hlaO1Q8HA5z9AF4ecLjKdjSIlpsaFWa3NgQ5sA6G40Q
JUEnXAHCNTApus8B0k/ZTQzG9Wr1lDKAYPKncaAmf7BguTnGbYCu4zaKB8zZ4v2x01bz4p3Z4wFA
U7P0zKYDySjOYGXxTtekCNaDER1cqcm+pBwZakJidUJDYzgiZqv8O6vpkpBq1FjvLvByZudACtyF
gRl2lTu0FjjFE7fzylnjv/BtVYIQx1efisGb4qMklZAP26mcoxbbWDTPsrzvMiOpwhaZr+toVfiZ
GXKRJrYOhPS5HN3XYb2GbRUXoM0hzbVD8gsP/Ig0rBGOpuCRa31m3KCQOuQaoK/nQmHXz7qnQwLA
sZRj8vdOrSOOzWWe3J0XjqvwNWDETI17YpyirOnb/t4Bd3CkCio5Fmzv8NKpegA+JEkxBnGdFXRt
eEUQ815PSrtS0sHc6/EGSvN6P4blTSefyDIdzTWktUboQRx5BOX7kKDrMCKUZZTv5qab1ELu9lPk
0cxsasUjFJHqxjZ7fgaafNVba7E3HdFPsij/gx0nmxfXT3WjBXXCkITCdl4eCNn+g1GTjHIiJcdz
us4PZW2qdxiMWoUc4JbpESjnVSRU90C6hiknvd2wcmWdMhHN7Y0gdOcbVYXscc5Kc7BjconpVEGz
LW+u9dDlx+rLIx9J/Cx0mHTRszlUlraE/+D6zdW6Q+3g7CmDSRVP2QVEMCscZHpGKpGtK6y2ztq+
PN5zWa9lLC0UKXY6xHY0idLtAt88unIUbh1v4mQtLjel5bHXMmAb66GUJkt0pyJMDFhFDWUkv5fV
DCfcrBvP1G4Hnbf2UrOKjm63t5bwzAvuQZyHkY/gG9ai5zr2nB3FS1eoZgIw8pS70aRFHjMm/TY4
zmkWbXDPm4KN4vZWWO67ZYTpFfi05hgyhWJmjxEq5yoY4nJmmzbr1aHw7sSp1URFGqNgyGqusLJX
mOTrlAR3kxnp5OLi2Tbw8tAa45uvaa/hbyXHAQf0EslsZu/wTY/3f7Ugw156baoM7+hm2HpWJAV0
P2KDfq+tuQHYRYvav/gzKw8TM6ugzwhw3iQiUE69L7pUYfDWYFVzJnJsDosgQJ0NGUAd/J3Iqtk2
MxwXCaRPyQdz/ZyyEApGgiqWy+7HfRiUchgZjSRHZJVXtdS7DWdEAxBatEBcr+IbANceOnOtCWbB
TXV3DyXSXI+evUOcnTGb5FNHADysOD6i0n3QoPc4v7pwUru97G5h4g4IvWBg9sS5rEL+1cI/7htN
WylxerSCjjpF9G8CZOuu1HyfIr04RaEAV+TQta2/u9z8m5+gYmNKqh3u0/gQ+yl4mlUA7Ma4EcCa
LrKkMTvoxRdTYrJXqb2lTwaJMbKPLt3M+sLXGZOSSik2Ip9f4YGeMCwEPJTHBq86t50co8Cj3ls4
YG6kcwObkUI5Ax1SjWLn1arprw+pdQ/VXDrhx0tzp4xnNb0WAm8ylt7Enyj/jXfoykFObu5nOmlB
9O3ZT4/1nYbBw8DRPfP7L7TXvZJpCUSGsUecoFMovvg7R6Lg9QCnu7xqCptnpN3xDPrdjT9Ly/kP
w+r6HrGdqA6r2rKK5wbyH7rbN5Y23aBfJpBNlG5tW+xKfF47XFlT5p6NW4OjwhkkyNV6v04xn80Q
BAqZ2iw9UjVwLSqWprEhMvS5vQmpjUv+VPlI1eEwNEWmgu+G8Ih6q3MC2kwnTkzhResDqZaXqOSy
9/yjGVLhWuH1JcGzmBeRuUR5+adrKZPU5CZ2HphKrBj5heGNH+6HlkiiPN7zPVwi2G0fDJeN/82+
0DxU4tUE/16TENxrlxGsfBWiMDAVc5qim+NcguFwoHapSBP1qPPQlG9/GWPR2wfvg9mpvumBSjEf
9VflsPWb+4WBozSnNgcOILSt/Nyg5E3yokCiprzuqcZv/1jN9J/CU8hNb+CdFzSU/fUAc5VcLHXA
dCkS8+aruY4RNa3yQsZ9jnt4LtFErdZEtEL0Pk/6ajuqAeEtLAObSSeZTwzTNFXn/3H0Tqgx9CH0
iluGlAUdSidthcYPQScjZRZlCj8NBu+Kzfvhfz26BrLw8YEEtEXFxFOeCQs/Xwq32xVgFEgT+AWG
vfktublxFh1iuUSIhL9WoD9dJ392DSliwUYTkL7CKl56hX00qIxCn/S/wr2vID+HRFQMxHGgL3sW
UMSmzA8JBc04CnRKIcszuOVSluF3EVEHrV9afoqfdCs+ro93HLdAvlvWZ7jaJA7JtPTgNz1h+hiP
mcXyviXkQPePzNmrr7HYGgTGiB1Hs/hwsrHh0o2zwnDQRi3tgjDG8UpX3qMHrE6Vr0bHtayO9UvQ
W2bi3f0dZ38kr7Y94dJKv6dc24YxlSeFqF3NQaBZoUBRiAR5SMzps+OfJrtvZu4ffRlVyVSpXIyv
dyd2PjdvbqlL3YjVqIeCSK788KMA91xhi5G6CI/Aogp59tJP0xrOqZUODF4mS+i3SYxEb13B7Ofc
8eCoOWm5Q6Rm9ycY0GsZmy4nGOuE5x9FSE6Rdn7de5VUFN24HOnuP4ZBRABO9mtedzHZGosLjLKi
XVSm4VYZBrc+J0xx43peZPeeK0f7d29zPXo24eedI8g3/GflJcx0OcrPTpqZEHNDJtyyn+scOP6N
e6xsyIvd4MvK1edeYcH0sUgJjn9R5QfMUTPPy44Cc5NcwPBemSRYbLOUZajG0a2ekCgTdhj2Og22
hPZFJa528ZhSzQrqxYsjAFXHrXqRmz53aVCRsI7vnkfg/psB3yemYRIAPIgR6Xt94N3SG/5z9pAU
bRUG8ojl3qTvecAi4vT494Mvz/zMkkRkYyuMkOv/wmHgXATBjn4qrfCY4jEEvAOZuYyUwgSFhDh+
T4q1hfjzFAwL5g+XOTIAB1UU7x0VrweQ5+7PgXKUbXNcVBWFSNg8s8aO/8CtfVXci+2WGtkc3Jnq
Pim+bnfwJc1T47S/lHhp1SwV5k3/ewIHe4gclwWg3Dgx3V79Xu4pLIakWik4byZD0AqEgaC/K6ME
KU4LRDzhAkFhIUUuG74UkQjQ5CzbQDCvXGeqt4yEFXE9sWVzOP2jxe6GfxLLFwGd7Kbd+IQRUK4Q
SikHAy3od1FlRUW2lW5lUtqYhiJ9J0XXhbpYux2fAYUBltcEFrrYZeFpRms/6sFRoQ7+Sm/Seacf
CyeRUizs7HSrmqyjH3ihILgwZwcFEf3ORx+LjAAi5DZxppCBkS6/iAoCl3qXaoGuYNa91hI+3U0X
PzL4jW5EpAMuM4nhERWKazi/HGvjqD35hbwtfxgwCu4GtMwMZzmLUSOQIlYeItIgbhr6O8K1Y1iS
lfZGS0FcKTvJnw5/Ju77MTESrMytzYYJ+8R2AHF03/IgRXpLMjgsxx8RCyCL9D88TkeQ1qyuzjmC
nqMO4HD7+oIJIx06FEKxTJxEuZTSZYhkr1mHtEMUMS7KwwRpTCLxTvMvluupoVMycyX6AUAGxz51
Dtap8hWZ8gefVmnd2knbHu+XqCeGE3iGgcODDDOCuLbPSk7GSImViefSISEzjixVdAImacMHQgBf
RvR1nQvFiV+YFJU/QUoT6DXCOS9gK6VgJKd92OusPx8tbBxTsb+SIC7+mX0lzfZHTxJz0UPNjI+Q
JJQMXuJY4s1R/hoUM0QGKd3U7SmF6ns44A1l0DDN8CXceL+8Ek5dObwUCo6FpHfXnmXgJL/u7Rfi
GJN1lyePyvYPp8n8Y3sSRJ6R7MUxm4CisLMi6e4vgpOdhBRgG5czXTfu99nzSbuGrR9IVNN2D6pG
083pXdxxYFRZqpPZAajUcKkNH1QoSYHyvzz1OkoKHJ+WdNLAqKApEMz8jqdOuUjitXgWjzhfmhXp
SQ50HBXSniUWjaqOWQgF1o6oRt+vwcLfH/BI2ZV54WeJK9xUPB11MLEyU1SW/sC6M66hI1SiW78a
l7NnPPm46E6jK7M0YqlpUZwybYhJmbe+vq4rJnqYBaACeX6d7tXXhtZUYLr5jDrzmypP34L24Ub7
8wwhu8SGtJ7J/68a1lp/7fGwXuwpEUWBUp4Nn1eqNoeyG3mhJw5b3cU5iOriTh6F0PQR+3UqQMH2
YG6Py993SBuF4ewLENpdrowdnDO3oGs/8aVmsKli0iOGNIJp7Yr0Pu4Wfry/erO3Y/FPcNz2CwPw
wHs15fjmcOVSx7LdEZTfZNc8KZoDaRXz0ukX7L6PH1qaMpesz3u0oKWIZyOAX9OEf450KDremY9C
3OJ6dGG2ufbwkF59AVrLFWxcHT8PuRbxd/6/Sqjr4TMobITf2ZgufAEVI2o+5dHS5+E/hm1LB3nA
ufrY5K/hXqwcggXhua43COUlLJjWTUwCGE7h/fs2mxDFh2vhI+BuwAT3alirMZLpOBIK/63xLs6W
YUrSbfXGBPcJPXX888zeGh9cRpTZt2/hSlcx8BNUip5U5iXgmp9Fa+xaK3188kLUbRZOrMxDvN0y
yO+JmXr+n+bkQ6DS0UCj5CLu9smfF0ZjI2iKUvyReL+eofjMKc/hTrisxZsCp8xlgx5Y5S+PR5kf
WFj1Qaus7KDMbwVyVwz15N3iap4uj7yAl47Dbf8HHg/lhzuRhV7BdxBMN8MxQHAsBEwkShQUAdr3
OJX9g/FcnE1AZmxsk4UaZY+rY4oYHbBEnOwne7q8Vvq7S+b98YcPF/s5pjg6xUEZJu6nOc/GbafI
SVDo8dodrmI1pcSY23oxZTVoqWFgIsCb8wf+TsAmV8uykL+JCwoIajju7ClJ2hlNkulc5aTP/qkw
wZ/2s9BVD//AFq2IxuvE3LryW0BWqfQm1KxzhK4bUUSgjXdO6DYIj24y0rNcGODqqCiptUs1O3M6
8GAq8RirwagcSvwMuvTfFLKoLNtUEYiBZ5K2AFgXSQZcSAcIbocIuXosvUZoIHJ8vHw1bK6LkRev
516OfI/6qd4q+S/P03rZuOHkgtTB5V1NTYSKKprkBxsZNuDMNikKxiuwpDA7zD7dySiUDPIbpi/T
E6guYqvfpg/FW2OBG0tGB8hHSuJZt+f2J8dNTfO55AOra91PWsIzezrMPX9uQ/sdg+YeGTYdbiVb
EfldU+WZvDbgGsfL68E3/WOxZTrhz94td/YdSECPzppvIYpFVun6VqoEq9N0pjgo3WH2WtoqlF0G
pO2A0hy4DxqlpCcllYTWl4GBHuTjnYkGx6FpzwEdis3ZZSia3Z58R9ETaESumwJ7RrxZnziRpd18
2rMHMvCesze/8HcbxUo9u3Ksajv/3qd5f3nHxHPgg10/olKoPq2TfjXshRN0fIrI6YIRUqHNn0s6
ETytWoAeov8oYFYcnqW7cfCA+2UBLFuaXTNg7DZUSK3D+OH4b4KT2KylmFQ9LUQwECzB6Sc/+8jo
7QBmpXaKEgHnElRvLTxImQdkZkk6ETdL/bfpuzJxdSNN4OCmAc5C11CIH6KcY9xrQ75BpiEqC9Gq
mS/31kddYfNOipmz0AG8kdxwric4nHyzYInfHDQ5bFnIgijd0sguvYgOxf64geqZflOh50XKPUSo
LgfB76eRUEGPXpsUwSozz/4dtWLDw+FbLF8u4BVv5pScZ6kK3Fm7uTzXMmPrv2AqUCNG4TEMJA7X
2x0y09TevoE/7O27eCp/AuUDj/rM8d7ZJSG7WHdzyk44Ap+8fB/ZLypyb3M6ze17jKM1w8SOwB6q
T3D+uQZsOzVpzP9bL8cXZpRqhsn0Isae4dRoIkswfcDWyGHJUq+QB/n5XNFCpj5Es6F/t9QBfLT9
lJfLrP/ZQxLcig0P/+Ke7yh2CLBSEcUpbc8cEN78s6ZV8e0Ye1E8RY/WVDZdoSGZZ5Fn/O7TEjoS
VWYdNKXezjkICOBxgyY8GJjXjlx3MhCRZdyASKzrpu2AQpTJ3ztDrQjPxrRyYnLYy0dr220raWmX
6pOHLaESEB70Hdg/tvBCA7vmw4zxc3HAqOivJG8FaPvTJRPiEzahb5i+VL2UY7GaYTs9wtPA3kRE
/svqldppfJfH+VNBR5LQKerIu/GJfhjIAyKkT/n6fUDArerGlgP9mJ+rBJXaRwmXoCHXfsYPR+9x
JUF6SfHpPps3P1HHG1fswffh1kTub6ZFwgk93ojkVZ+2oQGGxGej6DCq+XnYLtoCHE9tACF7VIAy
+SIlq+9Ncl2r3xMVDClst5hQA+iz1SonuWgG29kbGnZzhcK9gnpHmIkNLvZycq4pURquM35DqIfn
WOfRM0KuVCkdxBOa6H8yCqLQniGtYpogVo2CNJYD54GvqCmm+wit8JXJI9FfESTSim+ix+Wa46bM
Eo0Jy+ByJjX5qRxrKmybTZ1TPMMOFrD/1DxMToCkvjJ2BC3sIN8K0xbSbL2EgptiPCjinH8vNj3v
orqsOwuR37yGiLrk8cqF/JKuLctm4KwQhLNJinhwcxQVHeCAEF28yDKIcR6xhHh/LihBTJo+/484
wW8A8pMSgUMurOSUEM9Ez0uxZM4gx6VoKFuYj4rNO/qeN91ZU9cYkXm/ih/MdUj4iwRK9dkLzY9P
7pNSHHYuIbR7gvf42BMI92r9amydC9sXocIQilsnS91Xjzrl2e52lXE3HXSsywVEZfpqwmXQbMmR
GEu+oFC52qpxU3ir4a0jXLwVPhllMBEIgzJyoeMxZilSmG2wYb0WOu5LbgOd9SEarx37uS/bU96/
byDIhc6r0kyN2PgGkedsHPKXszIThAafjgq7fMm6H+fbdqdi4+0pKcQIKE1cLNE284qLsEO1a51u
nj53gVotmCbLAK+UnAq+n9aMvsXDo+cpQkD1fKMncQiPqOXW3LI775hkp0iiBAoROPc/lqJod3ol
mRct7/ydEfX5HTifjW/CiM78XRDAePamUMSMecTOtikpWBb0Z5SPxmsIVi84pLtiVDoP2YR9v+T1
xXgNPsAE0MkUrOMtHZCs8lt9D/tlrupVtRbVyCrq8mL0cRksjivSLJsxi9HMdgxIJoEkI3aeGzib
9AkXBhQ6VW4xMcMgmmR8ICakQr7eEkS186pnvTWkiWFyKRCF0lPBeUm0XOEdWMv102F5zvPoRlDW
KofdhiVPIv3IDoBGVRGzi+rUKeTk6PhXwr1OUiFEbRIYwpw5e6VIeY12XbeMUVWXD2xa0uze9lEG
i8dKsecfT3Xp+qDXtsrZwAN1hXvwVWo/M2ZQvePTdns1ePFTFkul0v8T4/vpTDL7++Souc8Bxfjt
pWjXFr3qCfgLv5YiWf29euktIuM881vTAzqL7dCm0u81PosmODqBrGUOPfK3bXR29HztW+BJ/C3t
bd5cWllhsPgRTAuacqKfUpOWQaYA8y34PwKMWm+wWJtdnDHIHoIO5KeXlf1FWsBLAtwsNJna26W3
zMv4sZbrxq0fPBP1GbBNBiCF8PHgM/Z3khh1gmF4ky4rsvrkikARGEo29n8Faj0DZCWwQRS5H6Wd
wS2asT5JgKTOml6BC5nuvKirGM4DU/QrWZMIdQl9P0p0OHB4qOR0a9qvtoQNaxLwYeeGKD5uUsVS
7DUkjDF+okGmt3zjQKinloyttCYWwWTL1zBMcqNRoIKo5Syqe/a+lsoc2k66jSSHoL5SA9tpoWt5
Zoyhuo6yZCl2VpKnq3zjKVxHNnYtjwHqXHdzmCehn3LtxE0RPx8wXsMi0bCwRZF6MGoidJm6NeC8
Xv00+NxSUMEGQjp9/CQPeoh5EmwjGCMLDGiruMzQpyyKRFVAxyVqoFq8a4a6ocKkk6jPMbg8Otu9
r/q9kd1ZfWPeQss2z4o8QitOysZE4rIxJPepEhLiyfqyu8YCUR2oqF5FpjySzNXkuwkXpwt/rZsZ
PGKD4vo+np/IS+zgQq9b8hLaek9jvcP02hsDUXyiBkhWl2qplKeNUEs5OXPPOzXIi2r5re0LSoCk
C+50hmZ1RntN4GEk2oik9IA8mCkVge186vNqyoa4Rv9ecmXRgaJBkKfzeddIRdE1Yo3pXuh6WYim
eeXWfNMMB1tN2cnHmKBvlNm7SOvBZPWWR6YSff5difHGbz6zN0D4jNrQO0kRwJ6sqrdg9VXDS1mB
lS4P1kROS1RBcDAE65XzcGIceTsrCXTooGnkNKi8Lqpq7cMWBHsX6wQ0QPs1a/fXAwVZT9xefhQw
JeKh6RUrGu2xpEV2EOKpQsAo2pDrfDkRAxnCITIpCPR8bwpxSzZuKuO3i/eEkO7t7UK/hm9q6AFy
4boAZk71pfAfrRbOEDbGwfffaq1IwX9QeDlX67vqypmkN54nhogugugDiv7GRWxICn/u6arVVEon
3b/xjyrLtSqDxV5Hjd4gps/IdGqY35R2/x4Lfksa/CExehKgfvY5bLEtntd5iFwyrrZL7K/phsom
JQq1nB9J41FK8INwh/B2uKc93eVt9ZqT12jvXJb1UNybfg2xwmWP9RtykO8/EALPM0CscfCW+xoo
96qbUH8Dxsx237VeEPRx323/VyYgNTW152gJG8GcG3LUT9seaMudDm8/S0WKeRXItfCOG0WTcQWG
6xwXE/w0Z+OFb+oSbZqh7ot5LFl3TC6eZ+Vel3KI2UEClYCYvFgP0slXDMaWn/cDdhzQuLWXNn0Q
+Nu30PfZ/Z0N7CG7OIkmo50tbC5uEinxixobQdFcvW+eoJRqHa5lKYesNlV+WEEcG8lTns/0K2Yp
l2NZDFgdjgV8XzivwDlHYsknPGBRji4z/DdHWdJObA7aR/NVIBjWr3cffcvdz9M+MMkUsnqz5YfB
q/YT9x7h0JjTpIOsoyzLoS1cz0ImT4uRL+rmORhY5VSAqWQ/dCvrZ3mckI1t/vkZ/huKYW6L6rVu
m94wyR9jTok8HPbY997927pNCuSBOwUJ9c651JOrPYh8okGVYSFZcb45DbTdYYKskD+MSpEUEbzg
K7X9heowHTPFL98Y7zpxb4P/0Krc533MvqpI6Zl56d3rPwgCMd86QnyXO8/wt06fb+HVNl+IXoPM
ljWG/G3ln5hBmNFE8yqogQR9fLj0bJrIk1gsi34jBJ1yrgRbdccKjgnp+aY4YNs/GBgxAJp+vNcJ
bjn/2d+sSBtJL6j7DZ/ZOAu8Q/rFSiG87bw9uPvbOkaLvEdFlqtLIgnsIYpG2SgalFNuqC860Pt8
0OxHqcCpXLY2AMzryWu3QTk4IyeTlkezT0yTmhWiYQNoejqdwCZsT+Gw+Yk6irKrL6miKLi+DBub
+EPlh5umGpbL17SJk+eN1o7E0DEx+11wKkWxosIMKnv/lKAxTPzWUaw9C6a2h3L5lbizXCG6a7KI
A2gQaUMZrDVAYzJiSvNVB9Lcf7SQ/bi9E2u05YnNPLoa8lR9sTaZklMD7YllbilgntVFk2eHxlPD
0F++wSXFlPo6WPAU6wAqEjP9AXy4B7dUYpUaLjOq2gMkdklAFf7uuG+28acEfnoSwOJ/7b0/V2mo
aMIH4QMZ7rpQH7y9z24f/r6b0zP2Ao8qvQfRTbBxyXkv/h8cIlZnlV+Ur9oRsTD5/y+YxuXQoXkz
552Mb4Q7d6gjDMS4RCtnJsmF2FA2wS9Wx5/DAKutzoRMjWMhrp10lVtnMFyaBFDZsKdeoyqFwheU
2Sj2tJtdn5abY7+P+NiWzRJPHsf8r6Myl0CYQuFY8TjqhmiUh3dP5aWefnQQHHTfru07eSvkMBUt
TiyJhhunO0sCDucIXx34C90QUsn9PisS5bFYNvG29ePkYHO3kSXJXmHIHbs8hydMef24oSIi0Dib
/Z5HWOtTlt1Me0jVYa9OEve0OMdq4kkTB/doIGvzYTstVBdvEYlCgE4Ta7nABGm95xaQZ+jQe4VU
eZCASfCarP1OLW808JDYta5y1B0Bj6bN8hgCJevXm1kVhXJYd3/IrizoP+eUXGuozbPcjasGff48
m5PS2NFKcp68dV3vIA/hDwPqNXIkCVB+UA4/IlPzVbGIJgtjJ53ZDz5gLguDtAJSoyz1db3o9kt9
bdSFcuwmXL8vOFfmarOeoh8YXvMxYQwF5O0C+tUyCMkV3O9mt7pc5/PyOS4Ypk+rSaHuRtyHEruI
7DmM8Y2VflCByr4P300/kYixA+GLTY6L1ZGf+prHD9+5mkdPUpRfTIkOW5cf4lizMilWEpy53wpy
fqUyXRu8pL4nd0AEcewP+Kee5rFYlgOxdfUV4vud+dwcPwjsfpkJWujUvNJ3BYdKMmALyE6IbPxB
clR5tH6XfJ8hgekrcsHPIiPHyOh6/RJLMqGOMUVGV6h9htrfS+icvQq2B0sIKjZjrEptDdBy9/Nm
pn+12CVPlcDFAegK7XY2Z8Cw1NcLYA6yBH4yT2c8vDvD+rO5pIcPXPoAOAgUpT5C7c91/87aMAFg
Z2uqjBPp5rMWsccPlCIWnSeh8wubJK/GB955lB4bIqjF57GnrDM6Eu+E4tzbjaZq3O7a82AmRchE
IYlfFQJVYHhtizv/ufPEu2LwpIQmiUEbjufgQOt107EwycJ9abVFj5bZGSokmRljHoPIoF6rd6r5
dCYEoDFdfJaODjp+f+KuMnDWHMitR1QvHfW3z/08f6hiqNbPcHf1FVxSOJwFNNjR8KmUzkicU2Mq
oQ7N1qCvnUcff2q+rZvK8V930a1lxz1r5dU2N94cyfQImDEfigfw9kHKl78EoRv4f5ddpaEFSHCo
3KKoExTj3k11ALuq2YWiiSHVhvmjU1x1T4x2sEp3zCeYd4l17O5SBmakqFavqOfNQV/QwGT0rfSF
qaMvoSRfMYPusTPVoKuZiTXnh8V9vHg9mcjQtVsfjwmmEk7XwI6wVLXeCxp25KFTjBrjKsGSkwQd
67llCsWU4pv6wyx7cUTy+Er/WulZOohpTmUVzAR2UJPvGdVhPok+8Y/AAnIn9WSe5dWk19rNOQFA
sZAOWZwzWGFPhGphZukCsw5GhOu3Z87eSIK9e16ti3LGIE446DSupTxuMxQFmZBHRpRikTYfoV2+
5uQZuaAWG/GyVslzvbw5O8jS4yjEMRvFTR3Bepy4SxeokFwFB+67Hxscf3BICixQ2K7jjgu6RGLa
brEaqKjSrN3o6Izpz4XCp1DAwxH8q7a2XnnI5CaBCOmBKRDetN/isfHfLQeiDNXYiDJCMJteuBkd
+IwMrr1gr9xeOjZwMxDPXWAlQp/nNVddL2AECp8OU+Nm7VhyJSu+ZiuJEACKblbXN7quQHmTmSxl
LFNOhcpSmG+ISNLTebrSOSMAy/cj4Hlt8ylE5Oyqh4ePE4Id9gYeZxV5bCL47vYH54sx0u5Nwa76
/AskXxyhRn9Q31Zd9BNiQLLT6diL0kdJ3br9+vqF0C8HnBb4K2OgGQUVFW14xAuxUG7fVta8p+Bt
OSmctt/UdrM+pF3eI5Rg/6rlXTaN7EgRipR7SvumkWMOOrl/oBF/VQxXi9OIaewCmrEJhydeFN9m
Vx2rqtxdPC8TxHzO+vJ0pUB0yW9vGbudyjjx3NBJE2gyI7/1LN+myrSyUYpY3Fskkm3FOmQCkM3O
BlsVHrxmMfa/zEb78/HewP1n4xVt2qx5F4SdYmRxCOTlruIuRtxS8IncFs7FvOJ29XiirJlseMb7
Q9snFhzqBPCB1agZ7PDNsqxfFcUFnpySotzFlOdkTOg+wrtWAX30BKIk3s2l97GcGPlUMos2nQ8t
MlFUpKb3xTEtsJPFLazUPpudCOXyxZmMEyLQzh99u6UZLcXqiIQYK2CBictSM3mQUDa7bWrKGBPP
/6FtQwp+s7NoEJ6OU16k7MHkhJyC4NXX2XZDZ9MWoMJbbKUOlvUlidy0di4RsTEad7SVtGzPoTYv
2mZiWdGLcKQUHohgeTP8PALWrI5ioHNFSUzj9PccbmpToP3MrJflbpFmwFwPIoVI6UaJCKOiU9iT
mPX2LnyrcBtd1rfRIUNFmyBY4ReOscAnSDC0xChVc31pY14kG7xS2LjKXUhlDckw3g2M4SKgIej5
SZym8v/bMP1oObyR5nZzp+bB7dFQ3DMDZrZ79Mx3u1Ess3zrx/zovlmuOD6mkX7OUjxoWvQ3mztL
prUa8uLvLYNdQ7n9MkPYltfpq0uMw3/p1jeq6JjqxndhxmJchSggVZZPdhURez+IE1UMEFNSlnb1
6mededs1LS0/s0zOmM/Cc8h+ZOecFU5munixMa8/twNOPkzfPvRupHsIfo7f6Z93ApEdNvox+lO0
CQQLEG0ioiQmMGZayEs6tXl5sSxCsa06W6kkSkDuwWunxDKEo4tjYpeOQcAB8QAvgKy3zLJY3apF
uhMY1sCPJSmHCdH65HzDAWnQyqyeIua60LonbFja2OrX49tZZO6UzlQz7s3+ByUHpAIk33SDiHrC
TeyF+ZHp0886z9ewI+rflH+jtQLGg2wVclqA9iIoLsLAwuoV72C13lwZ6o+IRrrvCUNPqDskNBuk
j6g3yeILMBNgiZzOuHZH6DenIQM9kPPDskhGnee2Jla7t77BtLU8Xxcujqq+IXqw8/NNg3rAlWh1
aS9qJ0sz5ewDEdiUFDsJG92tF0HMJQp2DyCNEjWnTSRKVo4+lLjZLGh/s5npmDv8TA8tPkufpYEx
lzfvY3p9B4UGszuagZ4/NYiqUkH/GIKzSmgpK/900ro8Q9K5t4kZZhYo8XoCP9HMYaSCVLz6ZvhC
3cCHDbYAi5S+Qwduozk5h1nNWMSTHVXHuN3tpZJkE0vUVW8ERaJAPU2XCPGoJ1hE/m9JccweAVRE
lLQVnqxb/IvU5xNGsilYTxzmwSCVHVZPsFm5/dRP0W1QOIE5oLDvfiv/Agd7YcDHnZXZlPqGq3d/
8ksgQkyG/fSBH3HeZUjp1LVvX61Z/qy2y5w7K5S5qIxcfHkYzG0FvgTqpgBOZwXCLK8DDTtLiXre
hFvNU0M28qfWlvqKpdxOGw1/Mde6Urv099a93DcQqexkqkB5gONnoZuJh+PKcGlVVzRVlzA8AXPx
KDZKaFN5vwnmQDTvZUrW+kEAD+/LhADy6SkcLumRRtb0fbGq24xKeiSPzmO0gT42auv2MZp2U1DB
5l7bJq7UeE1K+PJyNd+/h72c5uINurh/pjvoJRF/i2neP3TS7VYkGPiQoDmV9MuSXhM+llEVRhuw
olmX7BoJXZjJiwmFUPzDEYx5ixkc/h+sq3HzFu1QHQyo56F0hz1fu8b45H8OKxqdmfv1zWcS62rb
O2Pj4mdM5Qba0P1X72eaG/PwPmV4jppmpkMAvZUrJTw/8qG6wbyAcJiSThtY6qAOb6wsTNxa9U2H
+g4e1Ot3GveayEIczwjZR8+IjmZoTAgCOAsRCr1YhynnCFk2nMk3PQRU5KFSv8z1DNl5X+h16BG9
dJUi+lXCNQld9G6nw29cZ52yFPrTvbbjyOBzvXqCyq5ns62L/9isKojm7VPbEo1a0OynZGYcvkg0
mxQYVIcVB1FJuyqc9WDe9OJ/sv4pbyTiPsGBjYt3R6kzsAaRyPZTjNYjwO5bk3UsxTJu8OQZ+3l/
/+PrC1k4nERfJQtAT7MiLaMjm9xLKgWkTkI2OfsIuvGghGMMMYZPZyGDnmbg5Wgdc5SE8KC2PBWV
hplvJCr3cdil5sI5WKuZo3Pd+Jziytaw49+JmmVjcGplU/KATqb3h9lGLzVezWBchuJfUjuXVpGY
hSBW2BaKiZD2ytVEvRdxOkNffwHghjjyXdPmi2oqDiJ5K9YBeuqubl/wL9hqT+vJNsylAySvA6W2
4U6wPKqPkPDk4Mqi79m3Du4Ft8gQH5N4yJu/vMoAQzs64Kx4AOgItalYk8QDlXTRR9Uk+IRtU6GD
vVfpKb56zcAAjTfi16L3DNk17iz0H8ImbMDXPHASwW9AiE7G3Prcu480C4jvCSRmb5IGt+4XOCWR
uxkl8fznm4jI+3LDBVvuHSfqicvc/kX/9APXJO/1GXhAotm77JTcjy33C0GolQpfnYr8v2Oij9IE
LsSAm1qpNF4zr4veGzzpu1njfg6wWxA5U8b/08CW3KNa9fenwMApC8FFY0PNK+Vmur1/Lco98QeR
HA7rEUbbrDCVQapXzmvvJMq2fx7utv2dAT99HaiLwmn60HHghXMHYBZDW/tHMx7f1jas+J9ZJqNE
n01vn0VmCuD7MlcZektqEHgzz3bFz7M9sfE5Y6ahXD1rvNUMTYQ0rHcjAAC0CU99eXpW7l/Fm/7d
jYnOwn+5mMXM2t1ZxBLXTg0j8i4lM3JSOa4eP3dFrsmSCGH+VKS+XVEh+hiobBKK+DCHy2prGsHN
PuiPT7zTp2rXsOoiOwOkReankO9N+rsct8yEf07GAFZ7JCQBanIs5D/6rIQ6uMT/DVwOcXKFfh1Y
KyGv/hsftZGNKXu3DiM9HD54NmyMlmvPIoVIk0kXnXopTyhva0CMpA1iKTkdGRXwqwerN3SKTJK8
/15fzxd4VaUw96PW+Vwuu7Z6fvChDKWhH+eREF1n+07Tab3bB7+voLB4mWNg2TkEExaHh42NUfuG
/tnQ0H5g3c/wn3A+v8dQZTC1kSMrw9SEP/epJ7Z8FLt/f2HNLBtYZXm0VkhAIoP+csnHTtEhsXsa
wknaGUBJqMgnAEFbr0bUktNAn9IsMNE5HwKVXm8FNz1sMdZRoMsNnYZkEEhSq/FgmNlS+hJ9Fboc
kO6oqLE88WS57MzrohuxRMrueSaZq9zqi5Ll5UP1ff0myOPHgdZemUQphDCdsjwjd+jA1eZ+xTHp
jD2dQLYjNwNVOiO7nnvfydFuBtheVK8R25PpXtsNaFN0sZiyb67XXj7QEH9C7RzRpIpelBKlPQKv
6XA7fwhqzjwUIlgO5I+R4k9cbtw5I8gpsEcNvmhjtAUtEqf3IejkBF2ll9dKOOG+WBcqfeKVphfV
MkO/It0CW1oDnFNSCfMNPx7Acs+4LWYLxVeq+7pEmgQbkxgr9ylqvUTJb4LZMycgavD9ck+Kxpxe
+vf/aK7Mb18fJ6g9WXJ1tz2DXlenir1Ujz1Ge1AEknDxiZKjc/FK95er8jNzjvqxOeZVkg5Mtokt
3srehHFOTlHo0qHZseLJLsR6MsfGrt4tcsiOSmYmZxMqw/d5VNQ2bhVInMwWMFEGg804Jz9Zbl9C
Pmp6ZNpAvvHU9GoftyjCeVkrMDr3zq9Fhlvt5AYmJ1y1H6OERi3MYhC5I5cekWHSFdZTLDpbRtK7
KlJAg1mhzPyDf/C8mtlswx1yyeV9dlJgDE5ycpNaJhylHcJ1z4iphU2XKhKGE+NZyuUlKQKz+Ift
lK9uh4yedDF8t+uFFN2ZoN4Jcw9CyWGyBgrTliJD4jZ7LNv7fDHpzGs6ztKF+iBC8+lC2b8m8rSk
ww7cn+TX/RbNgVr9mZMzwe3MyphcqGL0GoBTE2FwhXk38oM6obvF9FRWiNuykuO2cy3zWUEQC6He
Mb+dPVkEfLQCGxzrgl7+YsGXV/qJdCMWgJq4pDPPBYBd9+EgHNUv6qYoj73V0vh1b8L4ZF97QRwm
AmcnZn5AWBA29VAoMPLv8vK9zOwxnhNATfBUo18/5X7o2guOujKjWILfQ9Xe9GqTju4qis6l34R3
pGt3VWgkwc8e+0Bl06u/98UlyPAFl/Nqy+OWprR1yr3JIrZ63vfMBCIJjsg6wCF7eK7IidE6VEdA
mDVkjwu+Ja3zIkY+i0jktetyRDjkLJbOTen1GG3NZ4J9/QTkSZPtUnQiE8mbcXHSHtHCAn2UEe9L
jr+4Ye2yFm4jMq4M44VzW4euGKw2sVFR7cA4uSLtvL88l7aLaZInYAfcUkfLQA7x+zWn2qxUNDW2
5yF3E1KQEPWmsVgp2U4xqFzPNMrBhsBALu3Tn7oNmkhGXl/OqaAziXIQPpsdZHYoRnCMMILUaLjT
d+52CvEau6CVa/+X3QNMyfGmOz9OhOXjcSGCnN5PIlAScfsB9sllq1pww9bgnIyOkZf2hx9sJ6GI
cZChiaIk0E3NuvgIDGHfoHaxeMF+lK8bXUrqtozbVyX2xkH+GOUaO0rUnDIILU/d6zxyP4IsRPTM
SwHCfRycAC8bRXDCQ8GecI37n195lzPU4RG2UQm+XhtwmNgn+ej+0bPcAG+CtH3jvSBzJBdMcW3T
s1GsufbovNT/ICDaStqOhhipJFxxfVMcWDj0XxROggOPoNuoiHEpVcp/fB8prkCqKtazKOApcJQY
qAOOX615I9nNJBZO8P9oPPOI6v1T8hwFjTPqDaX1xVu22Um5a6nuYLU6M+sZ8whuwCyz575cW8uw
hOWVE1rQULPzP7f/BfM5Pg1t1nudxJV6t6NMHHs+mEi/8KKHgNq9AX8Ij3N0elQxn1fjw6mlj4uL
pda4pkwgTraFY6pZPDid9Wrgo3PC84qpjXK9nOywNavJQzpEmoP8exlnejECV+EGxOjc4Hznz6Rp
yJmL21i17BEepGXO2OJ1gbVemujjJN6iDSAp1J+92VkT4YmUJCZDL3daGC3g6zFOIH6LvPyURMCc
+4lNW12ROFdCaNd0Sngdb7OJkqJuw0EqXTOHIvuRxivSeKsy/Tyt//VCAjUO/Uj4fP+wHXW6XXPF
AfsX6GOwRuhN7m979DpPruIJPAt3Ed/JqEWriWa9RhSovofQ34MCBB3uBziM5msQ8SNRcpiJCT3t
947lSJtfqNVzau5zRsIqJ0otfDb8gGj9CVzPPm0OlhuKkwbxCLaEjtwpzZu2I+oy/5SVOSAjZWuc
V+PMKG8KG1n8Z44JcOly0L+LLlHOy/nSE5PBDXtHAOk2N1AKw9Cn2zVnvAu3dJ1SEy6dul0NYeMf
uzoxVuwRGHjLAbr5X+4qBvoEy4faXCWDOIueRFPAbisgv2UEvoFd2KrWa0GhE3CTpH2OUKMYVtCX
KTelcqln9O2IYYkF7aBvy7XP3y/mNT1aFVsYjv5HzblZaxpKmwOu8c/oHbiSu1Iw6j0v7fLWAn3w
sJHC/K8mRdQVSTDdWglKCJuvRj56RTL0tilPiVQswfGYy++uQzxyk0kgnCelDdoeAmNnEzZcP7hC
hUSGa8TSOIvxcv2RrnEBPU9o96JtCFf4tcardr3rJtCJWsNhKuA4rigP3exhdY8KIlSQn5SeNMj/
4pCmNdtxbYglmi2SJEELaV+Ni5JZ0ONFLVXXbmIMdaJdaV86mThdiCDRE4w3MMVAckcZh2wPnZLs
OFQzmC6BTSW2+KP1bp4P6bIaatWblu2Fxf6rLnP1siAy+jT5x6LMzrowqMiB2up43VENhh6FA12I
BBAKnpke2SkVxum8iIctHEyDwbhTH+izdhvdjpqA8KpN65DUv4iHU/xR1i2iCFSjpa/pdSqzk0Oq
GyVdNniceL9hkv+wOLgHYsmVlIzIEWyh/G89R5gCVJ/gk2bb1OX9vrjhJDJgn6Gan9NYaNHgRAYj
KYyu2vJT1oywNJT9LSqfYNjXKCMGl5IDUONJOoaOoutkwlzrOebXXTJ+dtIe2puNgcZ+x8FTexq3
sH1TVHxf491qCTIIJr0no4M3CHo/6poXHbDF5jmHyGRv4KJ08LZJDTr5YoARwuqW28R0p7KEcsXA
qoEyO/tL47KEUBTKbgJFjsphFH5Yz+RMe3RyjHVMB3HUaIfQDBghbLLHY4XHWykY43N+6iTwFUX2
YkS+CiObmeYQDjikyMP0yW+yxHzi04s81VD9VUm6v3NVV619mSXU/Q1tAkmVl8BENzVR3VOPfA7J
qz3uMpoHupC1ZVdURvT9fgrH8N+bw5klnCHPlwMFypqddeK1C/VXwumpILL1v1aN/MvSDmLFJvXC
uJ44LuGIxBEuioMS8IAF1iSYkXM96z5hqfeKz1bs8OEVNWJ9SD+LCQA0q7miAek2Iu2NuXN/J/K8
fEYRemRmIoU9JR9fwPTmfPAiyGwZguprddBi6D3ik4KdmbTtool0RwgBqb7SPrTLOb72Z1SXsFp9
F6x9khHjfy3WdwTJEPo3zpeRbvMYnDbAaf969qr1gIFFJutZhI0mmuEcDoamndAIDUU3IGYscxH9
aqk3Ip8CKVkpBCPP0WDCCPPVb58lcMHIIsDYqOkPgOcqvlycrNvc2Vx14RGdxYwnAZ9yXwwoN/bH
9DGYTka96YrFz7Ada5RNOqp+uWBnCSxi61D/Ti7kWDmz4t9ssC8BGQhBq/zCEOnZGOB4nJavskrH
q72U8ogOzu2I2y/TWFhhKT7uOw1YWUAfnGE2+2pFgZmZz8eCzaYll8VH1jlC9Co4dFG7vFBtS2Zf
9bPq2HBacKdJD73K9GSrIfdf8dnRXvwmS8VuhQkbhUS7jDzrGAFOo9bCpxz0epbwY0YTG9OdeHy1
DHXlH7LbmQoT3gi2z+cZKT1j2wENxDH8/+ZsCICHlVkl47cS1CRjbDpK/jXaBO/CngDsW6T+EZyj
b23ZFtVYbGW09ny+/HsZ7UqmrY5M+FSXqbU4sAovNELa9t4AN3MkcFgaFzFiBoX3vCvRziHsqhpd
r5hZYd40jtM2H2tXnKhPL/jjwBy8/gGtR3qSMgBB4nqcd8koXjuK5qDpLefsWn/mnvkjzzaso//L
LCfaSgiU8miByszvhUIYqpZvz+fcGQn6PcdNhnt0UfEujO4iy4jzVwrs2lbjsEi1HWFmUN/FYBFB
5p9G2pFKLuFCM8Zev3/hfrgsJgBZAan9HyEXHADU28462BsZ4P0Qu9DcuMCJ8g9SC2/D3ufkMuFR
2GEQ4kOw74JaeUt6Vf8NFeaBO8USfS9IMtC3qRFmyHdWn0p9uh5LwWk7p8iOnnMxbtJKr4HgEn26
kL3ZJq28z7iLsUocYAtaxzrHZLYQ/mrw2VePeRLpqvIUsgmTGDMwXXdiGwqkrBSIeJkncvOQ4deT
IHf/jofaAg4xp8iP1bSWd6OQbHp5QiqiFtHNwgt1BN12c+qIbozt2RoCmmqc0rtwFuN7Cc4NOFSM
Wbu4eCLtxuKM69NTa+ZGXBWBATNpXYjJjb+LHZfml6QtKjsWP3QTPv7meYF+SYn0EqNf+E+cM3Ok
gFNYTXcDF9+jCrUj4Xmrr8/JBII7ugzn6f4vUxcA3fBVR8oUyNHloDINPxV/1xlHtHKEx4yV5ais
EA3jVN9D9Ik3Ug+4+RCqMHXdNypbPtOrA174xAdEeTNO8O9f5ouuiMOTKfdtPljO8pUhG5iuRSbt
5QC2BuuHyqorixVgrptDavgbPRPWIsYfYzvLD58lSHaHjb6Ca489C+d6I7vmfqVVj9OxyEln572Y
2+IHLfkPjsTrZjwWhWhZemT2ha2E2zt9tnfebDQ2AsjxthRwE4VLs4AhWlnxUNEF3pOKLK8wRYAh
OBm50zGl1r/Yoy03Azy4Llznu15rGckYoiMHCWyj8NBpW+2l8U/WczVpXVnIz0rSrkrk0MqsyjuD
JvUWu8XQIJ6sh2mVhnPnBX31ADnUpuipdqpv4O74FbIwqXdlAMC3bxHAmE27Vqax+SQjD2VvoOQP
+kFSfFlGb/3co+JXxW2F7E3e6jn+mxn6Jvdy64lvV1PbfZ3zJPoUPQ+EuYEc3q779IG2kA2uqD8E
NE5ZJiCvfuB1Oq296uXYLZpZNyY1/o0rRY9n4z2jnnWK60l6k3GFg/ei4o6XJ2zC+QxQMd9hxGb1
FUTOl5EL/E3aEepifyTTcW9jVMoXuqjCDozEbDj3zNyoO4JAW/cLE6XRhkiQBwjCCMx+tdzsVHna
q2Y0767gli1EIHwtt7wXGyXYobbxDDkN3HJeEr6y648cJJMoWorwuhq5iaYLWCSXe20V3JaNsOQn
0DEFfzAZefuZlrUttluwb3ttpm7NqqxxcuMrMKVIrkWXHcuKb4awj5WUC/k9eanWF+I9ufFQNvxg
mXf7XJp7FCMwAOBuZa+aZywFOVD/fwXSIqkwDVWEDrF6xr4vQU4echo4k4JJT9Jj1WuOs3DKorQO
YepJCT07Uw9Hy/zhOCZwUfG/k1ROjjxSybQnksO78xllI14mza9LSlGNqsIxIE7H1meLWGAIkyq9
8e/S/p2R0jp3ZnEEZ7mMMnfMdU6WvjD461UbHDtzgnhPoXw6YXbKEaniXxlTfPaU1RXxUW9kmiPT
PV0+XmptwCBbHZLUqKL6GALJRcMy+dB7ewHnLqwZ4cUkoFuqnBnWzAq1yq7IAKn5qrNOMmNsAMpZ
XCCNldfY2+dDZ8chp4ohoU1YATJMCpZ0Vwnm4K6pBp+TZ2+AeqJ2XevNOhCqqxTEcWnOmlKUQKC1
BOGN0PLBADC3g3L/cabTmnCRZdtFK0i2DiixbgUMTAf6jRzsA+gxZTMLvYL5xMQhByeKCup+Sdpy
94YGXqW1wm7bUysXqO8/6mMdOgkC++7b6/cCD/6xYIcfNlR52hHtIwlG7nE286nVhE6WWdc6AdjG
ipL4uRTpMHr9CLQS+lxV4YjjMb1vgQjDMgU1+PDEWRK5+JU6lhMeK1z+5w744mOD6pphxusglzlc
JVFOQ4731EWV1dxjZU8k0aHjavnpzguVUvuQCyyHrtHqrOqHRMD3nza9+yX/mNsSvYTh6mHn2rAZ
4RwcDBUHahX0eOjU6V+OiuevWBLo31mHEW6JBhuOPxzg9aYEF1KaFbLThuvW0+nuhR97K0beF0xI
Wb1U3PXq9VgOZsNZPFUFsMOY/5om/qV1V4WoLKB4tdJoXdlTNKfOO4de3GWKrDUQJs4v/jPWz/MX
vLX9LNHtyCQR13K52WcfcpdB9fhvHH+SgzxRttD6FvAoBFd0PrZyTnK9yeUkj17jBkQME3uFr/z4
PW5fQQrfmm45C7DbF38Lmv+E//pVLKIMhULZGak7tp3fU6rUDkRiNDv82itPwifNkq4h+riGjxP8
iW8TbEyiDMfH055YqBv2XUuGgESb+jm5nnDKeCll/DzfDV0anqQU9r0HMGhKyIS3iMxaa8355oX7
cc2XIWlOBm+RfNX7Obs9ah/jR2PSDn2sw7QGPPLT8CAB96m+3oEVp/Dj3giNVckFFtvZLwXgOmJK
hrBgPUk01jWvw5atupwHxWk3LS4+rMoxpeQUDkfXGKJ4oXqflxDk058nKObAne+3APytceD5OJeO
CoADWmFqWcGvedYx/AosavqCh2pTkqcEawKPNyaLniHhIGgX7ZQR4/xwO/WOYf4D+h3pD9j3lBSo
CSwbd4GSuXcY6kxgWk7jI8v6DOJbfgGtHZ2ZADRGyfruVqI/X/zTC6BYIp1sEWARMCk4QwOY/GIr
rrqD5BY+6+70y6nYwomJ3PxTiUrFTJEL3LZONHMCbQRlhUUTk6IpIp7dnbg9bMhLaJQ7LLe/ixwE
08I9wE50GRxDJrPF4MF1WBUVsLVRRUUvm5HidX+TgLJLi6dn2e+we034HvNAY/oxrAolz5Mhl0+I
3NoO7Wv2d52fYXiidXHgVOk8gw2c5UpAgZewKzKtSbZ/NUn7MOA0GimN5olDD+hbjVMPnvs35PGs
P2VJ05uq7A7qbTN/i7K8y0opuRdp3OLSj0p9NZ/RDKJtdQk1jyIcxlMJldpwd5d95rK1vFvIsASy
uWc0LJREStK9cvPoeB6TFVAreiP55cvTCqXdXQbxol+olh0IKgAWMbXpdQI5W0uII2kUEwvs+x4o
4CvHGrhsVhsOU0NZMbLtlELlPDw8gBneg7zcYNrwFuUxw/1JiNq566m1Ibp5AO9HQMP13E+3xLrV
7KT/PBYxRnTYv9qZz9smv/s069OvYW3dC25gDJ0KnJIG5q6WlHerSgLezjX0/rwasrdElDwdT2Jq
ac9P8c4mqRg7klv+kzqOx0rPTdOTG5svnROWSkfN1m+QF3/J2IBJrDuL+lgOuyhw0TgTP9aX09vL
loJ7VIDsHS/OmO0XLK0HInd17rpUaeWUG2y8hQyLUke/d/a679csLE5DGJH08aMm0hLCzZh6/LRT
wXK5uHtomMS6ce/cRTEa4DXyK8tK9TvsVTGjB6otLk86uNX3K10uqKCWJMgNqtsxbzjo6OFX6uG6
H3AY6mTtE2piHLeZriegKrSR946QtQ/C0UGLOF1bS3ZwwraXBnbr3UMQpOpZaHtv5m30GKUnQjjT
Ki553hn5kBiiTskbnqT0+fBtQA6bIE7maCxe24MpbsglEg0Zj9uteEryrTlQDuy83/MYN72wrZr2
oQrRpQS6Vwis/FWKEFqJptYZ7T8MH/ICn0RSdYyb06hqf6cpPPOQ1YYHYZ+XEtZ2chEfqTzu/Wjz
9MhcVWHohy8XKHEOTwl154H1qwfEl6hmFLfXvCNa6h3PyKLngyPC6L/zgOduk4+kELhs6IvFzg5J
21XbziaF82ByVDTtVlTCSCcRg2TMHu1LlO/faLUgaQJ7BhoxZBjXYQ4M8lN5FFhkD2F6u4izzJpm
y40cXjcGevcTEDN7m1Qpo3Dhb3bguIuwHEKyyoidlbRMhYVM7yv4D0AIGEUHZAmbIX8hcyPbUOsI
SxznparKzN5yEa7ijuhWQrqlKKumuSTj/ljPNlPNeSaOBZR2LtThvKBC0DHyJIEtGyIRXoXgZtnP
nbrCIfOsPZPwLOJg9yjtBilZ0oF1YJi2SzZHlXnab7fcI3vVO0VXH5Ahx0rCHIxf9c1TspsVAzU5
SI4gdVM5TI9dZh7Nx+n28fFXO3jibW8+oGYxwkVVrfqQPbfOUELnXm+XODHuAnBGv6GUOQbEdLQ9
owKdZ2wO+VhR6fS0iG60xrm1Gbr/GpUkPo3q53qmCeT7ULVC0dG8JFdhDrLhx4XX6klIqsapOHYr
il9wtG5/oBDpZU0Di0E7o5Z/WUGm7boRKG5/SBWYFoW5KIKCWpyxVplgnJhKi55iDurrCmTpNx8W
zD+HEusSYEr+vTS1YgTzy7a8uKlJJHlugH3HjR5qukN79Sj9o29226Vo87d6bdR2Ga6EemiEvCNq
RRx3ygviooywriduh4LxBDSi2XcoZUY0aAvC+SREIDzS4FaBJuFE4Ck9L4j557DW8rGlmy0OTgw5
xc7SjyEsFVTCpZgyekqMvqv/8LbOPdd+I+VbG3wCdjWtgTZbyaMLcurgeXhKWtDJ7pIdjZ78vIpv
1BI9LfMSiQk1Lfw1kEQfRtZpWQFfwgHGrBNXUPCPeMLfoOkE/NzYQEg28G+zJDho8r+HNUhTTw7P
MCa7/ccVNLaYbbC/kEMkAlek+72Z7EH9UErYJ7tFrv7mP7zONXTMkzgkmUpNxx6mHk4LnUuuhpKq
fgqIzY5Ltx0gxcnB8BA2zLn9bccR2YqrljjdbxuXI3OhwzrazPnqYcp/uNcW0JVIbLjsTvsy+7WX
tYQ2z5HydMDWslnBDa8C4VBYAsO3k1//AxhJzGACJ/OkQw7S2uoqZDw98YfGCO4Av7R0eR2TE6Vu
o3XBC+qcLrnl0XtVsz+7W7fSOWoyhlJJLgp79Vm3OkUUonBCcTH2e9k6EQGT7Pphz2WWVc9L24YL
Vmn7sSzepbMQgqB8pK8a4sHjMFKbbGpzK28IOeZEsTa0EN4pYr5WSALFRlJGNbcF6msfo3d9vQ7A
3nAezCxpVQJaPtE4d7VRVZ1D5DSZ4EvAhennVC7qAcn4mg49VU02wuNJbzcs8jKlwAc2ftEWkPgf
LaVLL4tq7jqfbngz6y3zKGoK6xbSVUyWpKf1IaR9awqfYpDM9Qu/5TahgRVZtnlusVLgcPiAyHPC
kPIjgyfEaAk0aW5ybkouu9q8rhuMpNNpYvxzdooDK1b/O8wCCIjQAQ0bC1QGAZ9UsZaKMy2iTOfT
trhDc7pSOPq+flh5+0FIwjbLv80x6h4DVgHWISihLX3v7IEJRSpXvUshU/HAvpHHRlmxhyW7lALN
JpimapLsNhoOhgJ3kGXQDh4nkEHvmQPifFDefWrt0D2mJCWSYJdD9WDKy4Fi5+XnQiukZOHNTQCy
K7z0Soi8CfQlnwWpX6ANC6YE6sV3eU6Fx37r72H7QxvWfFsmNTgJtlFokdaGR6ww95x4LwwMOnwA
2urtjmjUnHF5kf9yfmdaTdEmxDFGEMYQZ7o2B+fTK2Junr6lDtrQyCWjmoxs7MdXF1jZNKRfrWzW
50QDT/ib6amlO3dcseXXMyWWSp4Ob0TZzLPcKu2IOCgX4v8Bcd1iSMk6arydscaK6mf9eKPFp6PA
qoSdmVZ4WeNwgoBU3x0DUll++GaQJmQ3yDdtDSPnZgTS6H8/QryUF/ndNkFpHx2m5EJ/742r9gX8
qeAxBfX6lYs29jhZWLYB3d8KfeHbJIzmZ1ZDAkljt0eEpZuVLV4Nfo0D15L6j7QuFbfG7FISPbyg
H3e0gNChhNRgF6N6nhsD1/Tl2CKb51dDsOPX0LtHWhVrN2j2UxUftcYqPpE1d6QckegYhb2nojuq
EgZJ6FY1XrKEosNyuHImdHIKpFFTrBlZNhGZTyqibzvxAz1VZ+hFKFc/d+d/KD4iTm6yBpORCllr
6ep1LlQhmowfxpvvaKUbJuCHdVY01xaEsRAlQeJ7SIEAZlvoZW5WzfJ9hXA5MpPUxvnNiLZej0Vb
deSLbenbaZ+o7U8+HMCCb4rPU56Cmq9keYQXGanPJu5guTNSarr4p9lSc+36FEm+g9Bomnfa7y5H
zm0o+W6esTD9TBp5BmIYDk2M0IaEn8Xnrdz4KE8Nn4Y86JWhLNMZxzOm5Kk5DCE5l6GXTLZwuzzx
P2M905oqif1fgwlbhLLM2hJImd6MVIMwZjw/bQG/R7MqULU9e4C9O/fNBa5ZSbeJFMTfZsB+1FqS
3SKSgrOPmZ8RCjxPKr0Wkaw/Dgyy2E0nudQIT4rKF2YK347V86BcSgYk1zDBb6nyIXChuR0l8JW1
HMSxy22VGKG1sQa3+scC0O9LNFF1PMdxuK47tSiChfd5aU2yv1KAG4OtmXg4XO8k467Z/KrEHXDS
jXYZlFgeYeFgt791ysTMA+Ua6LthHx01wANGfhfOVViYzzYHobIPjxhkGr5yZhDqFtjfGEzkVPY1
jXCVLakYnFoCPVLR6K/mglXjhPTmNaV+1/6ARnfcefaxynwIhY6iu76iMmeaEOwlXRKoTr7f/iek
mrFAR3LOvIdwalbyZnPZenMZbSWZki6b1sT4b5hbGxVQb8W6HzAW1Kjf4BIcuW6ovQd+50joXE4X
cFuasW9GiKcmw14Yp0EOD2WLi4jo8uMOyGxzGWhSH3pdMqy9GCy4bpt5jCeGg7s8SYG0Z1WAzy1O
lFDnysCEj6hgYrT75d74JXwKBg2HaD6i9m4l5Tq1HjhJXvJxvC0z83hjNNFLw93UE3Ueq1cN1Z98
6eOdFu2o15km/1UTnVNezAJsBzELnYPfRKX7QUD39O+Wc8bkaUpkZgZtydP+HhBFW+kEUVCQegBB
x8KQGqi6Z+9soY1QUDOTPbEl933xsT1Su58Mp++RBBKIvlCxrDfGx+aH9WTvzkpUjips6StEn5L1
Nm0RE56dFVVH93wBzEp3KA7gOhAzcrBRX2vJ1h+bDyVi+OPnt5Brk37e1BJ2q8rzkpGnjN0e/4x3
+Qf+w/FqKauQ6Geyhf8RnCwxuo3iDkW6EeVCm/dpl5UMpd826Un6J6E30DCiOgDssaM9qdfslANX
xfHLPv1uLx7lFVbFf4We7bUoBHAZBeIMNGIxvnfHpxylG4SxAE63CtdaQzGIbMtLUX2oULUTBwo5
R7Vk0zNylmsYTSR6kqAMEFhCOIaawNuCSWMdxjHdj49nthLaBySxJHk7JqSEX6/xAoOb58jAd5vj
Jk93PWMUr1yeBZjDOlbThevFqKRYxMzyOUzzgvVAFskc4w059ic+KavWiopI/UyB/aDjpUc24sGg
M9htB2NpVq0L4GWP8EljQcU//O5Txi/LgKgcAtzul1rhdAg5YyfEOVqgafyTEmJ4iU0y1cDlws0j
6RkM8IQLsXK5c/nn2ht6NELVJGAr78i952H5M9ybo9U7Evvbq0n1J0WaxL7+CXOt99acuNNmucM8
CKAnJ9jhm3cs3o85rW2XCQjyuCnJw+W51qtgtxldWwILvgqX86AHazFUcMuLXZLCHwgk3b5EagaN
tsELLXb6Am0+43rbGqK6AIIwzDVQFccqRooSMi81XRamQnTxKR2UCp7n/QB62obi5YtlNU6Gi00B
AnYD0NsceSj9vpmwNYZgbXeV6QDKjCpQgk/k1AMAmyaz9+Q2a6Sk+x+2zv29NJVESxVd/vi0dgrT
dCj1CDeA46iv3iwtvfLJcZXfRDNYnc0QORGN3SEC751Gbge1jZhFNAfxsGtdDQXi0xQDpumx6cZm
9tEtbXK6BUbXWMQ6j19Hcw1DpPLKvNhUi+/vqiAb+8beKSqqaU6hQxJSyN8Oal0SaNTEmBtBIcjN
IX6ZGxnt1vQaJ63imTazMofGdUbY7eJcEAXgeLD2tOqxxMGQan2X11vMMiNC+qHX/+Q03QSQ0rIZ
NJQ4T7PI2oTP4+xGo0ER0032HoZWXLJHIzMtLDRjHzY6VTMfCZQ2vhPIRqRSNTtrSEpHm5Gt4t4k
5acHVqldimfOk894LazrkcIrAkAyIn97eCcq1pF2wZTWIACG/HLzlbI5DVcwkTp0v7Ytm/LU272g
QzEZ8Dqk+IOTe35QzFy+c0+PWsEiVkMo3mkhD46DORm2O0YUhq9CakT1tAvlPPVWpRNhw4i7h+KI
emtSghKAOdOArOP4aviZFgGvLkb71sh9IF2zqwZRr/Lj8LUs/SPFN9PToZdqM9o58JAgrPqr/W7Q
a/lWSllIbPB7482ZXoH/LOn/JaOQU4wCbq2h9QqGjlBV4EQoVLUupesMDvTf0l2FAfGwaAnDLJUa
U5cAOMIn1+DB0w/eM3bTAu56QKumOgeUdSSIlmkxOio8XAvpb1UyfnsXt17Mm2F/s23uf14VcBhU
mRpE+uVA88yARv9BsIaysWbxMxmSf9Giv2lTsHiJZbX28f1GSHjBigYU6ozf1xBSrlF7+ZpZMZas
wBVlJUu8xhohnnH3RceLzA+QknQL/lBGuKCCLVlzH+P/yqC2ny6eeGNsWoHf7mxr9O5deWFSukg7
cIrAOTl+40c9t4cIEAIayd/gPmBfLdewLBrviGl2Wj1FEobGMuPZOfJo0jyaaKoYeaDow+409Bbv
jBL6E3xztTveYA9Y5QiScNDyRqBkz8YjzHX6v9ZhCaYuL/MhPt+E3srfQqldzMiFdD1hxQpnrWc0
koQZnQPtoqZTAzAZMyXlFA2mPWKSbmODBd7kAy1mooLPdntlTvqJWetg266LwXdElREPkz8pLfeq
MSWMD6qF0J2ggrYX4kFtXVjtkvT7YlX+epZIxgHHLa3dYAv1vVppur55WV5QD3PT/i80/ZKC799G
E2WgfpQ5ahR9xW8dKfeI7PkeanbQCAp75k6czkA47HmIE4xSnZlbQfIkwQ4YGtBxLNWi8QGNYXjl
UO1aO1b34lpGkQcoZubB0uTVwimT5WjcmGneZOZOH4SP+tKvbUPO4SCN9jzaON/n2lxXuK87s+8J
O7e/8ug+Hr31HvRqrUgE7vSKWhlkUUP5qLwUapJZ0xzBrgxTcxt31s6LeUecQq/BLcgNLQIOiVT3
5Et5TUFDdxmGICjufVfY4oRX1U+SHKmPr6GupRIJeYrpXMR1qkLS0gzQwqxyJ/A30SUDF7KbTMnN
WX/471oCW92L+ku+2rlOjWprohczSizQUA99RjW0DeAeC+TkaSt6mizt84rYUovAi0QxskIFqZt+
VhkB+Jj7Uq+zH+b/SuInFmCglG6EvQV/nBJHNd43jDo/e+oVMoTiyiNsNjdrJBHH+BjPM+wHDQ+l
zSg4noXY4iW1JUzZ16aguv/3RTbWhd+Z7nGcG22Ye+QbZtq7D9wD9HIGyOko4w5YE4mbJYg47UyO
Yh9aLQrB4ApPyaOb7GSry9UuT0X7KvprzJGqQ9oq3oq9xDO58jADrPg9I3wKANs0KwF55qIDHGSL
LKwnUy/AXeYU+0TLQCgkSu/cLZCj/sueh0K6rZqCoHLQxOUoNizlmBXPRCq3b5AzR8U7L2/BDCsp
ZAWhICX2zRUZ2vcKhiNU4aIdzHYvEowAOc/b9ASJ9NTYfG0dz21PBDHEIUjSZw8PTI0+2LkqKbXe
fRiNCaEr2CFinyxkhzARZVoOLmjL0NkDvfIovu21n/vkSp9bqmhTtsVojFmntl/k2Iw7whfNny0H
nansbeNh0Y6Isbi5GdACg+1l7F/nFch8I54/wvT1RJREKy0LYztg59ciRK68AFJkyQztI6uHlXPQ
HwmVp0CrbVpITlzKJkgWdQDIDFAYE2Ku5oZuq1KwtR92eTn9+HCjiB6WinjTp2GzzSAo2SuE5Yno
FQXFMeBOOc9p/BGAr9zndIWdxd/ee8cj+kVJbxQOYVZ4ix/sHW+N2/DydR3+uCnBDm6WldpO0GA7
/E7N3tIqV95UV+zIxs11Of3TJnGWaOkBxxxLl0WP/CYitebH8ri2YBTuBVt/zdJD7kki4u0UoADQ
S/LhOC2yd/mrdN91yZqx79q29lkw6KXfO28YLPFn91OlNbceRa4vkALD5nMpykTppmVmFOVDYYPT
dnLmT0UnnhiMr/QokTDFkw8ufsXYL8a9laUJXnwO3BBswGQwC7NP7dodHcjCAvgGMzfcCqBb4rCM
O79HB4OQ1vqJBSlpFSGv4Ehe8N6Ho1bsyuAh0zHPyZ+KctE1zoPZKgA61q5fvSreVqFUK4EDNqfo
1MnApizj2TKKfclenuky/kgn8oKffU89fxLqxjH/xtpsZ1ead8yfnsGv7OGNCM3RkC1mxcRc2t2k
pwTr4kIJzvP13fHpIRAwk+936OJDmqzNuFST0EzA3KUlT7AlzQLQlTynSOI5iGirKu/ehxcTpJGo
NDIhiC9JhI16xNvHK6+BbP+dQQbla5VtquRXwNdzyNMZbaQkgm6XvAyt28oTalo6B2pxjBKTSqJ8
2Ebn/uOIm36xHugOTlfC8QRKs+FPrdy/9o95xvtbk1LL17npxz1vLnjV5XfTlH0VIaXtXmE1ODsC
wo/4ly4hHj9CNHr4kNkFyDvxsBbE0cLwvGvsVH4Jm9jAWj49ndMg9wPBgESukGU5CTokApxR3CTJ
FZG6TxocFCLScActQ+NvCgEFyNCmj1KGA9QKuqrS7+3Audq5HgHmLbj/5Qh/JVqNN4MRbbf6YaOA
l5GMaKvz5j5rQmk8KGrFp+3jEM/wO6z08idAh6+EZMhQWRFp1d0iSzn+JoI7tJYy+78Y8kO0Pr1E
JLPJg1NsI+LGoW8RwmVb5iYGys3ywSdZnvE/PJ5wjBMvxjO5aqdLUo/AkpJS0ZvDqmOnVvBmzAmB
I94fZK4qyraCaO9Y3SHFwfoCvutQftIPw18n8YZm6ypQ/pcMqYieWxQYc6jFo0Mm/KDhK3n7tdQy
DDNa+sSFiQbGOIfkffiNvB/J2tRlYhfc6FGlKwNIJ832EzVElhMrmOSEW5VpTXPIRX6IUlv4EI1M
xiShlwktHCAnRtE5JvgHby52sYKeazKz4q19ZhNVvFX9vSbHprBKC3nG5Y0ysBaDM5F9yAVr0XRj
Ng1j21DKHCLy0Yq3wRAF8APuTdTgvNCattzp5KWUMyP+tTgolwSiaPZWt31cCPKjMFwUI5jtjfDD
Q0te1fyUg9iwS0GGEWih8LVj1ohMvTzPzzUvg9gzpDr24yrasqgSJ4zOr4tHoPjeCIYUli0+U8xU
v9mNM/B6xX2K0OUcaFtnoVnX4IGaAy1e4z2a/ygLh4ZyXzCAo0zJKgosN7LB3HQ/u2sngkqDCpqw
Po5asPZ4x0BatKOoc4to5psYOc4L+6iDBFGCgnMu5NydyOtJpyEwDElKp/oaXcdnqijSJBmFWCYT
Nbj0JxE8jRZ7gn6xpMCvqwkJkM5a2Gy3lNVyjOs2i+V2/Eart+r9/gdrifTTM+iQqM5/EuCX5aML
+dOMpnitbqVAbqqB+HIxrMg+CRKeRs0CR+GezwdfaziYgzjdpkUIxI4z71PbT6k/ydeSsCNHVdFu
AZes2lgGzIFoQotArq1Tlmeo0yvZ1cPo9iZCY8RQw1hS2zY3ELIKPgVj1RRHZBBhRjjQjzoexZVL
8HWvD8EfNVxUpUnZ4k9OuTZovERS3WJGUVvEguDrk7RzYogyPG/jCfDverbaVUX+nHOAdexWEMcJ
t88isXWEVH/CWO3ZalQzLTANjbBeJjxVPpMg+a+YQAFbNLnVEDkconucZZgRt3Q4tgq4Naqb8h7t
xVfSXMJoTwDBbK09FidC4Gk8XtFKJPv4HJYYPmYryIPopqIdRnjgMjvkCsGdqw/NPLR6r9iFqyCf
iVbRsbsTTXcUVbOIrsHg5FTA+n5NWTqbUpX0xnQgXkyaaK/lyOKfbtcVTxhf6a/jr4hoJHDIB0eF
17Mkz0gV/ZqHZKd2s3noMAsHe6/3sTSxDyXGNDoADU80AnsvOB2vaIylm2l3Vu4aMsoHynCzYfNl
ofw8AN1e1KPL4sN4jXEQUUQ225K1GDTssMt+SpUQvy+H98x6F6Pjgj6rksMFg5Ibxnm6z9U4VMu+
f1+2rM9xeTg/b7qtfsQYdY5WV5zC5ccJOqecBQuT09iYB0RyMf1b3OC89YOrYJgJIuXJl2D9b+1d
XljLP89JLHH63wo5lfHNWmOJuEuoppbz4U7oi4MNHvqk8MNJHTmRfk0kZxHGCHuQxk1oQKRjuOnZ
HPU2vivqbdplP4LcetNf3dOW+hD2L8bcxyJw5Tm9j22IWBlC3m1EEPkOFDWn5TCGVou/pYdnvJbT
RqxaIOe2gbeSJQVoJFftl5hflNQ68JJscVBzXQpJLvLQNlno/u3RhatzhUZm875PW1IlD7FpZETk
9ljMK/Q7ov3AR/qE4XNSLXRC+ibFpGJG6JDWw6wUCXR2UApfEKAwBf4WeZpkABu6yuutJSXieWen
uwx9lGKiKcCOTuAvT2nKgQvjGBjxgxc4pOUR1kiRdevLI9SMPQue0OFhpGFxwGX/RkrqLv11UPob
akQGFECgBc5jWSX6ec3T6W228HDvRXl0xoQFb3HMst7mrxZS3MAFCLRut+LCAqLdGQTkWTidu8HY
NrRcxs9jM6vaiFt8ODSKzTPHRj/vtKz3BGOiJmetQO1LaK1GjjmxyMdzQYl5a4OFu7LYWQl53Pzr
kwIRD7GbFLg6VGr/z6XDV3CKYVc1FxrcPZcT+w+IebZgd4s3KHuYufmWJnE9UD4E18ukEy2SlxPk
lHJNwkAmqJfRqSbR1cxMOZGe2/bt3Yk2g8eTNZzegkbah4Czz25JnoX+aHQlrw3kf+0rPYnEm+j3
IlEmG/IiMw44q6bWHOK+WNH9cJBMnj+O0uyj50NzXpPlB74n9G2dGP3qX6Y32TnpCZcg2rJvmTqN
t+n/nVaT7TJ9m4hQgDS1EYcATqrnwHGGwr0NpZkSxfkyf89lF5QXjKrX2u8LsNPZ4H5Zy7gkzxWa
roETumYlGHM4pTCM7oKz0BeqO2E1S6B28PDlPDh88MlgoM16qwhxJZ0k0D1PXbT3oYiDUREUseAv
xi8HBakqpcjQgWNj5m/OPz2AavpBZx0+SworanCp3UW11qIBMKIxN1s46MAQYrMCiOVZJGtVn9qD
2m+YilNU0+WoiEo38WkHotRRpVg/mBuSuDtjjziELESE6PbzG7IYnujMl3rh1JLbLRud1FzjFPCY
XuyEzmZFmmsAFjtc/FzmygNTo/K2cy8Pfa3/LmuroyzXq+cjyW7dsr0F7YNGlPCXkcIFGjT5qDbU
2VOf4EaPTkplxDywDSwwlZVhgUIz9KGhEL2mOg51n8c1/bUScD0r42Fzsx6odavyhdO85qFz18CC
2xO9pNJcZRwj9I7M06md/TrCtS8ZNpnlaZcoA6tLRqS7jnRpTWXg9yu8l8Vvww8ANCQSn8GLMrew
cE3R7vaBugBrss4fvL7Y3T4aTIduXwQQdtrAQu4nZxMoPUUp4SOmTZxhCuzsc2tJl05/Qy0YNTtn
xYmamgKLePhEk/KhHRUJbTbD+Sioroo3RnxnFRT4Mc81osBrQKwDIGun9yahPbGE+7paRad4sjVu
4pkchtsJnOQwLo2I7jekS/AOiOS+JiNWG30pKqk6FCkn9+4tEB7PPXtZS/dTVcbH6vmm8PXZz7EF
lTtTxKxNcMdDCF4HuTnPHazEboPFjKXQ25VkJp9XqiQNCUfk6b5tC889qDFK+Gz4Kh6EEidA5DU9
S70JZAwCJha1NrlptiUxc57aIKSCcep/Wy+la80Bo1uTaU4nfo2hxxsFOo6eHtREHkBkhUHXwrHH
/57/KjUSW1yKJDmEFZBEHUJKOzTwGvaMTjokHnQeCJru96CGGZR6viiKTLR3l/ZjmAAzJf3raLjo
tZezQxOJvWrUH75qhvPJNXH/mrGDN/eubQPiw+mUl59WfNZ2VdPS9vCOR9QAXjcRwkjo4zbKHKZJ
7UUg2CI+ugjic7U1uUhzw4teS9Xu/8HChXi/ybazyVX3nHM1O7qlm58SUNosAP5NGdgwRg8wYQsP
dTwv1PMx/ii8Ok4YByaXCxtRj4hEKNWWThmcXBHi0Z/BPW4/RQm5pDtMEv05Cy41ZtAAgZLcDqYJ
/wGSet0Nz0+XejYUfvzlZNQalnZ8bvCIxm3Y5A4m7d3ouKMSNh1EQbfAZS9aX3khYYNNVkOUcGEM
F/1OhIlUwKK3LxdQKeLj2WtlCrQ+Etphg1nDZhjqY44o1fdNgM9RKNnwdZRyoNZJfdqcaIp0J3n9
xyI8pRSSMpiZbiCBEutCwpo7bcjjUhWslWKT9qRMU9RVz84Jx5DWMYKbzO8Riruyug8aEguXDF30
4cHTzvZxUcCVriGSiIckP25k96qaqB46EjA+ShbXw8OgmWaIEv2iiqbJNvxuiOmw934t630qmAlA
GmdZcF9kX41v+ZVIvBhofms/KLZiDSGWLVqGmiCslemabtHb/YqVb82YMyqDcxY8cHCLTMpCo7UT
e+WLku7NS7QTS9Q50p9R5sL0rsiH8Vm4SoG0fWnzqovor/EF/dyL5fqDySHP66Q1t1aPjnAvqNyi
Q9Vq7KjIwMkUbFIO8SDBQmlMdU34JEC/yvibDiBuOTfDcObE6eHZ3v1UIBP3XqvW4wT6yZEYtjOT
JKAzTDehsm7qnC8yUnqsw4sLd4BftUp+gLncL7VwpG4HsN3pQqXoIe3n1gRPKkQIESVJWFypcB6w
gDufhy9IHwcCprC3tUrSg4/yn1TbhVAKQUWBQU5RHn42+/jRvse2n/ChaYRH9qyWsasScUAtu20V
B8U5DlSBwLfLPVkLG2d06IcOBA2APFew2L5vyrBz6ed4lrAnsXQFCvMQ7MlP60FXqE21+tchPCAq
zElAlmbxOhVm3nzXjDhmjWixcbguPrB4zDr5bKjG0ya1ZpWDfjmBagsp97gDU71Y/VVrEh1Zm1OC
uJD6CvlamEKd3QjAiSLzMY85pX5OV1bM85MeU7mWhN3xY3GivTQ5ISlCoPSwovT73ia6fJTdjPtM
7pAap02fiHazuBwx18ec63bu0Xtj7ZNyh3Nd521eicnyV3fTrFC1rOY1HWiRh1/m9LnavGX1MNUv
/0B/SzlEA+D91Hlx+D47f/1SP9uc4wVMvB0ekQrDoN6vd74I/4/q9xYuCb9aoWsrIotw13lhSQDa
U7o6TVNFBMDzgoMx7rqajVwtVVVDlXYCGE4tVjyHclN7evt6LSgFtgtJvc/++ZT0xRQV/f3y6hW9
nlY6y/BIJgfLfLCggK97/8RictdJnI3qXfDFrFn4mp3CZu4aidWCwbGYyxRv2uujT31oFb35XS+c
1h9Vmq6XVbIa21n3WXuqIhb9oZBl7DwBqyWZ4uoJdgy0zKJyv93PZRdlfk/V1JwxV+/pNXIy6QM8
U2V8Z5weJh/wYaj2Qqldmzcnb5nPbvA4oheUnzWM7qXA6Pok9fHK6z2f3pgMEH6oFI+J2xoAHqks
PlCMfAGKEk1UMkXE8diD9qAixmwizcx1yTTNkr4x+FjdYMOCT2w3uajXcT85nS7bBxv8JPh9nfat
ZVdI+X1+35Nj/Xh1iZmgUUc8AIwTtQiLEL/K7PVPoG8OVTgzcoRG7KYgZQ4Nhr/CjnX1tYQlxpn+
ETTyGVDe/b2w0x94K1UmsQ3QIyZn5hkBxo3HZK12hh5R/YIRvM29IP9WA9AGd0+dNz4INBz2lXN6
f2hij6PfeLMRwpogBPcB8xDCBut6GsO1bCJRxsH+LaTOf+j453/GvKUGmXLAKSDANZk25iql6DuC
FIaHruhllLymEKRYGMEbdqhNGq3YbJOeKhI+1Tfwb6jymsUrfDBaZJlbiuwFmVam5/tMQselTmFR
Jjy9Qch0kCeTKSTenwDlH5XwsfjRkrKLhGJfIv+oqYfCwjZufknZnXfUj69siUrtPqgwwd9ezFEx
iG4T/ZndVELZLWTxuqr5BzY9cSF0hoDNmQ+znuuqUxvyAv6lJK9bbCdHDMyfMy9VNcHMvNgdTeon
Jr664Rvge65FZyFNbas3l33NdIcnlk5jyot9YhGaX6Xh+J+wBOjHRlEOw4bNtstTrVE6CD1t/RgY
HyB26fJQQg/HKopA5ASgBj9i1dUDv5M2rN8QvPBlgilHhJHzFBZHIQRcKOUI7gPkp8ZwmXcR1YPK
QudJJtc/xRuKXYqks831qnMg7F2k7H880WEQlwegqLq1KFVjo3EmUL1IwXmlTMihyAKnOVGcVUNg
b6BiucnMvdlUahOaYjqaJPl7Z/C7ilkGCPehprn1AiMpiYpVVIFjkByp04lb7ST5Vws0pMth2ags
x75bRSNWB5tAr/eUJka25iaPpO9ppkCdBdzRn1dWfmIVWn1u9Pp4v1UV+qTUEDfPxjsqLP9Vv1ZR
bcqfvg/twxr6KVp6+fviYizRPqtudMzoW+CHovh8HVaKfQHNmlgjsxGgFu9fgeHPQNzbpDDGjoAv
MiIrKzwKqMTXwa05iLZTRKoM5kUa12P6X6fvJO5ThooT9jr4tSp/Byl58DKjyAM3A1hXG9aPQ2Ym
moxMw9QfbBiKR/VQ+HKl93rGV8S7b769KNeKu+/Mw7gmkzwHIC3lyCIOdiDdsBrpZAQMjoWGoPQ9
p2dGFSdVt/WYOn3vzw78BcowYjh7gC1bBA2jsSLI2MND+p/D/XMl2ahE6RpNIH2C9HMqo3+ZL5U1
JTL833CvVYM7w/JeGLzCPE/YmqhIjKH0ezW21DP00agoUmbP4k8TiY/zO4Vyrejrgf8hrgPUc/et
f7IJI1o6zwZsRNleScZJzYd1cCq4M36CkrWqnVCrJ6FHe8XAICqaUXErsOIgr16bElypYkyA7r1y
9pMnBm9pkyFfcD6ni0GJHAYOdR7s7OLkaFtMTAAo5eDJiWliN3CxxjeBW/cdKlPM3N/zoPZfA3tq
SKVISplMw4lvTdiuwMYWgNvqExL7fOtIWs6aasan2cRi1TMOuo+dxUaAINfFS7Q0556arw/H/pc0
nONIQ2wBncqGzUxpnkLyfHtNVgEAuNoImdQJzdpSumMnk3gDlleIvOgzJ9nEQwZXMp423Q2gzhRN
B2i6M+sp5zOJ9A4K5HSrLLXPq9C8v76v8iF2VFokSXyBBZqrCxLT0cucrHU0ghA7C+ePuKfguHsU
w5IzRh1VBvT/Kytz2EvWZRVvrhpYTzGbWFs65CdzZzcJn7tJ23jT8c2axkHpOCwsqJyS7RnvN6MO
s/LTTV80RwbcB4WuoXfbegmCDvFUWuyKwW0hd69crshrAcaqUwhPFzGemTHsx4qw6UT5wwQQQnEq
/G4suFLzzzDISwD1120e78lrzh3kpogIaXDq7duIVL6fE0YzH6cyclIkmfgqG5OAN/H2jbXAnNHg
vHHIOFGVat/yEmcDNUcMMyWl4HDLxZUwpnhtwxxbYGlMN7pjU6g3yJUB9n4wXxOuN/YHg/BGCM5R
EQ57df0Cl6jxinAhlCRGKsPdXVjcVAzNiHMQKR2lOSF6JFHUuR5mtUn52BSZXPb2cYFQmJzj6uji
lilCjJonb70LteUuvpuau3UZIeR/eFTfdjkw4qRSQeLX4orrP2KIVeMuZ7IC7qXZI7SyhXKQcPT3
KQDbs47Ewa3Ny0x56WT3klm+AcWxlvMZ+d8B1IS2YBIh4o/34W5YP0Gn/68mpGmFQyOm61NC7W4S
gqRH0uinhSTp1VcvucLvD8xifTa7Huw0s8kzgoOmmr6n2Ba5xYbxsFewofFiz2/gUQtEHHn+vMB6
148e+U3fIzrHRYvNJsrQ8S+tFah4vTe7Cj2TznozbkgL7ENZTf53GYObPuUjv822Hk8pH26xM5Oe
RomGGsKl1NBVl3QGbk7QFYpNigxePqWhO2vmYVTmCMTcffQvkdmB7p8CaQnmCk8799t+xgN+xgRq
7j3XjIp+tpc+yDRIeki8y/Nq/uGmwsafM6r4HlrKE6XjKUgkAxhWqcjtfhwx8zKXpRodksd9zkE1
Sx1zQtT2oc8EwtVlQTJTxP7KAwNB8yIBRcyhljsX1K9JyKpNhZhE1ybhMMb1iJdUph/RirVSkLkI
n1Yxwt2/MjtzjAcgjTsnuxwv7MHpTI6xsM9KGhDftb64QjyyR+o1wzRqY3tQmsKI+9DeZbrX0kzH
EVWEaqoqjSynPxSiklL0O6jSSV7MJVpgiv3zKu6pgKCEzjbAnEDns7YqfPfT0HW/7On4yiespgTl
eWG5+LOmaae+1NiTrtq4Sxj9tfwEan3Qnj3nlIs1T0bid4bjBtG6hnvWHRLRmBHThZHJLka9V5MW
WY5Z9rV4pGMDJePcLkSugMqpLc5A7dYxMyr9ES3NBZw8ooT+IpGva1UxnhS47yLdQUeYeUFtdKJ+
pdOl9wQtRbyM5nHTIL3EjV/v9sL7FnFft46ouGKtfKwWLovrkX38lNSyzdTjZTH+L3gx4kwcCSka
b+uyWTe0LoC3kwBopjGyoDt7SIgX6j33XKhpphOsUMP32a1foee0+ahTKee13EWp10nAlHiv38d9
skadUl6YkG5yGomakaL90JlgYaZbWnzLhwD06d0G2DVvpdUV52STk2qa9L+A6D4+BUNR6CL29/gx
GKOUTd0lTNJAzppWo9hI/LXF60Rqvekq/lITX2swjjlBtXy2U0mS+ye2xFhbOF8R2TadpaTWoRvT
BGNxYfMbvgAqi3dKo6C3QaYeHc+sO2axd/q8/SUTxikeFZMa9ku7wlj9XuiIQHwOCVOGYQU5IjyM
dijDy9Thauqy6fXKLYEkCOLN/D+0UdyKUyMIh1HkgRzBL4dBkCjSnzwv2mk0/1BAxa41O/N+DVU4
jFJx0FyYN9IqqWArCZIAU3ptPUiVQuEH01UoVsjbWV3cHSPuWItJKMeYihHljHsb8OAgEZ0KWSP3
UeiAbI9V74UsFLRWYaEdCqb216ek+GPaU9Qqhtb2fanYodiSo/rcUxjTFT5E+mhc0W6b/a/K9W1F
Tx0X5jpZ4I6sPxcL8wJdQqfbefJmmCVUgigcDrwtczj8yDUTqXGfb5+krg5RQkhP8856FagfVQce
rHVepxS71VNWUufLyZdqSFfbgzHLrNcWipl7NsFPCfrDwSTiAOD5XVBWRFf7ladO8tvXg8ZdqPyK
lknNRwXHJiODnkcQAvk0LmSAci1LzLFLdF5GzvrZhgZnqpw5KKNV586HPMjE5aZW6VieRhCvNBAj
GsmSiDPRGs/EjcCP6lHTsxUjLGBTcaX9FK2ahW8f5eM90LgY5INjUuwPmBqE4PlVRP9zbzHoGv5v
+sti3beEDY21GWnRLeK0e8Vkv7gcUJHNAPmN2MiDjQqc0Jmg/0r9uixEkifHoLh0Iunp84er4LC/
aK/snMamBKjQe7Qk4sK3f1shXmILJvsWjpv6YJLh0WNck2QOf9G2uFCJQ4HLyHveND59+bUi/0kM
bqDPDoTEXkj8NM9gV00dCCgfN1Mgobbea37fcxdKEag82xyHKxfkzmzCCI2ax7qPlSuTDJFJcsPl
AVLGOZs09WAlkvd6xmcxFyCIMypZRpE+6IU0JJ7Lj2f2he/jKVvAQKPvC++1DU18NymloVAhXpvt
Vnx43x7Me+5pcdwfUOvgb6b24pZ+UrtBu3AEEORyOfMJJUjCRd++VcU+jGdx23nBYN8AoWJqgBkZ
/Ne043+1PITryy5r2yv8cMDywx5eoMVFSPea6ELBzPuTiuZbTg82vTLeSqX/Vavuca2J0f0czmqB
JdKR5Lwv5Ve9qpOszpcO0PX2tAQdKQiIeydTbUAivbSu+4ooq0XjTJNiMBgmfCYj70OYAcdFaq9g
/D8D+EoWvyYIfuU0cXCkP7cJ7GWDrHMB1Al7CmTr1VS2ovu2d/iDWSBnhZAHdmlF2y6sNYfOCKno
ISd79zU1zaz30ci++gsaOWN0rVMmQ/vYaunuZhjBl4AQbzQsYZ4ddH257dZPBhupOww9rVkon91n
WK+Pnu75Zr2iSdqXgyXh7Oc/WGuCbVJSb2wAnS2ARKbMKnEor2Aa4KYXjucFoYtl4Vfy749qFUfl
1eAV3vYcGTVHAM7SjJVnCHVEQFF980L7CiUZSFtBxV7Nl3pqPIram7DFRL0ID7WG+2HE2VqPJ9kZ
GZv98QQb/+UxLp1hs0DUoSEorGbeo9CsaryLEAUi8vB4nDrobm6zcPcoXVGOyJOfna8D43kwbK3/
9yH8S+0N4lO/xvmuaYayh3VErcI4B+zl/FPMvtPSqXGds1bBjdzIhxLpffIM5Iu3SPCGELArCcse
oJBiwMuy/AhpatV6KgMUTL4384PNngX0KQhaf2ja+Dow5AFaE7+jVqRhit9fKmVE5EhBNETMb0J0
2UuX+72aBgv/et0j4TpF8g0+GnV1tSoCBG5I925ZAX2DtcfDWdP5DuTPzhQzPbxG2K/G/QHwrwAd
4KPL0ftGPPHbdEBVAov5TKPafb32nc04Va2Xy6+bIId5BOCiXXfiODobdVlfeuw8T2fORdISiqfX
qnA9KeNJ1Z/Jj5HpCR69qzxKKPWlumTgMOCyzH6wWvUzCnD6o1aUluPF+/k2twqaFfnqCoJWte0Y
NKtjryhKjIKloQMtdWLoi5XU8B7y9Yd5vRyDFTDHcAJrB0sTGpDfgGw0p0ZX5kRA2uj0QywaELqy
/bbl1Exv6fyngNi3h7cs6KAYY50qrDXMjkEAro6D9xbKc+nk3nkIEZrIWiBQGir6SSRpqUf/DIKW
fbPfxYz1/30wHvBueevqya9mcH36SMA2tSR6hfqZ4k8UQFYvoJViez5Ik37cKTuvx9YsaMgX4j3s
14ldrHT5Ya9j4EcAexwDQ+scBqL7mfusMCEPtaEuYHrhX8PbOfepTvgyxDI76ILcfnyU0qmfsomH
bjdMmMJfMKgqlpnIv3e7+/LSC6i06CGctGKV6NWU0n3SUztn4jJIGGUuNqY4EEOqIa5TM5auLJ8e
VPjADpKob9aYJHPhlPHxrfWK6iC+v1FTmgyZyWStn2chJAvNxkbcVYHVQ+Ii3f8qOFPZguKfX/P4
sQccBCC02jQNQZkA8H3jZR7zkyitoDNzJOZvT/eN1Z3hfLpXbwFsuqsBdNpotoJLnqarin03ehUu
PQlwiDDd0w0AosxT+jfCyg1zq/KWEgDJ4l+BAZyq4MDEFlpCXzi629AVByocKkdxnHdKKeY4Oy37
b9FWgFmjXRMWKF38UoMN2ZRkyvmwEHnGsuHSWcnAoCEpGpBQkE6xJumx50wJRRY/6ADTvK+9Nwa+
VJpDXPNX2xOzEDB6hLp9W9ptJ4eSKWk8EwlmaaXlUXfbt4P0HuBDYbCNLMq0BDJ9Sdyou/dV+xLr
+yiw3iG1pmDO21xOxTPvoEZMarIaApfbebDV940yG6l9czkU6aiJdxamYIq2bXaRboLy2kWQbdCh
XvISSSvg5ArVmUIAjm7J6WaFT5YVoerQyThC6E+Am7XiinuzalWMiI1KxqQMnqOnJNaxmWV9LWcJ
lh2b/XpQBvm/d9HWHFOsNepGf+Fcx6KWeVWiOQFGTdFZED1Vqo6KOgd4oGME1keoFKr/OY9DkBuK
npaMtdD+VFbraRev1pzDjKo2bBEZjzIko2GMXKnEtbaenMfRMnrbiMD3VO+X8CShxuze41Z3lSId
OPna7lEeuXp5HkAihEfyJy1wPPio4GJspyZNPR+16iGkzGa0YkfOK63jCZr5xIiRxmdnt1d1PTYY
E5DNA7tfvT/wL424fI4vWF/ei7ZT5TG4hRyWs3slWttM4WnaNO3YYHF4uAWatsb0L7SzrGpdIN2B
YAtyIbLzGaSc7giYKB9ij1SRdpgzV+QEmNw3w6Qk936ShqcU0lUsri8mH2f9xpFbI4Mibcqjg8JU
G0SPGyK1r3cO0wopR4ogsNX2E5phMqqqv4iBCNURLYibbkU7TEHRMOUw4/KfaeLTCQ2qddSWLZJ3
F8QI+5dugj7j5sYIPJpNjiPQPoDzv1rd5RVg7Ok1hK9hrtSzPVtV3ORJQUFIiBeqn2CJlAKClOsL
IImcpq4nyRqQ9t1Q+QmVFBzXdxTo5iG0xRgmbvvo5SaKqzIcXOn1BVaXJ8NfkMKoSYJPpH7EpmbE
TciUxFmoJvYWrRSJ8a2bJXAHKhNaoEise+Kpb1XZvQ9e+JtVTnnA3b3tsCCgssD+LStGEJXjtHyU
s2sbSs2jBn0UysxY1MpGO29U4IwXCdZZNEcJNgJgXvIubaFw/Wfqto7x4XybJWqhkQ17038WDlxR
jZG4e8V5NICuwhVZXo+q5WZHO+X7I6JVW4HsOs1F4IGFkd2IA43NjLOple4hc3pNrmq9lw3yyWf6
aqD5eqJE2L/ptilPNSsZMNeXU2+Ve1MU20DZ2BKyj6yKo80x+//6BqnI3q71+qTCQZOBB9iE4gQW
3n1XAOS3qPY0VdFVbLTgiyCi7E9xQg3ikgJ7JMoF2BAowN23gxZI30zG9Xjvnd5yg/PVdQZ9Umh3
rYtf9luHItOZBl8C2mrBCDK1AaRMCCBowyTJeRue5Oi+Me1kmr3sOJcE2CartfmrFNQFGX7jajQD
JQstbbirkdB27xFW/zWbMMMaOO1xUomB77ri5phvKT5IdrBiet3AVSxZDimjrFK1nAyRzQAIvYW1
5kXgM5SWp1DDH+Geudi5Obyouq+gy5snrAsRZ7v/fMbXRR9hFZz3MUvQ1zaYQqDlaIyjJC3reDI9
rPD71u+GpJD6WN+x/7FYei7QNEcvT/Si+V/bQiPd2pdbX6oul2sDqKYv2q9wZ/rJw1a7OtxkRAPp
NMiq9gFVVyE9hvlxJCZz8GV4uVAmeUokZykLuLiqihqMe/WAlyaiTnw0WBUh6mZudFzzKywPtRfp
XHOji/vezLmVq0tvX44+EYGGlKFZplSFdDBq1xeFxLthuauooB0R4X47SgIyJlHMJFb+THLNo5l7
3LC5nst+2Ld3ZSYEeJG4/3ivb6lqDk2nMkjtTiCdjNHAu/5fp4ujC7bEke/tN3vhvtEZJJ+tZ3h0
uXkAwiHiDm6x7E4M1B5C5Mbjhya5n8+Yc6Ow07Gn7jqMz4KA3OE2VnRHOjctLDK0BqOabHCNTPD1
ZD8ZBSnbeeKtYK/vJo9hZgBKqWhISu6YSWvW3ns9rcrz1FzlsomqPc0aU9nJ3VoEthpeDFPKU6A3
6ruHRsBgA/oxJr+3gYpQT28FXNedakzc8aSYYGTOi/JBAM7+ziSn4nhDA+0TQHPrutqJsmxuC+PO
97FyMl6276X4zxhmtBo28LUB73j0X6sPpasTnUtbx7FNsjvKvBQ61b0p/KA0GjNvTSfukUndBaNd
DPVOHGY3PcoxQMl4l/KNc8cA0Bhs9Oyh0H5OAEgPJkvPxqXAhaiMMnZoqxKQ3YcJI4/U1bi1Jqjc
CYaqS71VaL4zgm8MaLZyArB85znJhU9wGnic06CwTuunhDSYDdAyyxnwSUMsjy8LeyPbPHYNQ7Sj
A9O1Ap09orM4O6Xed+WqAKYgREWCBxIHkqaCD6PniZMQCMu6lsLoKyjNb6dRHr4EQ4mIhOClcM5q
EpvYpJlcpFTC1Cb7+i4WB7Kpw8D5xoKhq1jupa6Q4zUF1u98UT6FSR5HrUYGVo09SVVSzNpWsxbM
8CWWLNPx9qOkZZoHJOoKrpdPNXZ1VHNfQi2P9bdxDKZQ9YT9fkFnGuSlYUX74GOujMemIQ/rNz6V
d/F1SDeZ9MCdbpYyIjqX3bnEL5ze8WgHfxZncW4A3FCHoSuEIhZ9KdAuHFZH6UWTb3pmNvPRdxw0
UgYTBE7uY+m+6X7Pj4TnpcirIO4jvYNo6OsZYWD86StycVNOljdwavhtzNu4omAMZzd/Ykcswp+J
YUuPbE7xscqWMdpes9yqbMmtkhcjWcgfSMgSVqWVmC8uHjDXFfumQUEPjqrrfFRJvAWxWUoldyiU
GE9UdzPZoFx+inOLfVKBSGnDVGZdTpJBiYE+EBde3Y/Ippl/DPQA28CmrvLfBjq9UsMX6ok4GOqk
o7PHD8EYgYndus/YbrvJdNutW7PjTaylUuSSSR+liNi9XSNcGx7+f5tywZZ5Q+SscJRdS365RCb3
PCUlFP7e+GdTc5cL0KtblbLMj44bJNlSHq7UJaKOg4FTiHxVQV0ArlZObWJyAumxHESgFQXH9xCm
2EucACEcTumj6QhNh0gGXB7UP9soB45ceV3/p4XO7T1kTjH1SyKclY2fQokGFg/+dk5uJO/bZCO4
8+ArcYJcMsY6sbKVUtsX+wLFNn0hM03F+rcC3ILR3Wzh+C81ts3btpMJe3dyEVMXcyYbFwEdpLke
7eCBXy4oalNKu3aYRPXOLd8CguxMB7FEwTfAcWCL4OwYoCVdt1+IFRtlSjUCh4AltV/EDHUUbkk5
/XiQVTErBO0mo+MMUTZO3OtS9kkoF2BCElY+OpKvL/z+fYo1t30h2LN0UeMXJN3OkrhqrAvJt1EN
bmnUqzJzpnoeRkjIg+JkBD6FlRgYoMLoxqbJOM9yMygpEM8ba5STgWH8u1GH+6DWVuR4yxNuMD4g
sZ8Ql/BZcAhKRTxXGXRoylzB0fgNefwto0TqG5en6Pb70nqZs+5tEl433qU7XKcfQMUojFYpeOiW
L58tAe3l+s8aLvK0VgJW/bYtFxgMUVN/2d/BmpLPd51uGYmcUgInVGrlYMGcUlFXx1WFglzFb/uU
t58VdwgLZVtxA1O1ClX0pEjNJJ/E0fuemyhWanOjw9JJz5GXqUvFsRsoWbFqjOYnD5q5ya5FIB89
E2HPdRT5fiI1SwGhYLo0W9oTYjT5lw6DJHSBeGF9l9p9yAdXSqIEep1kj9RidswRsr7g1doIj6Ql
/tBRm/TGT+gcfHOmFD0sxVACvp4lqSsiy7cYKxEUqcJUUjO5wonFwwTIFbx2Oh7EOyAtcUkuRiP3
AqWPI6T3WdZcMHBYjuSwlxMaBxTXkGkPpUaG+7+E0vgpUrCJzGn0Adcmvyn4YuSOQKZeu1PrAVf8
MxHpvGwK6tbmTRTH8ySoFxCyQyAE0vnQQ+2xXJIYWUKoDibKaU2r2lDk1axwfnTj1Pe4R0unpDus
m7iX36j9nc1cQfP2LlpunMDIgx1Yd8mpStbAkf+XB41uEze990SS9HWpT1KC9CWtHBColeppd/Y0
8i9H8rCATPKfYF6nxCL4WJgZP1ocvH0/VsVd9p1Om24D9NoEQV48XCmaqut2PI+wtGGKqnPXcJ44
chOwSsAWVbTc0zyalPheOwpyYS+EmgrE4kjohQe8ruT58gs5yVy9UBuxVrxPY+5UX438M1QBuITa
4hQhw3sD0UTYetQqwEc1Gy5ykr72MhcynlJQloNBAqhW2cpqgNUot2l3cYuvdRyBAGa5fvV2/kZo
iRxBgCVqEg6EwW2meZiTHM+5lN+K4BuSqCJRdXJ01tQBzwaeoOGNTqhZ0R+SPcokIn7cmWEV6uGQ
UeJpW/x+wxx0BqAazGz6l8m/MsjhlOhsoeSX8OY1aFfkxsaWXxVIRhV9+CNlxnf9Aal1k6dH7MP3
+yIeTlDsMZ4PqjcCPGj500tgxoH+OsMDxcuKA7SPxueiXJ92ZwLoNN8lpdcOuxxOJkmAfU2TvN7r
SUhIrOUmckLVqzJLbd5J36Jchbj5xccWK4OboQQFjCL4UGrP87yAVtzHpmfz7/iOXeBEszraT8mv
Duocz3Fyb4jiz3g+G3h+CfE4j1xot9yiCotJROYcuJ51WxgUuhu+u1gMvAiTyRIG7TEukoCNjap9
jUwfLZnZaQMDpoBADGu66bTDWrLfUuWH0qwFw6OPZENzm/K2P+IkAgnWW1gpMyiAahvCVpyBLsW2
3q6DrIf62Y3g2QqNo3pyXUWzCLqi3QTdcq3Nsejyq8d1ETPCOJop+d3WPXZvNDpTIyDDGzWWaWHN
qKp4pZx2pY2JwWvav6t2DjpYTUdjbwNV5SbZp814haZnAgvSMScL98ZdfecIUWXgYw001LIh4x6H
+7GBOcx/wsGJ+WAu0jdk4EUfQeHyxX7BV5fcJs9oivoZ+S3e8oAptiNP3rc9PpXCtypFU5YaEZex
miv2Pb0qJNNARGo2h5EUkesj6avdHlpghlob12x/0YnrS4J8SLAHDqlJ3Uai7KTDkYJQQqjhHd+Z
9Nl0tkVAA7JE50LMoaFwR2sPoQ1HWpNUqNCBDk9tgbpSosy3ZtLs9EaXy/I27Cvnpmuze3ulx03F
o91fs6OxrNyIOupKcDQwDAWkknHTAqZL24jVeX/CJji3EPQvxaNhEVLtNO7XwMC/Zknt6PjP/13a
BvjHtssu+VcUTiJwN5waz4h0esX7YKCsefZ0TwDvOoSKk25dvZM+/pJ1tMxP+GIVWrsNpgGgGLUB
a3y2wQrpKHR4Ev7ToAFF/J08UIQXJGz+RmWDsg9jp1ML9tVn0vEac9PM/fcpoEupLp5R7EdNHhkU
4PwVIjwwUolhwbVq2Or6Y7EJPmqYzTozUja6hy+iy/uj1Dq9fg/2VOqTX3LSViMudy3Q3sswf315
g6sKjeP/mZWtDo++Sg8ayvqo5nWd7Q3pELGg+ofbr2ppHSuB+cMwugfHdPPjAGMBIucGRxfMI8iy
3RaBgdZ6w84U4oyN085J0qJ/ow6QuTrJQI0Q7gYf/14G3EIUhf8Q+oQhrCklzX9bcUrnDlfLdAHx
b+v9849otjizwlRzASfaVWX/QqZT6E4emnRS2sMihCHOI18tOm1MHIXv891aGCMLZmsErey/jiJu
bvSj5I24Cp1CYgriUb08iySbTIS8dXPLFsEojXlNmH194SviqiMko8NaRddxyVErhbtOsndSp6Zt
0UHBsCFT96ntJ4eDYgEUhVrNYdcJ6yLGGPyneStpLgZQ1Wsf6APnwCCurcJwS4njO/ZnRayPhJ/3
ZW7c6VykZ+a/jjcvX3hoRindRdY6s0HA7mS3DWyNLbacHVFFzaoJLQ65jtaRshD1ml2aDK/CnixM
w7XJhNRf5oCgHVYTf4PU8qOFl9bLgXYwa/0X1A4w5SZhnEo4nEQx37yU1ecsnZnATGqiSr35mMn/
c36xVAS6eZj4UeFwfBfVwUOYDZURT4LRW4EB+Ar2fvmHDDl3UZO3rzr6eXrk/iwdUAQT3c1LO4E1
ESY5HCOAokSbZFP+uuUNX9zHIQjWD4BuELBvEapVHA0/98xGlFMvPxs6Rg74PdYcgA9hm69g4Z2h
93r9soz61w0ka2OrxcvHn6Xl+EUO99cYo8jOJt5Jg8QblZMcECRvhmqw1oRJbFzbLFpOEXBZpGr+
gnluKPlQiDJYQFMX/cGe9T7yaX9JNRx42r3BUsXHKMlVM8pa6HO7HF/PyPmcxNIkuu3T/WvpvkJz
2d1Lv9a5sRom4qKAlCoh8wCa0uWwvac86KUF7VJxKPjsaKhxOsRRGXenF3P/a370KJMcQGUyV78t
z2yDSPOxExFeZ2cgimSKPzJzsBh1XoGpQj8ggv4Jx3BED8T5bcEczasuvzgcgv1fnaqejk6uAE7w
HMXW1GpnCWVu4nJO3vnHNNYlAKzV7hzwQyZHV9r5qI32StrterD1qNxujfOqiZ7PDNGTOKC/STqx
oNVp8HqYoyFdhEsgorSxaA6az5t9DxYOCdQ+EnjdLzdwoCfBDR2Git6S0ZSc6rgxda00iKnFriBA
IMhaG1iXd1hIdW0jFYZGaWgs8PuZ9xVyKuuFFxWK19IJvsU4OT8I5fnOAi/It36ES+kcgBedZbQK
0QzpFWqzdu5mwBUJ3hN88QA4s9sdeN+U/jZ6CdU4eLY1O/D1G1IMOqOA0bUehZtCKsyX2f+Vwa1X
+OPX5m2GXXoCd/E7+3ShpYhfdsAXLjuSG142o1jSCpwel7X3uD3dO3TY9NdfcdJfqzxZm0/w/Kpw
nxJniNzL6reaVgyGW/wgaGwegSfLwr8SlSRkgglOBEixeTTcgYOxK7OAFGYqM9ZRSBHvjiVy3hQU
yfent9Opin0Qqh/JjlYsTGkzQ4hsDuaF3nPLXBVrwct8113Dxo4pfStO8EjaM7wZjIl0X7viXcJ+
bXXL25UfDdGcCE+IBsB3RxppL+FR6jtTl66IpeRTCEgymPLA6JDD5bjP7Lh6L+ibLdjaE4B6Q0I9
6EC1ihXJDAbwabkDHBZ64mbvRxkjkHVp8/j6Zz+onk9gIKXxEDdIGh7Ci5GX0yy7MoMkK6I+kOS3
vdU5dZUudullYm1B6zay+xST0HlmSSB390RESOUPUkiIChXiJKPVDeCN2IUhbWkjI02/DtdpmIqO
UVFMMA2/B8K8YbBOWLOJ39LGMErVPrBKri2UpbBSZVh16GkjpSCAK4nA7mU1zqolhAXRre8eTCcl
nnlUsBwWTpSHdx3TAlF+wYY48eYRObHR001t2PslrqCwvf/kt6okogOVrqs7JIZwovB7OcRwXb6H
7lpf1FOs7TrrXE97tf7/gi7J2GAyCGywwvo3LWrng+MikMiKbIzq8V3ggUh38+aVKNyZZwwUM2I8
min0NlBVVluH4terwlbWq4CJQ/+k4jXEQVBTP4i3zN7Tv3DwEjutTm69bWRlXYybifrxp+8upb//
P7b6exB4RD+3nV8WRrUWVKDR1HaROcmZVaBeh0RV3hX6VFqxgVnvQPot8psEWvvQPJBwUBjrCStl
N2Lsp7rNPkfJ06Dpb2uI+R92Dkg22+M6J3mKmNcTeAuLq8oDZJctouOzY74Ilf5OeAUG7lyhMHyr
IiVyw4LiI/O/GDEFvLIYLBunminhHEJNI9bRK0LUZQi/fsJNMRmU1hb/QG5//MmKmMqZ8NNLJktw
B7/aAnSB/tFtWs5aUpUE9ocsDC9+lFoQ8aKIH0T3RSoEqjaUHP0YrzJFcTb5NK63vvMXDL1Ikx8Y
c7IQUjAgaXPAuVspeYiGvOl3eiDxgkzAAi7sPIMaF+VHM0Z6vOFaNvez3zxfKV5VW1sp4oS5gUh8
kP32lz6mvQXTR/JYzkhg4LiZh5DPxI5yjmkMAESxT6JpRH50y6QKPlq83CFL55VRmAJ0MXYb8Jos
7NDPAf+YSUHGS+PWqRQMI3Fb+wM/vwl8K9b4iXJWdbAAqCoKMYgish9IYBpK5KMrmvHZEGH8tJWY
u6XsNSOroyiXRo+zYDp13CLLJbJcw8jZUJYuGURtjbgm9xcvMnqsXcwQkIBeaHrAu/EDyStw0LxB
CTjgN0gRM9+22+C+jM4oJonmBbnORWmeB1LUvZZ0RuZDMBvMqUTPVLi5vd7t89cGnG3yUPH/tXm9
UCE9ukfR/IcEpuJcVYkyUAM9L+taD5JhdfYakB9ovwTPhP2xuFUuC/rBzx88/EUau9OuzCPyG4wB
u05P29ZMZY8zv5JXnFgzMZKXMCnqti8cThP9sTK5Emag6gYts1La5HDuUmBi/H8+YTH9irkZa9VH
ZJwMX+4ae/UC5k9oPpzPzQFwFnautOWvyQwfie/euhPlDHtN4wjvSeKTBcmHwNkW32tz5MEvxB6X
N+NTsn2Ql350BsNT0n8Asbl2XkNq272QMUjphG7iORZhh/G9ks8ZsnHpfoCLALasntS0MVwkqJan
0iN8dgQG3imQMUcRk69u150bw2q0lImUQuKaAgNlW+zN7RveLBCncmUfHyWYHry274SWYN9uLFu/
UK8jgnIZgRhq/rGkTsF73OkkEZ9GgFneISGZrnvtpcSHna/dlPZ53YW8Bw5+aME8wDdR+iVVFFLA
B4M/XGvVVWsgMWMtMzaKiUiHrXQPAkGUI7/xZm1OeTt8DeemUhMVDAGmr561RdpvLTpPvmwGglxS
cA05OslXOaRPDfiuL0f2BTVpxLIYEbFAIjFwppL4dQn2qjznNRwBfRjdTIMZOEZHXQujFy6K6EWT
1xgUT+BC1Z9VVtDPFsE9+YTqyU+2jEyuJFmtGLSqCZQnnwWw44bQPMgQBOMr0h5Vs2MiogHbh2WN
E93/3DKNZ6kFi2cqr8fSxlMOWq746Bsbb0VwRdDfcoDuI3fM9URsXJ/4Ckoskt8/6jPijSgZTooB
TiNVCBJmh0DsUCsz0Ih7/UHMY/eRvLz/fNYI1fzNupx3Q8POZ6mRPkPxZIP/KPG4dI+an0Q2nWpn
/lUHKUWy4PhvopnhZ2MBrToXR0KksuqE5ScF3TIgJD/OC2BK4p10mAb3p8/AeYD+0JixLEzcbJyn
YU/CkTJx5thk3Pt3LoMiWFsAnWafbYswkoTnquY6doSeA+RmhIuK2SF9Dj1NzTcKGY/gH5TOUnOJ
tlfb5GkQsMH5VAQlKmUVONf90J6CnwVTn/RmT1/z1PXjPh0khhKJGS6GRwYevof5X+pMUNeI+8++
dy4r62HKVUq8ajWcr/qoXWLu/VZlOrBgXbL6k1LpGeWEorA7AE/g7omzhDq232ddLSJJe6Yj9IHd
ZwxsUdGqlmn6VlJooTVeL/nds0lbUUWJjy9zOKt4j9d4SXKqxbNtHK/Cv5xgS4iGPziOyM+NHdDA
EqENbJ0txoFp0H28FUArlz4PBd4PVg0N3DLi6J34lPI9nltJBoPZ9reXetuKRhXQf9YVYU8tORL/
SUklsu0A4/rjPndPw5BQSrA5QNeFkS1NzZxDcEH+LWdrPoBptEEfjbh6E7wBcH/Q5VNtr4WaljY2
3kj8QglmaKynmT5f+JZyy9qO8cuFInNaLGjgFxA+YrR+imBMrf+0HN9SOJd7F9dhnvVzmH9Ezhmi
mLpPmQJ8xo3sHavBc+x39nI6qzZAxueR3kdKWECQfFM1IYos7ZRVLL47SMCliY+xzoGCj0UXuL3a
9QHBQplAw/kAQq2l4Rz2fmGL04J/J0Efd4MnpM7zC2jjoYk7+lhiKKVAWwNkBsPa6lkRlRbcwNq+
GrGZiEFux0C0qW650CF2p/E1MO8mUBD80kQ5wshr32hLgizB+N8hf57w5k4x2FEKaAMTR4+ULGyJ
2ubVI3con/A0MiAbS27j4AQeu0I+JfE0JN9x57sEIhAcY/T5Slyf/JjJJdXHJVn9HlwK5P4ovD4U
FXxEf70JpdIBN5QKfNDNck1GoPvA0AwpSlTCURQCYtV6QxuMW3xa28geZw/QEaAGNW//Mn14syqa
SP4FJFV8iSzk9JoHWOEPb7ukeQJ6ih5aJGq55Hm9uALWiUMAvz6XaVN8PTER9Hl5H+zYkomoqvIz
dnrgJMxPQ22c8GQ9OqnR4yPyIdXOLQlFq8dLbVniIFj400U6iYbWv0JZGFCS7uJG9045dJ5Fty1o
GB5P10EeUg+uuzsEsUGZklmhZKpJ+DNn1XrYYVWQqJ0e6yDyWaohI+aMnAXBuoRXk9Bwb08/0OvS
yjJq+s3U9iT9GXup66H5gzpogjkxqvbSU5cxTFy5nMTcX9/HcsScchEWYRQEqCuCMuQaxsHl9kub
VJeAUqJsqE9RB1wKjk8aMWOw249JajlHOQrz34QY9Rha07umvc+lStdOaCAIHyzay5huU+hATrqB
1253puqL6MlMF2QMNRgbrYvoN0PFnVcHDgiQUJdcuC99/FWfr/KxPehsfqtvsO+aD9x/0yLRUk2S
13WEQXJ91ZpKajx8nvxSMhccV0nXCLFQvnWwBic6LByBVQeSj5VaHki4vE8GPjQdZGWLyIR8twEt
EYU/xdQK4oAkhVHBW71onxf67eRSFUcgtlpGsRrBUSYaSOd0v/e9w3NEcHNwHQ+ROrW6j7bRwdwR
btaAz8XxncSwCbMwtCVgYFyn9qTJMkBsqhNLn/WFSVR44doHg23wegd/4q3bqacBfIAIbQYJuJYA
b0Q7zlVq6tTMHlbJ/44gMm8ic0dgNjxM/lA2ajDWu025CNTnMgOZfiUKx0xQSvSAs8q6ZaMMOrCF
Ra3esBKZEp+f0ohrTta57/g6BliJPen8Tud40A2iz4dHkbWOvVe+Y6sKKJTLB6cqITpRgMuHAynq
NThBJYZdM9mSH/nFYcrCFZXx7K5VtJ0QH9wdzNWahszk9tUZztgVkuLwuTSEwid0pZlL+wfso85D
ljuAfdudIzWTaVsNrvAv3cFBs/j+5wT8K5yNs8QWUlqetcFx6qJLJuMP/b8pxqubpvfp5bExJACX
I78PXr4CSzH1LB7QDOQXU7tZzb3KNFFp834Q37fqQPNCdsSRwyWoE6hj/csa9tDq20MVDOimuj3u
0hlSp37zbt8OUypvlrSpLEQRyzb5JvNUAmxlGuV0ygtLJqLnBCqZHPuCS89UuEBLC0YXSj2X+ZQe
kqP9VQ6e/zwZm1/RlrdLFCCbU7jpKdWXZYMFzlxu5iVnu/NUPn5K4++FAs8nqvSyeeHzgvkHILIt
9c/z0rwwGGU+hCLmpggMg1Jlw0ycKKKavqRv4O8OTV4EibwrymOW0Rvq1e2iavPi4Y8XDpd1KxMT
LjubrJ0JXDXJAVjTQOEjq/YPTGJbHZZ9kZmAXbEIfdnVkcZTMoC9DwWYbGRH0XExQbSIWUKIOU1Z
pWmcLQuZIZH5kM9LlYL/HAqJaLULGfAFkLzOcQt5yeJ/f52LCeSr9vodggfW9UJgRotY8SCHFTPl
cAA02bt9wLmeWwR3Yi7x1hRk5QbU1K1crBBeiTZkCTnLlH0hcMukvmYgbfAamdFUcHIyHrlb8bxk
IV5UcAeh9llMYfDAX2dW/7QY3YdLxu9fXgoAYh8/ad0VuIdNmsKIs3ItIfzLxOlyhKiIZl6O3G1h
vsrQbMsn2aLFHaEpPmgspuo/QZ7z81N0E3569QCHKoTHrCOhkqs1WWcB1T77z1S+K45P/tnzEJFu
gOy8JW3bA3fUX1t1Zpht8w71OcHUzyXa+9xubbOd9qZKEs9/uXhylhc5wMOo9aXXK/l29YdDQSJx
xzus+brUxs1lAIAh6ZViuKa8Vcq9OBxPSQWXZ720jT89KSFweDGzd5G5HMk31PpxddKG8UQf5MlD
9MILMdOpwiRjyzQR1ENDoQ45kGBnIgoVfRfUwIG2ncKN/oW9sqSj+X+PEmpjWCnub1eygdnDFdIL
4nUQN/qbZuurl6rDurNmyCQtNcxsnptf7nXydEPRDhlZJJJczQFdOTOB50VDLGvt56rNwXI5vDUY
aPTynwRRABbZLhJWAo3lw4g5NsefAqRq/eZSI417DvmckSHsy3rLxE44QYjFYem2Jvcp+QxpfXbd
kc9OVOKrztiFCq+aWH3e31DJYrqhwVkUyPHsOu+SJ50Wc5vku9s5R0cKQe5hfNHhGtYhfePb4nEF
mUr39x/fJMIik9Bv4wAerKcBE4m0z3LK98VAHYOYQ6ic6K1UZzO7WHT1DbRjVE07ooDTXPwiraan
tREJDJvrtXnWFNlHjG9nTxlXaPb9GNw0S0/EUkXYrOVlqOgdunPVMRlXbuG2z1GYBN2nR/77bUGH
hpYdXoH1XT2+Vjf8L6NrkFd+88gjagVIcD59VOxoLRjrCwrFddd99V/00d/ivsWqiE1YX72FIHsP
Xd/ALmRrBS5JI06vRV0q8swFi5PunX1D8qtyfaZZ3pSkyVb1fGohWM0SunrtT3YnWuMbsP70bu0t
zDtckdQ75YLyik9X7Sa9C/pFI4WzL5PHGpnT1ypMO+S6Ti7i1xJEu3WHye/S/upJapOrlCCPx/N1
ANq8co76bWG4pOZplogvAuaaUJCZf5XVDH12TeI51G7g/M/Ay9T2aTLE6fWIghN9f+6qXbxLUmGj
gE941jpTF/b0vinJOPdPK2nbdCgKswvMcxj8kjlPHYsJ6LZ5JmUQHVCvu9/JBwhHJjoHC7n0Zo0k
HghLpl0rm841byYOs3PTVcU7M7Tk2m2jbI1vhLBFmAVnvI6BIv0JzD3TcpI6YgQzqe5RbsHx7b8G
q/3s/gmMdXD/XHvz0tsuCv3IEjmTv8U7wqDeiC8ZgDBuo4B+1s/LbtF+bcMuS0eEXSHBdIsFTlEX
w3kzfNQQyqAkc1Q+eYWz6SsDcD+tPYCF4sINcUWzT8h7weTS7L2dk1FrLEi7c4qjbfOarY2YTkLE
TOfPUkvHSKPlAEZFWuhpVA/Bv8oF1cwhl08F//SDU9iUDStOcchupCNl1rgZ6TlqgiKe35R4LZxH
o/srhfn1jKRgHxT5hmJvXwmdVM1SElh+7tpVu/fhU9YeYm1KhlAsWRDGzJw1/vgvgqRHcrieWuEU
jkE+akvYK/TpZkteEIS2r/XeiUSyV4rU01n3evL9Qc2TcEa3RtOLtuvGdCwxj3qRH14FHHUJlsH0
j2D6+GZMI6Y+qG+5X+PLHKRY63f97Rl34A1roKaLTqAWqUXmbYnQLojkn96B6TOJVbSUmdZgIlOK
80ngE20AJxqYDS9+So3FTOiZzpM1U0V3LB+meZa499JT+8LvDARz1vjZCiP2XZnEcS1MZGd4QmSd
h9EOktQs/NRu0bub1sOgR3WI6NNX8neBFMvKwNNNZopoZWE3WIJ+yTRLzvFQDBgc3OCjSySaxLzP
eEdq/P8XImAb8i+ZarA6wNJReiV8i+MTgNU5+sfw4NdgTfLlCVkoITzTpcIW5papZeidLWmnfjjk
tBYQkvZZ+AGR3T/o5A5/KuilRw7OfaGKdrxpSJkSsol0OJJggEvQwYnDBuVcjS1xr3yiTpXHbEY4
s+TjORD1JLlO/wzODiFMQ2LglNLZLU3CFUuuSsc0z3TnIo5EmKFUHX/tTcnEq9naBA9d/VJqD9ns
8/31I227ENw67+LxiSr+vOKYUULpsMyvyzA8CzRtQYO2WciPFnWNGvwM9oCXLCdOP6IHymQvgOnn
2icu/jCVjsMZ4A8H/AketVmvmX/5hKXnO08b1pClYOhMCDXWNd9E1rxh0SCpSlD7ajKgLv/OoVF6
D6J+LcrkWs0EeTQmr6T1vnVJ/qzhlB/sB/IlE7JFEKPTfMYbqHZU1Oo9jaKp31T+78VgKSSFKBe+
vIisaEkF/QQiNYMjMHNOlQPBrqG1lMpJTPpgjjtezQgY8nRPejKau0c9Dy+feJuFNKO1ABBtSonx
Y6WwIP38xWLhjcSBRAS2ctiU4R1QW+T4CWWxJQ1u175ZlVz67gjnO2z6KnyhiUb/3ZEZeAtPsFcP
uxJNCH+AReEw+hTTAYx7uzxlRZCSl0TKsxtSIF5v3frUDoFlipQVrcQa5QNic2gu1VaR1o+SQUku
xNfsobTSpNxF+95VtS63s2wJbOSMS1F9k7t3h9+yu0ECH+J36IdEm6Smb9h8mCc5D/sdhrhZWenv
Ry/pT3u1glH3xmc+0QhdXcpjR5CEbgxc9fV0jawCfB1NmlAM1Fy5KaCx7AswCrjy18Ijem7PRCcc
uuHNEowduEtAqcEc1n5OneJYeA1yrVI0qfEqyqM0euqcM/BFHHdnyZgRbNcpWCCnLq3KdRJ1/ixD
JECMwKNp45QmlnTjgx9luuSRbkzsqIHiyRLXbla7DpgK4eNHGbNeH1NSsUcr54d+pk3yq+Cv4ee1
BCGVVk9sOh8xab08AYXSoeTksN4o1w3by1RYfv4imXhflJgMCEk4TNArrYmfdrrRStteSihLkhIQ
GJuQIeDG6C6b11hRNZwlCHMy0XWf5wBoHkK5v59Bz5/bWTS3EKG8QQVG3fb4dk/UCJeK6d6pfhKb
8KBDrAuPV4u3/gZjp6Ml6+G1nQ6N/cdefNvbnyncw9Ygggqb/Xrj1xaeBDJZlBZsYedgfTe4lhsn
c+Vs312BEoWQ1Ekaly8XABs8lVBVxBq0zYTRd7kt3n08Vadq6bp1BmFYNJLNOFoPp7C/8xhAXOYj
h81s3MDNwyI5hwO1xP0PPRYw/6+Jj8351ZHVIH92+lRA6H/mArvlVj71/HR9pNkMwJMl17J1wQZK
4seR0DbDuwE6Fac2YCsAcQZ9xTrzTJULfqaFn7+rVB6N6feHTVy3SfJsLOhahFgEQTVZJ1vnpimN
tbR7CsaqriSZaBExW0yvgKEHeUVSSgB1u346hkwUFDaPftJ8yUk4YHzJd9uS/vCLZv4q4P9GEiP0
zOfE/cOrITdJE+HbDYi2aWLnYc2msn4nVNslnkDtgGWubSh74JuVmpPw3MqlspAK4HnQ4LCp7IV5
f+H+1b75SKFRRySUanqRm6EZjSj7D7XJ81wUrlOmNoQ7TAvgckjGN9g/KrdMHu82SDl9WQyq2KpM
MfgZCRvaS/eCcq6giUR+3+0kojIHaPN73ajapdPOBEQU8nwmO5VSJ7dQ1rfBMbNh3mQclpWnifnq
zxW0WP7bKC4Sa0jNpEaW+D2NLyC9fmxrlwYt5/BqVB+HaBX4TuXKDAIkqhVImivMkChTbmWELEf7
sOjQF5VC8vOR6jeXzXALh2y4IftH+zAvmuSxJsCEXuxl0odihsCcmwLqueEEj4UEBCuWlJsObZYx
E1iMeYmwZazxH+lfwtscAG3FnVLVoePz1xBM316MK2Z8WLkDr0vH+u51ryPKrLJSPpfx84woLxK1
XjCLhbyK6I1Y7FbOjawkvZlV5R7++hpMRc9lnorKr1ZqBZiTcTMMqk7hNZMUMaXJgdZavMrxLq1V
ILuNRO7n3xlcdv0/naFU0kCIia7NSsnV/Op1BSYVBnSBlFADMItuzcxCfjy8mC7mBnuK0kjvbe48
0ToHtMC+M/ynzPZy2VtYLptSVdSLsqQsB5eO9micN31JAZr8q7HPulxvKp2yPDjgyBS+yZQ0xAjC
97YlP3RBQ5GQFY4jyR9Bj2OonOzjR7lVNA96IxbMpSxAw2O4UyIfXGf2ngV8xyXatjbvVVvQARab
Xstgu8a4+xuyOZ6j7p8DwkPyDdsWqLetZssUPO7lZkrpt4Da6gJxNluk9GhUlsNo6ihMCJ5WcsBT
7xm/Wnx1A41/gE2uvZyP1+OeZVXk7j16pkH52e6Y8/2ZZdFbGc1M0qRqtYudseG4KHuSu7/Lv673
zx1Lfs5YG8z/NA5K/vOB9KgwE33Z3O+XSuKSSZliC+9uA4s4jqD7BvIXDgg2K2z1/xvAJvQQ47bc
fmIZLdp24D3mcxbk1iESruPDn6/v8u9A3nMtvqQNqRT2H4Y5N7Fx749O2XszhfuaABxGBYRRmFp3
Ppysl6uz2db3PgjK7r6GXfvNF17S+tzBHdd6NOUax3O6X115Lp73vsnLLl9waTQYxUSBLvjRuGc0
VJI/vbGQavM/QzzCd3hy38NtJ8NReYPzheGcWAdh8S6JJCRadZ6ijE+P+F7mKCxli1RvA3CU/TKC
Q1GTpeKJVi7c7JtubwbfBZ/JiZ6Ka1nMjSRDw05CK21hv242EVoPyvtLwKz3XQfT1SOsw8r6T7k0
spctp0Jf3zLq/akz/Sc95oUS9KkCjmsCbQGm/BToTdKgWbL3PYf40YsbG8QECQFwNWzpSRPpsAFV
JVpJzZ+2Y1uwSK9bnIeLNnacNorLKfIRqcgdy37Ub81R836tiwDzpquynEBi+tnmeWbSGU8DscP2
YKwshAMEGniz1kmZta1BNk1SYkMWgpWFueyWad7F2u3NYlFqCm8W4FZQGtYlWAP24a51z9dkM5YI
Lpje94a4s/n5D8gC0lPgzFzOQn532TVpEWmgd9NJcTnJzYfikNhWGP375yVUyV9jrp7fGFh39tzY
jNd4/Kyh9gN0bfrIHoC+X4uVz3E24ZV2nuDY0A4GYj+TjPCgHSqkV2DjBfhXB/4PgyMQxT/PcKiG
SVm9vAJsVLsjzjoA0GZiFwZ4Su+AXoea5IFBZKr0L6sRNYIw5ItKAe3Sv79WGiVP+KB2YXyTPssS
ZAMrgukknwByRZTGADT2u1v7sN18htiLMjCu/Qm21ASHShmFDOmMKwl9pDhn5kzYf0Y83wzgcvpS
SwXOf6uabaNhUxS4RN2++rvaOjeqWEJbF1P1zf4la5NRZhu6x8X9/amDD9uBcHM2/T1KkUH4Hjuu
8OjBLzzwK3C2vQGeSY+sctrKf0tfHlpmd+6t0gtZA/CghKVsVm7/WRYgswzuKPhPJtMnlS7aqJbk
cBNp6sjgI4GGmL+RhMyJ42dvYmLkwvvHbMqg1it34CJCH6lxXfoPZ+MB2veuDDsmv+fg1MHf3xU7
EIS00hC6JyW0yfCXdk4We1lfkYj/42KZ+/gdVXJ67Etz+UayQ7C6ZWGiF+vpjjqzlTS7g3x2cV7k
ghS95sc5hcrtgRkGAsNUG8qYSDZNZF3YNRQRqIHfA/iCgqrnIuuVliXvVJ8BvQscT+xkvXv1Bcs+
1QGj4bC0uiLtTz8Yt00GTYetQMGuVJUor0AtlQS8FTf0f3NZZaqxTaTbLmdUcRt0xIgxlLGcys2b
qzxUhddo0YpoyXoGzHhpaRUGDulqLPfbH7BqNDVW6FFOo7iGJMmIKibs2X0dj1zRp2kiXEC/iYZ8
s7N5w3PWBKkM7qgCZ9SSSm8xi9KyB4meeoKL7qdPmD3AGnG5OYIZdnwG9bErnLqMLShABFdd/7VT
ioxYyU4pDK7x844KRAp0peGc8D1ZUbJQzUha5CSiR9I3VlT5xr+ZGpPtb3r4Fc2iI6NejzO5zKA8
hvVmYm3WVw+2iGUb6wK9kiMP6abcwkOAjW9wnDAR2f+l+Q/mcqEHvQe1kbTX7sC7A2Hty8lDjOnT
t0A3fc4YJn+VIZ8vApx3li6SQLl9fRyQ2aI5HY7dJB/3GEnk1kk0g+5H3dPkthnTRSkwMYvPDwaT
b2O+S0DdmTjQfOPQh4y2AX0uMR0R57IdjdGeKzTRGdi79Ojy857b9KwGr0vLamz1o60vi5fOnghH
fSSBKGiCwyE2eOxoTLW958f6WRtB1V/3MaroIPCR6ZUrcuACuM2WRQHLgxq27xXMEbMAA8K6ygTm
fFRTLGiGxVsKq/1PFFaO2MjeDg0Yz2bkgxsFA+RFgh8KeETtI1Fl3HIcyvqvpJg5hkzT/hLOX8KJ
L8WAJRzkJZCMBOqHlpNtTf2/5SZH0BPmUYl7huf6YHh1bqHCug5sMLvo4i6IOBQ/TtZxHD+zV2aG
Rdw9XtXrqf9TW1+PmoFLnWiIYSjKz9eNpCxpmNpG12lWZ6Hms9qyvvKmV1poeVbGBboMAJgLieK4
QOp5i6FG6lHXuhJrGG0TsZwzwLAog2KSPyQUZyI4eh6SM5KlMDdm2sf5Lt0Ydb85eiHiTmlhdc6z
xrag8qBlYgG65xdl++Sxu99pjz6npAkQMIhU4xb7C+x6iFF3nLBsZg8t1G9JovOxjfvUyxoLwDBq
y7+OIvV6YaZgarEYuiUiNfvFRK3gye1kIwGj3B5Mgr4GNzue4P2kQ0uYZvljgq/hH97sjqSh6nOM
DuY/5glKHOkmd9WCETk4snUdBT0PZ29yS5Xo4tx+W7t5AUA8iIygBAGOEYbEm3iXAbDYHZlleTNr
wxr4mhCpRiJ0/1xTJJ1saiPB8W4PjxbPGz+DVbNsZVwImj2DafoCOeI/icY6ruhSSo6BKAuCrC/R
Deg5bdwdJaA0fbqBEbZGD/EqdP8fupuPfC69Ipau7Ap6BimSDFObF+fuhLLuc6eP06A4gV3vDZ4L
xYfVzXxuTM08rFu0hADaN4VNJ7yHElnqytzHlzxA9CaOErlM25ImTx4bSpM03WZNZcHCRrIvXFgF
qdxzyiDENdkygngksz+W/BvsnXvWz8ad4L8hXWYI+q3RNmlvlgJgImnluZb+sRphTTrx6ic0UnCi
X6aKKF2gz/oTKTVxLtJDTsti0UowViTbgcNlafxG9g6Jqr2XFR1sUtsVooxLcLmyvucrdAF8QtYt
ohzZSOw3nalmcvZXE8XSblfF2qGKfcXOX+PjUaph/NLcZ03XwADTvh7N+zluG1PdIySgefAN5+ZQ
LN8GNueohR3KXp2WH+O4WrCDxkznSBzv80BwsQS+ZaWaR33U2bkaxgUE9GVIhIvEcZ7GtXv07Lof
fUVYQNARy51W3t+HvvZVn6kPAnP9DCvWnwDOTJI/VtA/PJZC21i/o988OIYonL0PIKljsl3boj4Z
3p0Kb4qzpebtPGIZ9NFZgfpO5Bpae+E1p0q1Us/wjT4FySuXN9PGJZcWJAgwSHgRFTg+8Hmc6K9h
6knNBdgQQ/Nm3YMVuCcuq1HV0uKDOznh3XlvyL36wW06H38hGbNQPCntWJ13eTkVAWGt8SrPgNuj
KbfrdHJnbVjdTIcNk+UDKHEGrvnhhCj3NRXwBLlolY7Gz8ZzYhUiLDPG7m3H8Y890VTzO41cYLCf
r1QRD3qFyGBbhAPcNijPnKXsbmJDISAsQIQP1auh14eMW5tJyRNlcbZ7cycrvhZHckqQIvwK1H/S
urfdTpsr6Y/QK6AlUJfOtKQqspkeI70MLWg7zhsTXfoI/+0fPPDqK6WjXHRIyVFCAWVQA8RaEurZ
yRch8QKzoqZLXH/7ogfdpVOeq/9h4IOGl85uMQwTVsHjxjDAYIMli9uHd8XarTuoM4sbgPWSE9Hk
bfpP4B7hrNrjQm/KxJO/8VGlDmJkwTT+M/19RKW20gFOJuMK8AOnN2cCyoblaPGPy42N9xBfUSYv
iQILA0L8xwjDZ6c7pQO23Qruyb0R+cZTi6QPA+GxKKJbf3pwsaEvE1nkElrB+v9kc8kmME+oGuFy
DaoSxaUt5EHS+Ur1KMmjyHPOucx0P122U+L+AzbZE9gAJxFNQZMUxEZiiI/Z/2r4tweSnaM/dPMx
wVihCMCJ4ABxGRk+Jq5yOWq23fNvbRMIeenMlUcnVYFyPE3LNJMcvRDmKIEmptfwDLLxHQ3zGFZh
ivKm9jwB0Mgj66tpPrd8UlyhdvTZOTPCy9FAcLw0jaKjSXAuw5EwY7v52gecobBTg6oFCo0lLIi0
pbrjW5P5vq1yjYgdef13v76FhDfteD1BrKBT6L82p09d3eZE+L9u1rHqAE4UA7yWTNbQnq+bfI0N
A7VF/cZdFDQoLk1C24ORgX77WIJQzCmCl1bnXD1r+uKkS0KPKoK+6lPgeBxNnioLkDw9nGmp7R+S
H2Nzywb79TWdzDSthDBK92DkbKQOs9+0wTky1dB0bds0+WoQ5A9vJ2h6C6PSf+WBNTeyV5nFjDbo
kSVmM13DJWRTHxUAuX+Adm/LgBgp0jTaQKN9gCxopDHpSDsAk+ltCjOR1krTC0MgZ2+ViYN0M6yZ
CblOzEW65rfR3xO6TSHS+bsVQxZQDtUtjjjyghhh0biTteR5S71KUBq3tlVWssCtddPuXuOOHtnt
3pU8MIZJlUGcj4sGCisPHh4Pg9BiYRXNJFDhMYVF/mLrSIPOc14fy3oBS5pgnnwWMXWArL66HwpE
KWhz6pBaid00kAACWXCrd1xpUyaScPHyzqQzMrMltpSQVqI62BdVDfaMvqDccZUQ3tt+QD2iJ8BM
r4DCEl2D3rdeOi0f9/VJaKgXimX231AUQk9GJZox1Lz0aP3W9Gav2e218RvkQgJXYc3P2OEqyYLw
uHVtD7CvJ55umnytHh5SkI7IYOcc9DZwrX9j3Quw4tm8Q2ID6c3fT5JMLGergs1ObqITX/o7+bIv
mhX4K4DnSWfUiIdSYL3iginsaT70o9NcGg0MZrIhAU+PB/BDqt0QojrzMyrVeFxMFlXXTvWka1GS
w30saeYtYAjxuVJCUL4pKWLuNpzMIgz54IK/r+3AUq35lVFiaIQ2Qg0PJYAgV9vtLQa9/gfeX3AU
1wl/AQxbgYhxUI2DSVRorYvxxuU9ssVAnBTbbomqaedaZmhTsQE/6pHk9oYqvb+wfqKDuBLnXFU6
OFuA9dVg7TDwvyvCegO0zXW54V5wpgTkG2vCUXcYNwQXWLR+ssvkgy7IdPeGli72pLhiphH3bmjX
wnG/+vNTbJYcQ7fZFHdfzJXSnI5AW380klloIpFDqfoEXqulLGHiDug1FQxBrNTFcudnJG3kpHYI
dF3TZ99neHtUgPG5oLExEHbrD97nIB6JmxsMS/kYlsDXt9agQtLl+1SSlLEEgF12IsgNnO965+TK
MxaClLNVp3p4EXskNhu5O7rIqTvxz3GVL2Y18n1dDB0n5UskTL9+BH19g1bDkh6Kd2GnfDYgYaQ9
kWIOpemBvzn7UGfHRTexcmL+XVgmQT4HPNt23OCuJEXMZdtbSiAOL4xwwVkDR118uN2fNF8MkqQh
GIpStWO4jYn495B2/bUy55A44lnVxZYdc3ab13BRZliTEcF0Ryj5BPHb3gX69UPXj5duuyzfXXJ/
6CHI5wFqHD9HjYHw75QJ4QMDBEUIPWT6Mv2l8yO9Cndgpvg1+IGemk59IyF7dEJ2uo7xMPVBpnOa
fLrZrHz9qQu3rG4Hur3j/Z7PaR6GbKCPwKf6wRqon8lQ34R9JdH6FYqiQ4gM64V7lzj0crfJozU5
2swzQBepaLwbiKjzI/B9htgEIee6cRgZyrmPkLJODxL4nT5tcj2QBYFcOshtHLF1iXZvQXa+O4Fd
4abmI8oYaDO/R1w9hbWYof2ByFxIOoteJ51/j2wa3RZcYXMUvQH8lgXWkVGpfZOxALU1dist0udd
auocf8Mek39IckWQrEPPHjEezZX5UY7Fu/xkS9LpwF1iT2KKQN2klx36cB8cIydiw0WT0A/FY89l
NFKnD36p8/Z+TD0SoSiJdBs/Efs9VVawxy3voIhd3Q9li+ggJYDN4mNu1ZXt1yqckqXPrvZhBHmi
2VEHTl2s3rAoYawcVRnuchQx1luT1SVFnzMuPJw075WkpWzkb/64q57l2HJK0m2Ac8F9JTS9+o+M
f3uGHfkspWHrCyZGuKoobWWgKF51UbTuwowKYEkHnkTQO3ofwxCOANtvOqe6eSMYoKLiCOTMDLfr
pmxJ+I+F1cJoADwmub1LuGEUtQczz8AsbLPHehK67YSfbzZRcVMmagDT/RdwY2dmUYh8mbc8klx1
udlb7rr46VtpYAHr0RiWL7WKKauwSKrYrkg5to5TDjIuaRD+ssTUwKhtVxKejV3kEMOumL8yg+tD
o7WUA0PGof3xTYs0hTu/asfsbh1FBY4/JkZiqKyTPoIBo8eMR5Ko39eSHvn5eD3RPgPWE4KPr8Gq
198aEFIHJDDt0JLXgVIQ9iJ8SjqLKMYNM10qxf/NZ6OJxDSQVwq3tUTzvQKcRKXICBQgvOmU8Gns
89yYRUNowliHue+NNb0Jjl48jNsKQXx/L46O4uvjYvSFNOx0vajo1zqc74//1xDPNycUQqJarC3X
8zZvyqAgf18wiewvVcXEGMk+cD7Oh8baOmDqviVlItGhkInOMvw0RbgKL5GmqTtMfpl3ZhLYPBuC
RVLmw6De+DdKT++vAtXPc50gMu37s9I5gE6mF4ufw6Oy0CQ+bMuhCHiNgS1NfWSKzzJ4ObKmqzTz
90kjdXA0ulC3kuavonQLPAZo/PlpGo/e0Em9FtCmAaJD8RsUjmNL9sBBxXqrNNoFjrioi2ou1OBg
r5EfchpzarITZyraNtb4QtCkuvmL4ISnRKXo/hlkKJSVVBhpjO7/THXOKObSz7B0P7KnQgsPCebP
f/OapGLTCQacsbr0JnbWqio8Ck2V8IHYe1mj89AlRufMz+q95ZgvWO/5jCT0s2IjRJdrBgDVwOPc
QLneRf87M5qkg1Nudqjj3K+lpL+FvLtJWCh6x5SJKb7fSD4kpdI8jeMS2439sVeZctjnft8jT1ze
rejImPXR70lmGWQboDniPG++q6H6rUWeyh6+ScIehtXO8TaM+iZys2aY4c/0J6tb1FSjMmPYl76b
4goMLUEOwk2b+oL8amXuEdIA0I0dpjP834TpZ0wdakUiQ66t9hy7TBZvEGnjI68vPxuKyeMvI5p7
GFhSTBxWDKOk00kQt9oWeOI7F6YeVUHYirSdhGFrb6455YzGPV0H65DElwL7Xz9hokTuKHuEb18u
EOxX56OPe814wY1/9VdB7OtYCMRPrwnLZKI1zgI+WnIF3wP/j/7rUIg4tl+T651Aam2Tw7Jq2Wgf
Ci51JgztWQe3OUh1VA7JsQXkIU06/c1h9daqfFJNSVNqgxCv900nGmhiPcvMih0602Bzqc5MXhEg
dQCUxyhfcItADytGPme/7hH8QKKNsC8Yo1VtMiv4r9pnyvoSi8n2pw6BklhMHaVSYvYm8zBQOfgZ
+kg8RfaCq8nxoGUcBmILvdfO3qi1IJ+/5ZhgvQQEIVxZwUYeXcYazVkySWlxqCRXdICMJTmWLPVV
L8Gn98wBonofTCft1MbezVoUAfBRJuSiAXPodnU81bk+2RxGeLTZdwY1+ebXNqpdP8qi8vXy2DFI
sYuyTWUa1hfCddBjY0EL6E31aAb6CiKLdR+f4w2gKC7uBnnj1PywqErDlvzworxpoZdvKc5mlW2T
bjHKrILEzFnZOn+poB/k8eySbfF5Ivgmhl0/3hmJHu8jcMVsZ6aSfaYB8MslzZMAyRmP61kAD20J
qTgWnh1qrmiIw134cyG7s8eH1kqui4cPSnMWkiITzKTgxMKIgAif5CBcP+EMm4zZk9BXwSE5u14V
BNf1w58WbRqGlmSllHxBRK7qGBXmGKiRUE9KFokK0BmkYqargYom/5sBLd2DJPAIbwOXPP9SeD8k
+SDchMDE5UlY2pH8B2eUElaUM/UMrb+Nz3Ync1ZVVI+qLvyyaNNCxm+yV/Mjoo+idDBjd8TmtYEc
Lnuuy8cUi2Tk1FgsVD6u0MAxMY+FI35Y9AYzlK2Y/Jyw311ApbK0ojIfROEaem0q7QMU+Nr2O2NW
Jz8hUS6BL5rc18TDW+IegOSaeln+lzniQ+1BzYedfjWOnj3E99SNXsEQJq2r0R6YRR7wQ98NRK9f
YRJzSrsTIcrMM/lOj4t+R4uAHNLRlGx9zFRpIlG1g4H3y6y3q9WNhas8XoBULzPuPbaBwzib7BtY
Wqas5Amiip5RiXrd8UufeNQNEiBmFzW7O3Dx4gClVYdjLpTeh3Nj9Hns6Ww0IElYuyUGeUMggKPB
DkVZ5kxaqAP8bVHhB/+1ldDGblJAcIO7cHeN1+mvCC+A6+KBUwgptFcI5ipONHqszMOMbXzQjUfe
O994XPVvEGYpVxahqxht3PJ+ivYbwjYEGWhYwf42V6OL6FJUgPzQb04OPUHPOSKTNKwNVyMXzOTL
F3+f03gHMu2eWQmZ/exH3trN5MWQ+bsqRWVJc3nMYa6TFJlfr3Lq1JDOroTiTlEFVT7qPwHDa1m0
nEDfTlnpe/c0dF3QePEvSFzij5UinR+VUTVtA8ftQ3UK5xakczTfXbEC8vnhiuYwriB04RSDDJQv
EUsSZK+RvFMkv9jgIJ+6v1XUBlxxCRHcMt9rl4U/xuAAXnpJdLJU8Ogo6o/2kmNjQsHEUG8uDI6r
cNIIOCM3FWDlrqeeEc+nHX+9oVRSGXwi+e4bSl17m4+EsIC4rMLNaoeqcyGyJEptc/e5Mm68EgW6
swZkIF2LIrvh26FO7ts6/Aak7xgh4f5x8cgtcX3tZlZlfJSo+6Sdpbu79YyxwCjCL4Puxquix76P
crqv4t478AMc5mrpGniMnDjKrB1iPI8pJH/u0SlNXRIPLRdDBO7QlOCWuzSo4WYYYh9OK1p5r86N
py4d/5XbDIluuTPxqZ9nSPmcFm9b4oZbsqtiWIx+TGNMpnrqN+KxF/F/5As6mrgE2qAUU0YfnqVD
QCU6ANrHB3YqUq93PVavBKd0oIaQKpq6HvxaJUT6UkNOgkP+QzH1PZ+U+aptlxywk3PaLVd11CjY
nG2q5gSmEa8Qzj/YWIckL9dMt9tlMpEZVxfkx3CBgGDZZcjc/TjPf8vr5mb6DUHUZi6CMtFm+IM0
oKq+RCjXcxjDNC3dp0vyY117hfaFmNrRenSU465Tj+FmRwFojLUqnSsnRqH8/ZLqqoF0VdnR7Qbx
sJmovatHM6GkOePkaHzD8fM8pypy2N+rPB1bTihs6/b50NGHH7LW0dHM4YLH/0xlCE/4Ov8dIW0K
1dJmvpIpAZwXxXLp5Sl17UADC7LoIko+Xsfl1W1BpdMKvhzGN2FU6WhMLJ8h9ExYLPvyPj1KKbDh
5ioxMHCx6nHA7itQ+E8a7kVP5qPReWFyLnSumZHqPpIwrBM4KwTx/3+vqA5+zO5u5g9iM3LUgPY4
Nvo/3EEGWLb+JyVKp5+HZ7/is/Zo4wjhQnZuJkbdYyBsOUAe9nWa1O/3ctQo2YC8f65cF333qCa7
GE+HqjwR8FW8eN+IaExZCf0T0/kot4lN7lqQl2jw/3YTL7iePSoEwAFKuf0kyLHVvHOhx5GjzP54
7ZiIpJXFJBbM+ZH7Z2UsvPgoQucS64f1491+XAfMOqO1iZJVmsklHASu0Sp5VgDPfmHNekoyH7W9
J4oUYAb2+8Dd1olpVK8cKdJ0z1RNBSukLtFvYVUc+0yal3nNElgWNwhcrq8JnYT7h5XETNagVbBv
v6wHbwD5952jv7N+iDqxt/F3SaCWi+ZygYXN60rSq4KK07bFV4dt/rlzcCsx0LXN6cASHyL8zqVX
5sr1ZGmLFrntjWz5MMKglsC4pqh7ZfZWzOm2O7soB7Px76jSlRtx1shNb+GmobMThbCw4h33S4+D
A03M6MCBRYwa9crLmyZM0GgY4zkpEMkJ9OQUi8njyGWTkalBWdz4KY6cDZJeMzAsMsxKPpFNuJAV
sbC+D69RM0xuq0Sl8UXggufJZaAnWJ/oJMFliHCW0ZA9jeeYwS4yoi1XFWssWon/AoNx4j4JrOiB
ZnVf6TVVLyFGyM7ozerTtfZTatK2S/Aj97jWaz3qpYNHy6PseePDyWrzhp1K9250qIS1ckc5IH+f
fdXP4I+4v3nh8ir2d5FMo3L83CqHIyuP3AxNNipI+/EdfG9vMdCw5Op57PAuJ1rYe0OmGKU/rZzM
oUcwMKtmEJw4FBAUJ4Cif4SrP5pE6EJvviiwblvCNv188FjpKWRucKg67oWpO3jMBzQ6CppeekeE
aZrzyf85PgEqn4Tp5WQq9gzpa421x7tlAjLPTgh6MlJ93oiBW2LfFxrDhK01eBlq85g3rb9hxiNQ
jjWODnF18FUUtfPQP24mi5GYB7hrr/+p8+tvvftk32T7ADfrskVeETcbGi9xFr86JCGaPEXo/D9S
t8xpAIjPA193vY6ieKGFpfru5qO3wPsIhV/rW44kQCL+vLxlfFCzh4K8y3JHRpGXSmeegaq8LdG5
6BSMyQDY2iHJWOA2bqgXXfEEQFCO1w89/mwlZGWPf2nplDXx/b//2vN71SNxR+CULWq98W65YBTE
SdOdivZnoF/XEuWDfU7gDRtRtmz7ImG3b1FixrWDA+gonQyd8w5ZWEjWJI6aKLIPwRPtCM0KJt3o
tuFWIdDbMlO/O6R0pDXzIjFkyZ5dvy91b09Z8TqaENWcpP903w+htSKda/XXWEuHPSTX59GZxGcM
tKk/KF5MPFggtTsTBTIpRbq9V3O6fI43xnGbz8jGtE7HhnhT5ItMdqVk2yzl4oFOiaabNj70QnOX
XDlXgQnBlMFceEpvS6lno+IxdLpXzzxmwH4IQMtnmVuZKr/1/Adq18oMIL+kMvkr4ZGm3ZMwH6MT
+/mddrRIqJI0FiC6/Rse1MokLjPSUQWpF6zNtIKPyGgjKPVWJ87BB4R3Wkzu6vbn4pruCQNeEANb
tvAWi37ub6+LUWIFKv1A7K2HIYvcDjD9FQdRiv3AOZAfk7BtJXEElq3w1UrrperrfmVUHogaPD5c
D9+gArwntNZDSX7KG31V1OHNLeTC085l420J4lTPBBKGWQrneATEI4MBBNDqicIcZv63pL0auWNC
S/tX71Bjw6RUz/GFoamr/TDmsQ8tqv3+aVFTj8KTBp8l+CCktB2tP5RywCsw4UroMnmNZnvbrPZ5
gNzDPC3wSdA4OJd/2hLLEK/Sz/YuMDBwYRqYmzfnH/dNaS8UeBbqdHF+G9sLNP2mWUT9m+rr31va
sQhNW8Dhb5SBQ3T5eW59uc0Q1ZZ5Pl/8QOTcCgNpSjiWLV6J/+JwlDG1+jRFeEsqqBddEn7sR1aY
vSj1odQRVa6H6BIxVxd8t4DCxwpcIjq2Wq0zpBCJYTeEnyjb61QH+olFoLQQ8eusaDsW1hH6dNhU
VsfrRb5Appq1FbCh3veT2ICBm1oE4I8Qi4ZHf1BHNK9nQYF+wngkTau45D62rU6Jb3XEyEon1/Z2
7EboU8ZpABiGMRPgnZ+uC3GSavClBGFy6bJFrwsEVU3VHzEpCYy00WxeSuWeNapW1QkO+1y0pTeh
jvgzqPqLl6n8BXijgCMgLEXc8i5F5gE3AzbMnZlYXWEoiYGN/vFNPOJ5gAj354WRcUmslsttFtZm
XeFKSXyH6+MYuded6Wm0OvrXeEZM+w4Mi+fbdtXt3yqML6tdZ36laU9cLD7b4auVs2SnZg1h4vbb
IBmfy0YUyMJZRfmfrSembzRNiHdp9K4CjHfg+lGhC6tbAPzqYojluefghoHIxo+s8SAg2wXBWbY1
YqpcHAp0NG4KNwJw4OIQbJyZKwZid7U9cjUP0kjyeQB7spEOZNLkdUJR5G/X8VxZSoSk+Ffo7gem
etE4Vev3htY0naUG3xH6BUZRm1l50726tNsiIEjfU79fqY2Mr8gWj5Les4J35bTalbNzp3trhkw/
n0mSY+6Y63CYogGiL/oOiCmG6tblQ7dhSwQ2xpM/ms3hdOIwlQU8d4f+ktCC2l/Nv5+S/oWFyG3b
TAfHCuo7q1T5Gm/1+nzcAoojSeAcUzqs7/RXoZ1yAxl88HtZ625QYa6bjRLG4TJvvSwp59i7bpE0
7/CS4BOH4bK36RTkXcRZyKLCplJx20njsr4gn1KEZoYAjOxlMGpYY96PWhMTEP3fhc3+6HPlI5r3
S/xpIPADuPBWEvI4f7DX+G/yHxWxxsGc+q/2G9CESnfGmmLnuQrq8O20xnhj3HRZZgqWxjSm3O+u
FHcXCHj/q/LVh2aeDeky/QZlegLSrS4WaRUJ6GoUr4wFQagIaoZuAF1whnvu9h8PJWMfKwdRuSOU
jXVlySskhr6jUMmcKk8XyXEi70ss6akOjvw33AOUKchNw8tovOiI+GNsYToL+0Hph25WWF9XwR6Q
DZ8rmAqNGqbTVcfHnSbQh/9uxI3dB0jTtPkZWpmns4AH8hVYc5Y4hAKxgZytzKI3E4w1e7wAfHUn
lWsqgfD76FbUdA4HZ1j4jRj0imXXNYQ7ya2i3A9Dpvn3mgJet2IG2VaFIfasFysdcBRhzGjBtonl
3ZeuN6dp2FCc1Ciio4omzbZFAcCLKMW+apvEl4cHkqCG+lP9Ob70yxCGJOIl+Bq9ievDQ5cZzx7I
2yZoDW3vzztd0rMgi/6OkDys0wXDThA8c17+GB4AFCCcTryiCpCtG08Ga72UdE6JX4hhl1+3irTM
ky1o2yaMtOYMXKL7sMHgPRJzaNb0WFt+g8ovAZIXkcNjd9pbPJ1t1CGorODCgCUGJY+kLOo1CZ76
cG06SE+h4f/3uOPQtRvPqTQUzJnJUA2eCVKdybEDG5OKKI99ZyDbIpPctHFuvAewzslfjmnCHbxV
WegsEgEBdE53v6t14EP1MrD3ZrAt8ax2NI70naB5+r4t5aPVoBkXK02Fb3/kDcks9jZLghIXTFtT
LZCjVkDmUtiSR+LhhkjaCb0YdwwyVLUnAyLZLbW2oIjlZ2OglWZXNWtcBCkMbqTklwjbepM+rXKc
+WVOUwthq8924dFTy6jFDYSsnYYyqVqweOlIbnZa9LQIEis0Y+7q0ooNkkpF/hwMm3W9uFKmv0gW
8cznOgaoUyidQ9lNclpn6b6Ms96S7JBR4+fyb4irlbTsy6zBYfu2NPRyeqtZP4yaL7mwPfrGI6UU
MWMUrrnI12iHBw4TWY+n40ICkHdga13W2JkcRjOdBCklSGGJvfe5XV0BZ1QJ4ZEZSxjY2aSDhi5w
8IfEtCDi5Z7uI+yFi3iUPxPF6RzXz4tcphU1xyhz1k/rih/suRod90dDLyBf38kSJ2GRoxlWfmeC
ts382PoWROhEp6YxJ1q4ddICJ3UaXt6HtTVmj4dbw9TFG1tPFC9HWCwVqW+oVmd+dxe3ATmIdn6I
3lN+JNEkvFa5mqdvSbOXXbduoRyxoUbY9lKj2r6ErvDNqMuKgIWBM+MvSCZaV8kcdSbCFrrl4wiS
t7uHant04gwzp8hxZ/p8JiBZYw4DHzjdMULb3fXMGaVX+UkCT+q+uFesJSGyn5ouhdCoSNzcgCst
SFeDAuOl8FeNesOhBd6nRAo6O3Fb/2y7ikHIaUxjs934k3/NpdGnfCZeZ+OOCpbDidlgyzplpFxk
OVCWDt7wIwQJS8h1c/CM6hUWRNQitLFv/DW9xm5p/o2c+s5jQKh+5Y3G/OmkwCD5xSb+EQm7JIWt
rJRx5DdnWMR2qh6ss33UDAnKx0AQXa7NhBdL42NijtOQFfJosuRDWDLRPLuDJzCHsaeowQbz3u9v
chDV/X6vdCM1BYcq86wlbxfIWuZ2TQGpjP4SPg/wo7MILH0LaFFgWdawh+MubDv9kWjHEiWWPkT/
lkJtXaFuGPFt97GaEbUILD5glqyP+Km+zBL9UuFGA5OXCYaEMFFv//hmiOzN3IIUAMY6rg83sqIc
tXxSfd5hrBelcEYKyFDkwFRa0xmBM4oLDcQftVk7FXrvEx1ZzAcXRz/VXXYO/CDdifjWvEsS2Mvv
2cjXZG3BJP4z2IpQFm3FCiHkCCbVVwOIctk9hSISKTtoLIZeF6oDA0n5BQWjMjGISt+QHM0Se97E
PKffKsG9vepmy9OFGOzqcb1YMMD7jPqbGLZrxmswwDYUoA/IiSC4m5O7eLv8F1BcLcuTXUtsMCtx
QTqyfEG/zmIA5ddB+75GpqE5v41/GNlXBVztCUrGIdQn9nry1gBahT5LK0hs5Q8NAEWxfa24y4yX
x97cF/tIIN4x1v7aWIa3EWw7zoQ7+hdrXBCmL9VT3+bPeAXspBMFro2L0L1FegNDIfwfkjWmYmuP
PLyQxogeE/B2JcOENdKfMH4Wx3pUKvWj4dGCbKZ+bS3aE1KGJ705PkPC8zD+gXYgqVZmX0KF9TOq
jnjyFWd6Herk7i/je4SC4SM59b6PINyvqFA7zj8dn59+q/ICZiAuJ6cG7qXaQ0w+fdVSoSGY6brX
0bbRQcV2tGHWAgcY/2YxGuFm7rJ5NPKCu5BFc+2qrUViSl1B8pVmWBkUZWINmSPIkxCxOtUSK/4C
Y1MMJzeQ0rJhpkpY62wJh7FYfIeFoHc2wmVia7cZbInI8ZEHM0VI3L0KBE4wiEtqSTNpdQoHPvC+
ORozINX07+lD34TJP89SV+J10sHgj31eu2XuLwbkARjZRs37LqHzr//p0+u4N0sUkeQe8O+16/tQ
r4EI5TCFl3U15n1T2nCy+KWKkeaA+P637Jj3/rGqoMqyyL4uKVwyYvpCNUfRAtrsVDaAyp680OdR
XaNeuC9dsUvW+hpi/81sgWigfWuMTLgVDyR0Dz8VYk9O6nMi9NldwSa/D0ZHjlYwwSGi0cMttdRJ
D1Q0ew9yGaphTUJ6TdP8eTRAXL1lb0kShV2hWNALHX4N514uKHNEU79sTZvRmSJvHb1OPxhSu8iu
MVRBPZCrXdGBFyccOBSh9V9LYaFfC0MR1rE7x95M8Xlk8yuoRdiWkKgpqmxcfNPHc9aKgI+3WJIP
+a0KCflNAi1xLPl8hcUuhSH5YisXOi8jA3g1UCC6wAlYCFbGeT389yJgnrO6i3Et6hyes1aa6PAK
VISqwDr0akQAmIF4yvgQEW+tN+lvNylj4WVyjheTp6cn3Dc9aEWISCBBZpTr169KZpJYfhbz906z
IK0Pk6hlNv3Qi/rjoP5E0mmtc6xxZ7BMzat4POD3hNqIPGBTznLSrHjfQR+bH2W7fAYZ087R3/ef
lrFeb+kT9eiWfEbLiWMbyqgrJtn8PAYv3H0xqcjDEtzOM9a491KNpzc4mLJ6+zyheVY7UwMli22S
BVPhIJOiwajCSUgbMEA6whOFmFKNVBBm18oukF17erBnhSOoYbmlPA0svTaw/QL6R+EuNTMlESXE
P/dsXoiR9IBELWBraeNDF5jtywZrI75DQD/jNIduk0j1Ldi4UeGwZejmImA2s9LrfMCFu05nrjUz
SVJ7q3htlYFCzaK5ZxL/LiVreBDU8NCZiQhmPgNo6rstGQvvCg1ErYx0BiGKCA3eI1GJreLZG2Te
xWEHzWuX6w4eaH8f9yY9cdq0uFaLM4EweEwY7a1xQMf+VrE9QZXdthaKPRL/1ZPUGXOOqp4HufPK
twuGXH9OqxBe082pYmMjc5zPsTzscM5LxorXPfy9xBL2AuoQnBBCrnLSrpA1+7IUXY8qWN9XCwBS
B/wVhGyqV7x6cVLeAVyg6uApe6koStDVImm7R6/WVqCwJE4zXw8+6ABKYRIDMakpen2ecqEUVjSy
ph+2oOVdLsMHpgeWGndb9xG75ZnDNdCPFJUo1tW4BA8aGDUFA6wM4ktXjxwy0SG/GLCpDZJ1okni
ZwBo8jtoEoo1nuo2kb7trgPFuCHxtmgcb2DdswpmOCtiNOZOFocMnhJU5XmnaeSxLtuh4ypIT6RH
iV0Y2MnMjMQq6EqAzUhMydDzrmkGTJJmL0PclvH+/BxUASlUJiBgxhspTo14/VJoTvf9C168UcEe
2QXhv+4p5ZVGWw7qNWbo8nd/ATtEfe5W5zOAvB53/9puL0Mhygag2GPMnBSZs8Q9MLMtrGTbau7p
e6OPmbe4u2h4g5p80xVKOOAJJRqxHxKV35U+kjB9QBOGNKBOyS3EBUQCBcc8OCtMePJLxII9GdBh
PrqagY+0njK5ua6TgpnE6CR8Wchpohse47YKhubQm0m43XLF/vu0FL6C2fpyb2LN6LuDiNJjftDd
toWsNlSdOEMDZHs6F+xnfsxHp7lfIJAUyQFwDkX4wlxwm+XuQuZ+e5GmagpjQ88iN0UaXLBzI7NK
cOIyEmaO/R3c9aGaV63LXtuBFLpmKBZ8vD7Gak6b6dbSgXIcp6uuLyTGBCIxyXWvpre1gNLP0hd+
hrBCiyNtAVHHNJtNAyHrlsBZteco1RT4lJnf0112L0zCSl8qM8nUqqtZjnKRKuSB7epNWipQyASp
GSI6NFe0pCbvN7hp/QW8fZ4Um9TmUPTHuwwPKYTYz/9+rol/p5AvMkt1Rpm/a9b4vqXbDeL5+c0P
xRGMgU3JX6d0iDnh+HFHJRsT4/kYXsTaWfx8CMVDKaFtCNqq2nhVVsWC4VxKHms7CnYc2tr0CDie
YJFGhiLao4qnyHnDAPPLnrXHZj4fh3iW0Q6QAof/j1X4mpfPhTFsGUH3liLOiczQAEIp0/C88H6T
naVr3vGxco2vLtb7SMdTvE86PVB2eN5z6heFCRc1SCt9BTm4mf2A2Po4W9dM1Q2+/QYkqtsSgQhP
kVnb6OwCA12dQJGQ3DcvBv2FwO/4hlsT1JCXfgXWk7nEMGA4yyGMPPaafyUCKR5MNcQPRa4T9Anf
+yNcNMqApfGqtEwoC8FiGA/AqOvvzQhweWCSSmR3jI9TDAckvZP+3sqsXLYy+lhwTfJq/lHmKM9M
Hqh87cumDDX5xLIleo99MZsu/M6klxE377DOrEu1je+kc4hYyyobiP0NyXR11T2tBcLNq56ktpWm
ELPUd7r4gyNIfGpNrIU1gsGP77sB4NBFlBcRNhPcWvmPovmfuUtn793JdLurMoDWtUJmeuvh1RSS
5uQSrMZXytdYIEVJqdZ5TGdTM8LXbCv2m5cV2pbaSv/e122+EqtjkwkzMIIzw0QV//+x5NFHYsPv
pQc1DSRI0TNHuepE8WGu1+/ZDgPmRTP95PJOFiwRza4IbRAe3xdBzAkZn2mkoLYN9PPLbawhbHUi
VFD/xt0osde38KFYvrOf+M6A4UjMkP1lZIMTaw29swJft4xFpnOkv/MTkYkQqbOd5N9ZFkQhYW+x
2BGt1cB5urnKtL1/i5SpHTVJwPyUOCyc9NJvkgbfeSZk5Pn4zjkrlgLWTm43VxaAozLKeT4NjMRH
EzfxlLNoaDTeRDsEg2EsEUeHWGZGUcNcFgzv5/f740PmA5D+qGbE+cIUMesva4+bsrjYHC3xT7z4
Wa0AnpyNpMXoJAMccqFM0I4oLLwvjLaeeh88+RnyNY9VP6qBNSghDdNB5BcgupkBIetZWljpn58/
abtYtELo8bsfpHy03STh8AG+nJ+h/Cu9MKqWD3khvVwwvd2++Ht3LBxpwk3yQyp18AteK7fF+1iB
uvh3gqCgBb1xqk7GDs2Gt8hbNzxhi2IUD168oRBFVCWipDK2BGbiqLsFx/qm0/VlOUGv3+nXZGUS
K7Hxl8DKOPepz0pdWAzRPmtQ/PyalICrax8VNQliNOpBOq/SDxqskxze2+G6tj7pn4VrkclKifyX
ATlBwZY7syfU+lA74naAb26lUK48STPu1Uo86Uc1ceyZMKKk+0RwzHDx3UK8Ce6BAHRcuFkUD28i
aOSKpnaGRugSAO6fiAhINS8RbLufe7khjmOKuHpTvzxL02B+xKRIvmLL+Iuuu6MvIE2XIsgCOK7k
MAQGmE4h9twhOkqb7KIaxg17I0C8BbbpULJKY5uHnZ/WCEWOQf36yF+Q6x9KBHlgiioI/97FWCeo
3S0MffNan04QNQ9A/KJ87zlfT3pCyDUPWe4zLiYtgUns4g/gnZdwunBOQIgCh5X4didpnQ2vgqw+
66dAVE6aflp7bZRwQrbA6LD8FoYe70a/zxGh8B+y6dA6PUH/1Byn+1VQukK++MWryo96CIM16FMW
uKxh23h7Cg3XR6wUoVZyn04tMuP2oZV3EWjwcO3E8gspnUk6n+ltad22legsfYGCUFc1GPpEel55
tSKYLPsMasiGedZty++ZYeqGnCVabDukziyQkn0HHaonoEOS4mpm5oItzr7Sz9H8XAts9Eizug0F
eGnVynKpTV+Daii9z2lQgndgoqF/IXsCN4IMdA2uwcqQS0m3rxt7ck/9Ow3HCRv/RSGEu0JfhKto
B6v2QQn7B8xukDuj+pVFNKCsrlNELbA7cc1CysZm/PlFGkIP6KTMhgOhR932oYraz5WBZHl2x9IR
G3XqTF4ULeVLNnO7Dsaw0qJIZpbAt6i3WWjFbffXs6Fp4PVnxOpNnsCdd22HcdhUUkD8PXIzKHaO
/0GZLzQPti9vz/KKdhPqEpTTitBOQJpFSfAMssO1eqDadtfFCgMrJx/Hbb8Q1wKc+TbtT6rjd0L1
Ws4XicAnxzyXd+xspiLY/vSSTHp3E+ZX/rUQLv2fBvwXT+4zDyIaavONd8vLH1Gd/6pkALQp+yKk
l6gSpx8TbCXkk5cJdZAXQ7d5T7HgY4V068odmkSio3BjUihGHvaHsq7Py4J0jdTP8ojuTrpJam43
uhnEBVpXqibKJ9Cj/dymnHZCQIOE0Wv9qT3jdiPqG482BTHMHLzvE4TPetamLh5OCnxV+2RysC+o
cwli+IDpdMxoWqOK0pJWWzzWuEAyt95aqTn5RnLJW4bi0Jn4wdTI89iY7v76rOhW9P6rJsCsqUze
LQ16XH5nrm4br2StJcVtKs3rCiaRFcHIVDXRsCYZn+xvrDtNNmQUiekSEQTMdmTAlSg0cFkhcOJ6
ruvsiZAuvC82whaAnD94kDEhi6tkKQLe/ku2Vmextv1e+I2qdXPOh77SvuNzrVUFfpN/o4twDFct
v9cSsLNEo8MBng/qOsOwZZlbt9XQPYVcBxx3TUuolqLH9xWdAFHYi6BKGjKHNiU/ADhf2HWHLbYz
uh2+wpvxbk/SVCwOnWg7IOjklf0e+EcrNayujcrY4w9kbg0xiKTvtWBGN2qtVHogZhW6M8V9ESLC
12aN7RAHgWYIktTF3lJc+FZMI2ALZ36TPlJXTTN5pGwsBwV/mpyX7vAIObFD8Ku7WbVPt/0dl8qd
qGVvW61JMVngMnudN305eILWwO9ewKMOPuNN+BZ+TvYchYZej+T17L9SY9UXe7ldaTHXENhUqKfe
q70hMeDWSEtngyYFxF44U/7ZdBpNhtUXB6k3xkgaiaXZMVPoLhGewqqsXtikrm4iz5K1C69iwHFW
O0y2kjyfklLzUdHq5AeIsZ4YIXkA5zdd6J8QkZ/4m7AoIs87zx3xW58pJdV1Ia6iJhA7wJI+ljwk
oWBMTgdpqebXJQsZWJrrcEc8mo7/UZO1okvCIBKI9W6h1tJ5fZan8BHivQCUgHULAAc+MTbgIFwT
Qzj0WAjchjuK4e7PwxXvrcFPVE/dFotvbvLrpJxmBguVrJHOe7ekyklfkHc6Y8zPjfH+ggA1YWYk
CBj5HsfuOq/cYjj1xKEcUmZODAG39oYrI9yPY1buOfBhPpy33qtehO5+qcf/zDku/ysAH9hM92f1
NWElwTWsGAgJjIAuAX08Xs9TbqEre9FNHd0vJmMMYsb7D7PZNG2A8ZxXIZsJa34oHw8ywXnxOfQo
q1NdghOzO64KfV2zzFxiQhn5PbU7FXQM0si51WR+YluRhqcHkWzXy35BCH8b2BhcqPGopcK+sAFO
arLrN0KBhonMkZpwGCIbuwkBIRvVP5Pgkqb+bRwfk+dMlKvDEi4x82nQZ5Be297WObQtRNBtyQ7I
h2Iraahho4ZkNfG1hQ/QerzsX871H6ERN5qNYFoeI0urYErPcD+7qkPhK2Kcp8uzxt6xwrsXwVDd
2zBQXKMZZlb4koQXntUzc/sJicGr3TGNsEgsK5tOBNcApCK6tAzzKZvetUwJP/o4Vqe0WtUZgQco
JjneM54+AgBNTz+KG88ijg9C5gex6dPHOjT8k5LoyCz0oX+E7FndOE4ET6z0s4LB8tTOosq/dYlX
Y+4LxbgFtiYxtEziD/oiHeibXqjuKnz/+QWaMac7BDxmLf/Aiwvp0XASA96vhSRvJ7almYPaLpe3
uH7HM5xzeS2ABNIwPd/F2tvaINP2GUQUfgJzZff/wBk4dq5c428tVWbcmMXtus6ru5MNHQ08nY5h
KUHfUkP6Wx1DqYkZ/SYC/vz76hQEkPyHMJdL+/TpPdC8FbhIV/VIXe147bhDOrtAdJSF7sH1lE43
4zNMjdOoRs3N0TKePoVB3yx5kosL9K8jPkbbsM3PeJJkXuEyv29CkyJH5uM+s3yI20wrp1nHVfWN
nLYAaup+azJK6CDB7HyI40/JAyVjcDVtDa9XB3br+JHxptraIHmCOI/H/8xGeXy7hxi8XoQnEraT
pEtnnLBxXGq1kkmd07JLdpkqAXBBKK2YV2ntkRXSL9QfTcpYTN0aZeVQzzSyCTHYpY2wGOMeNMUn
4Yfm1PiVADiIVt9JnJ0RTCL7AzvhIbr1wmjmy0UY+4P1HpD36f3KPuVHLrsANZuWpwWiFk7pLUCr
m/MU1Iu/xv9YJdsBzlTRpxf698YVcYUeshbe82XH1BuOjOON5s1ca9F/1KOWHdtDxcdxwtqD5L2k
9gY6mDnhybtLLaTy+2vBODDPWJhMVwC4lmUkho921ElFIxDex8bSbsqLQaHGSZQsv562BKZ8CwZJ
AVujcfjm2tbTr68vXMA+BYZ5g+LC6HFNdjHnreJBo9pFiBov7EiYoHQ2qb1dZQymGeWbiy3V5L6R
7629D/mkuaojuOfFo5l3t+ZTDCZ3zkV8FGK9RKmi4wa3hnwc3tEdU4ZcN0KHKykV7HwuT8DO4Y6k
+o9Trl6q6YaiDDh9zNTsVl+27J+s42dbwlrneZ/DObLS86cUVEdA59oGg6G5mGYXXIlgLdmsR3D2
Vz3PmRK0L/x3ZE90lDdetDVqdZ/vFwOUFA0jsK6gSp1qcjN0Um86aRhZzn/RkLQDeY/f/zz0P7gT
kDWJ5SVMVF5Tjoy937K9YCplEmNt/hu+Jc/7FlktfC3eMAW67bt5Apr3fYKCobCpGuLMRdl+bnh4
+8QnftrLLMlmZDMCcOKsQNhsFB2RgMMiUTkDGZQK9Cc9/B9HISxwP9tE0t56Q+efsM5tVoeOsnJm
MmK6Dlah4rdKUJZfFwp7CCgi9Wd/7GSafAANe/PODkdmsRAj+xdBY0Zqz+vEHcG8bNlRUIyZmRX7
WFGtGGZxBoWAfzqPr2+CoV9k+7s/ym7XaLU7ja9xk5YzDDHaU2VJAZsmbvldhM5bFfVE/apXQfP0
INf4qDFc21PZsFCUXCMxcKYDylVePKSzDO9MNVqf37660GY0+Gz+3K4Tuit5a+fASD2o3oY4WOuv
9eQ5w63Iy8UomTJqVIpdhxm78QBaP7C239X6KoiajneQLbGAETAdiv1xz5/KrLnJYJYsN0u6vW4o
8FDVqPJ81NAdjDAXzBx4B0g0YKyz0RoYashGsO9Tqmw6pBeWFsJx8v2iVHjavEqw2XZoUvsjO14f
ksGGqPu5MYeraQjyHGLF/JVlEuDDgf/VJ7obZHpeaGSLpmQx7HA9aBLQpKFFNd/sYbpQ8Qgv8GqA
BB/mGtfrhW4TEh4pBGmoZPHM5NKyQHGm15UWWkwKn5r6fkrcPnl7jyEM4GqdW8R1W6sMmO8KNasr
+yANppK3QG5BaQS5FsqRp4oybca3CLbS4GX4a1zk5N8dKHyPV3tYnJvVsxCcJYN4HJ8DN+JhjJy8
UsnFbg47Lx8sajzEwwbKPFiP+vsJpDYrDDmx/OznQMbxREkUqR7ft6KTAsDdH7je0ki4YQbSTTFM
GRJ1kcWmpZTY88giGq+U/RXEOQlc1vGqxxjaOTZjsuwfCh7U5mFFFeRa1bucmNGEpS0gh68YYNj7
CHARrutp7m722cAOKKlyZDWEw/mvOAqba4TTbhKHT/oP6LmIgynnRUE8h36F2oPQPxl8G30FghWk
iaphfX5At4rQ0ju5kP756DjLaHc6g04sgi5+me1B0XIszd1x18uiMnUNk90kCDsBT6Lo9vTshokB
hiiu3/z0Hq/+AoTG6/MDB+1oLp5rucqhqlQiyc/kGABP0RBBtuT7oDtljxRrZJKv34MrwwApTlTI
7IZfqhZM0nRLYieXrPJk0hQarRTz3hfFx9N51XAJ88/YejwtHtzvv5zcnRyrtHnEP3LOH+RyE3f7
McSUUE88QXTsJegVxmJca1yBiRQBWUEHdwhIxCyOe2PKXiUUrJw+HvuyTQGftcnwUkrS+zjfizg5
kFLTnCaiUklg7aLIEO4L8rzl57LRtYP/X6H8YbOIuDmtOsNHTOuswCRzEKkEhiwsUNMtcoggLSwO
eL8Ll+zC+IgX6t1Xoe+sLdD6HlJKT+cYmkv1MX6VATseeDo4l5DYaER4W5umKNajEW2ULIPr3gM1
0qXEbH8OoommppqK6dBvhGKTYLLWpFFMQ0yDANSX3YV5cVhGBrXGX5QiNF8MVfvnr+yO0HQnfPuI
2NQZJc7j+7K788p6NCiqAf66/TBZG4Wd6t8LRS/tgWn8FY+DFnowxE4uRJc9cnhwZ67A3vPqvHL2
GPawdWmkQNdenZEqLeXsIfvv1dvCf2KVGkfUJRLBDcf3ZMLDvSaENrH5fto729OKQy7jbfsPym03
PvTgkslDkKUDSjlMVhDhNSmu/oe7KdPOdUa2C7r8JZhH5jiR4Eqi86c90zYwUT5rg/RMQQQcgaDt
H24KmW8J3kA7G2jaVwCdjn8ypV4fZF2QsMkn74q8Q+kHU4r/Ve1oqZCn6xC5LpDJcgqb/sVfJamq
+KJEquHnLQYFHvmOl8O+bh3vqfwPn18ky0GrPq+ZLss+MhBkW2xRIudWU5o+IHNOFrO6u1lA7L23
SL+Jytx3PjWNpCx1o/A5zCRtT2ipddyDTRv+0IZI0d0SwCx/h4gZg0KCjDvRPdSWRgykcDufVVQB
ldJhVBKKXa7kaoOtflh8simf9TF+Ea4C0Esvez5naye9QKZTf8pS977WdzjTfqqRZkzTPw6wH0dg
rII8eM7lRZvXrCtmzXfn3dybnBRpkc7dcfEbdmWWUzt/uRpyR/kcNYPjckcO4GEjQLkD8VGsStMI
ETttnTPYT54Wc4XNbbcndPvRdmRw9da3X2wE3iNQBZ8wmymoMw3MQNXur4aH++kGIfwck1cX7GBt
anGbEQs0DfdFOZzT/KZ1khCjeI632DXKomf8KhFYToWDSt0EjDkPHcYc7e2JQomJ1X3/ZNXWBCWt
/+uX//CUFW1xZ5+LUGNjUZPklmN27/X4cE4Rn6TQoAL9k6Ozuno/BA6Lgi/Wfoq4Ek+RHeq9gzJ1
bU9Weoh9fkqz9F4CxUwyBjHJ+AAUb2DKPPSGQxZyEWpO5692z0zf2HhLLxIe9a/DvXgcTSbb+28s
0Ipet2kMSZPMgXnN2a0BOeY6cFdiNzW2apPBauEES4HUZaYessyiZDdGoYafxnYs4iKLW0xSKDfB
7uaSnQGblzYXz2uSE+ktLHBpo/do6Kpgu6rB/6ZCxF2/tAY4n/9Qo3bWaxCwte7FhamAR6bwyiNc
UBc4t7i0vkh6BOdSSM1NMeSf53VAJ2YochnQjMlHdEWjz6Wb3xh+jsgwxlTZuzUDaHHm1Np1VGC6
HTPTb5BvqUNvoI+GgJmJPouwZqWm2w13/jHxbpeg4xDnNfNe05Wk7g0WIeBqWOD6W6R7CVrf5qy+
BkX2kn9mi26cTBpJoNetNdmfo3u6RPnV+D1q0vsHKiBMTJsc846lZQnUgr6ETFnwpjjSjG9mcuFv
VMHlRaSvSCLTVo17kE1YEjZsPNF1NCAHoKiH1UQCLATA+zbizTdRkMoWtMbHNXvEfZ2L5OLO98EQ
nODRRfuD/0zF7e709CSYKHSMAl1++S3muwv/Yu/6lUhHuD1CRaLrXuYDHpKDTpfZcG2vMG+iO84d
D/vWBUw5dNoWw8m+1j+W6EWfSiMHB+37rZdhY2WcZKndHQKuubRDY3icbi1ZBQds1u2FLJNu47P3
0nwd30OUtKo7UqT/wQuoxs+Yc3n9EkN9OvWHGI2Y3yzsembEeAwP0LD0twAsg1E5eDjOAwnd4FeN
hQCY4JGM2o//3C4LjV/XoH+Cm70tXbc8rOMB2mzVaEYIZ+vHo0daNMcPwaUbt8WPlWG2kHwIC/Pu
HJDKA/q2+YoAWHBDGGnTRwdd/7xIa6AtIBztN+96CM26wsq4RMtaCsc/Nw7xIwR5LX2qN0KTGkIY
VUtVmBSVah7aCkgnykiGh6nktILHX7u4FExBDY0+K9XzN7LHwP4+kLlpjALv8GG/HeTg+wPfmAsO
rJGhOmvJuF3jpRtdH4HjzRJPSUYmfoumNUIwXgO8m4kWK4my7tMFyTcpSe6bLX8vgIRx360EDEST
h+wYxnHwv2aISTRysnJ9hDba2J6gKyGjj8648TcFKOHS5OllcYs14JNMTg9KV6cEIRPabs3rgZhw
eT12/6B1/SMqyCxIxd1pUZanKWBtuiAtU6jk3HVI0GriioMmD80L6TaoW1nbHNNT+JcrmgNKwinp
mFCGV6I/HNSkiMJjQWWIpBoQj6c5xMgFHfy4SHt4Pb9P7YIUobPV+VErPimaUF5dYBz8lbdukp4r
h4t7kAmW96LnZTshEUgeIVJdmkIJhaqik4EPrZWoo0CpVa52TQctsdEP6QGEw0go0AJY3Gb3o+lz
vaS/+JqLrgZAStSNqKi80Fj652P2tMUUb4HypCISLGyggMyNz3CvbNTpC3maTijU0GQHGzEqW67H
+phh5j+Xk9ldBI/HdN86mO/gPA23gfOnOPFIuLQ1GStp8eNK2MA9l7qam6HWzgdXhAgkd/CXPoCh
WCKBy2JAtWh2QCe7Vlq6KD+dc7U1aAiwma0Aarbn2/sXU+Ilk1rZX8ySmm+aIra92RdbWt/CYBix
M0L8PN80n++hhRc3Mm/7Orkx1/pCpq4TgMMP4aDJFh6AmtGkUA2YBqh34/Xs7ee7aHtPM78WWVaa
2va0MUllVYXrR+uUbkmRIPDrPIWilmcJh7HSidky7EKVa9EY75X+nXtx3Om7EAzdSuKPL4GrDVlQ
8fPc8Ww2r/E4rcA5Q+ByGcbLcwP3uoc8EzuHH3NN3HrTTMrYHzuA2aNu2pNJwjkv+E2T7iESqxs8
LSx1b7cIW4iT+UlK+2pRGgxxmjbJGl31QTv/6TqImhLYCDQkSrGoWC1GSR59sWq2T+GXAlkXV0oq
VdMfpumtWLP1M0KBQs33hxCVghLlkR1iJJmwvTRHgyoEQs8rp3H8fzzdb5nbroSbdWcrTt99W/eg
56TFCgC9kna8oB6guPP6Grp0i8jZm6oVZ41tnFRIQUdS88sdWPsBlpCXDT9DKQa/mMPlEjW5/d1C
aThk3JXwQHBPytc+pBdjMU4R9HV/P8u+Eq6AMveKK6/xOOGUTGXuh7o/gR4OBobQowmJC+fwvZUJ
Xohr+4jT/XczjC4mPW9fBwvSISBjk1tpzEHA8a71TzzO51II1wUcpEkoICQMGFP3ZGe1AmSqWsz2
vlQeV/owYjb3LCJxf/igQ9CTAZYzTkbMhM/YRaUCOlscj5EshSBfF/2V7GIyBtKluKX8tcXn1jr7
ZKxIrG3k2cPChofZmlHlNKyYk2IPoQEbCMOWwp/lLau2NZ4LfW80jxMDdIU7I/fnqGbAPoKmB2Hw
HmB6JXf+ryzrv+F93CkSfnMGwNV3o52MTe30OAfpNBpyqI+6yEKe91iVi7tpidISiVBqY/5jnA+j
K+ExbUgKmWEMDBcAqq4n2Jhy1DUuX1SfAM+5K6qJVcAa8WyickZHhbIr8X0AAkkgr8OGlLO7cB95
88OJKyPziS/oiy6OWpdvzVaJdoUAaUbLLBmSAuAf3oyGa6NDXe+KaVjgYSL3O4063tLKwAuCfJIi
xPl7cQl7HyNnWZlidODw7RPSbZYyTf8fQtf8/1eju9XKl6dtj2nMcN842cZerVLPun7nZR3Z9oOi
dpaoMH2qWdYDtRB9I1Y+H5O87rsXSmLvIpNYagWIb1A3FnE+vl4q4fC5FH+hve7EznHVhuVSCil9
EmCis1c+MUyX1BLLgaFwUABwq98D1I4sD2pYsoG4iXH41VTMEUI762uUkSegDKR/LxAvPrcpD94H
nYb9maEE5f8c0daQIeg82wMIahNpq63PyGybAEpjhdGGSfItoxzGQklg0KKImxbzNeX84tpodaRb
zZcGn4EuNH/MpnOkxi/r5wwEmcbrbMIkpFLUxNE18sYRHKea7ibChPNBXU0HLAUouJe0tZX9mG8H
z2e4oVBT9dB26X1HYIPYrewHtMJ50c+N0m7wYw7jNoFi//QXHgLsQ8yGxSBTWFMZ4YyBbhjuajcN
Eq9G9OUtn9u6Pqmb2DsQUihBGyyYeC47qmZZGSpT15cYhO+N9XTdLyqb9Wh6f3RK6Z/U2xYULKuF
Sn0LGlWv/aoHlrDVekgpuaRN/SIgigkwItrHzij3+u0T11pY0FW2SoL0iuvngsEel5gQ5hNSo4JX
mVPjJvyxjU218lbLIGY7Dv8sDIPIDDihdlhOA/yEfGEQ9oZQeQYEBsRzKeRu+1pvquJH8UKXCXiG
zvWqw4qqJf+K4Japll0pb6+FCO116wsDtZINosCyWz3GbJS0Z4qQ91pDTDn/L1Z+AGHYpXigfHmQ
RCNAaNTJzxElFb5bLFn5sIUA5g303DFKNGjdyiaqx0duafiV2AcTRkhzlioZgWlxistzvMj6JG71
n+pFQdW25M7K7n0kC4maT+Kaml3triqFarYSohe6sEwDjkt71gVhHPIVhM3QT3S+H/VIQt1vMH6I
6QVwJjq+qd68f+swz0W+i9h8zrTv2hFtXZwxQkXN+dF8Chbaqw3OfI2e/n/GOUQvZcSKc6P/2Uhg
dH6v/T+b1TIS20vAWSx2vwrxjNxMMN2X6e/oChMqXwQG4kl/FwDPTjJTChqUcx3Mc30f/qU48L6E
faceGL0S9CmYnuiJsIdWmBPnPckVbHFyN+Nhf4cdjbXrCSJClc9tH7yox6/Zx9YV+mFeBT/ODRx8
i+eYq7zoplmNMEtML8YgtOtN7ELO06tHf/gunInG404tyWaLaqRT+2vl8JgGMqbRyYvHvTxTW8qm
6b0e+0JSiY0tgnjw14E1QIb+s9JBSKfzG8tKnq6rQOniS0UCizxIjLz1MQ/+5OPvJSOtI1U1YMw8
P8bTyRYmf2VsgW2lrpi+/qNqHKb+5mOMZMEDQdeD/phk9h1gzOPsAIh78e9eyWpjaWaewqWXnkyp
upqBLPfUQq3TXav/Ya+16wvyfO3oBOYdv8dbRM1J+DovdPwNh11c8DDpYkIU+EdQrKW3QJNWy+Sa
75dFe02hm2Hxyyb3DSTU1cq3qHPkVfsYZcGDgmLqz+cIloXWDQxY978fJizCq9wbBbdl4jToSZog
xkWHxP73v0KtixRw7odIcB5V58hky9At5Uf+NfxggyB2tNa+AWPSBzZPVUdip++IGWMOomckhALu
coVQDfoSesNomCzCYhjoUu0GZSObA8H5dS6f1DyPqR/ejLBWVUk1It8+JZTYpqQlrVTK5jBdDhQU
3bSfCAPlEVqn5UCDEh6gvoaMoupNMkNiLMcySML5t44JEqrvprk0HR075cgv2J/vAG2UEMO4GeNe
viEeE/UucBVy7TQyNhE34znXEBaIAukuKbNCf355mZR9oyngb10Aq8vOE2Pdr+I8oZy7beP/hN8u
Lfp1kpQK+OTa8fmF8WEbyrTacZJ7Zk+AZp8wWfYDvWzJimSICNOt3+C1mEGnnBp8FVvZFCvgDNQK
gFYV++U5js9eMjPZhONoV/k89952pkwhdUIKk5OLDyaxHv+nrHrRy2J9EBhMTtBDP5Gc1xjA04mL
9pHyQmmov7Gi04bcy/5z4qLlBjJrDXWWOS035xgXIeN30mK46FQll32sDgrNQ96Lm6Dzriv/NFxI
bH/RiPitdGt/bPWopTNMc9zlojPaWrA/clXk287W5mSMjL8Xw5HWhazrehvI++9SyXP8BGG64oUZ
5gmT53JD1HDR3R+uYyiwa7++oIptyBzjaBX2DzRRLt/FFmMO0z3ZyYzKLqa0blkVUFcACWctvS+v
7oePUrE6oOg/9OMlhhZAroZlzuvkWhnUUl3Yp1lSkhss4FEfxopqtGZ95T7LxN07CuJAR9xPTxfK
gUZ+mZnPX6E0PMZzuamAUBUh+wb3P57V6p4KNIuDPejFHXGsH2zlL0MX99bnpQBqgCSB0abLFkUL
jLkXva5x1G4U/aSdbUG+DKNOqhqeTf3H40E0b62kwmfAJggdmJRuL3tVw+k4DCqvilF0lT3mQogb
bqNPEHvq3uml59Z+O0GK4tEWBB4Bj5r7hclgR/dI97wjOS8VP8YVhqdr3dmkBu80o2E7xcCyw6ks
OQ8LN5CoqNWjFtCLRouPWawSEiuTFUbeYiimpHTy81Olr/vxrS5YaNkMCCPfwEEkOp9yGw91hAvc
GxC3wzgEjoLbQ4Zqo1JuO1bMhH07ygPztLZe81CIX0dLPmOAn0HmsgWruUC0E400Qh3BKAUMjX2q
fK8yYh5UiMKtWFakDInSM4AotPDiIP9Duh6oLfAhdgop4urMvOEk0YB4XKruk1NlP37+WDlWh0GE
qO5Ap9V6L8UErnmLYRA9rlvyzl6FN1WGWReckb8gxCrSZ0+T4efu0CW71F1EZCId3MY0hagCWtyI
F4kg1t4KnzWY6WrUsggPUA6t0HSNaZTPK2pGw7eL6A2mXfNcLyxMkL9YU8jMgwHWxN6QjfZu5m6e
8BVGEmsG1KXzNUDAdIuU1vvy4YT9NHZpm1TXOI2p5PmB8pDRUIwBgrbsOfsY8SVIjB7d6drWBOeb
sRvDPjfzEqsXQZDKfvjtzGgyraFDBNYeAp42130xAeQOlaHTsrpBwm4McN/VcvCuShRnpQUEEYd1
AnAYc8lIxnG3Fp0uR51L9v+kpB1d75OzzpEIdrhgv5Ul151SovSIgqBOFSMK0JuKCtb8SRbzswlP
2ayivQc+XJAJMk6aBjPRbfN33vHlMCuUQY8FZbRqtHlazce43B/lMtr0PM+GaCc/5mQARjrg/2rs
VcsjtgC3GYf+/590X6BK/PRNt0yN5Bkv8Z2ZWt8LJRwak6QW4HjE7dLNq8m0Ua6IPSdkTi0NlLE8
RgR7mdxRW+Kk4Fa6jaska+3q3mI/1/fMUKTYkkWKA69NWaE9ExrJYwO170Yk4YQLxUykO7iAbDSG
qwzf+o6/E82s8RIpKBdEO5sJldPRnpMFVLRc4gzycqtwT60l5exxMi+eu3w7S+MsMXBjx0WXFKof
ciBsdh1Vl+PoJUmpFrXntJ+Ip61fuwccywkLiSpOS2jbC1JVnbqjMORjLwY+GtA1jgBSFWVANbE6
f+Rr+w5kaFvsXs/gH6OiFXAZ2scDSa2rK467LJQurxSeEG498jb39tQPc9ANNya5O1YwdEToP4Y6
A50Cri7ZWFEfVymaCShs9ilbO8WtS631iZo+/8vUajMSL41ompHbvuGBRShe4DCCN+hlAaIYXzdw
r4AIi8S+m6Axv2Cc8U9liEx+WLTvc+5qYrk0kVlHuuF4RFW/uhxvGLUs5kpDes/+NFEilfSTA7/C
GnDcl/pJgpDVDfHT9l2rQtAqGynaH4WAXWaPgGBRAFl4DEZR+rM7DFJCn3Xl/BGdLkNsPAaVugXg
9XzdkmYJPZeWcXT65K0Tv30yDBM/Vwg7cSSp1DXVeyxXLARH+WYirRLd0T5swyikXiiX5OAFTRX4
CMNzfdenWLD/Y8VStkKe9IKm7Q+m/tvVcOzTsH7QmDdm88xFXIKTeGGnRLGQCOxrKfMd0RCnqRt0
VPg9RyNrrvn7J0Fg7KDHe07P8exodBKLn4v/k7DcRySik0bPSaIZ0Jgyr9U8661t5b6Dz4RjMdJP
fs0Xj+0Ag686X0oEEWO3etHMYP82n+GpCvjX26LpywNVsgrRa6AGiJPBH1A2JWO5L5LaP9cFU9QD
hu+bBsyMpxlqb745cJph3UCmYPkWDErOXCRDFpcqyTYDd19hc7+4+CcBq5asZdJGTydMAG9yJtrm
31LmN/LEFi6bQEuFcEsYwGA9JA9pxmh5xzw9FZYCEeY4sgPx5hII8bL5yDY3t5VqTXL1XQaKMoV8
gOT7qKan1pTxgiQIiteRMQoRq2tCL6X47La2MsKR93DfntV2ARxNWdB9DeGa4pBMiAu99YshEs/7
wYCIEs2R+4jQwHCSDt52YbMJco1cz/T1QI+TvtxNWgc15VMlk/15cA6x2dcU7W1biGxGEuXu4IoB
NQ4/e8drnFd7/i9qL18NJPgoljCXpVw1OCPY0ak/FP1RLTKABuvSDN3UbALn2kb4khT4EieVEZIS
CX+IGxJA4IkYshch0Jx9BLLXiRUCiL3uFhCqaqASqIuQH7hyEFvdNhUByluIbchTqHhdVPWobTnI
IsB24thED8W4TiWhyrIEeyd6a+oW2JpWwvfva5GE/OT9VYnz6gJhGyhPTPEn12SI7Tr8RIB0At5p
Yr5pqOYpNLx5RxSK/FBykEvcMRGG/7CF/6t/2h2VFsHc9KT3C0blUWg2yqx5IjO8g5AOYpwNQpz5
+DLQDJx83W0vyIO7q9xpp8u6dhUtFXzar5fjAi/8tqV/XGvugKyiMtbad6zqAgt/bysLY0Rbtt87
fuwzBVbJIzXMS6rwxReYbGg6Y9Bu5sjQm+i6Gu/DdrV+7UIbOadyVKEWiPP9vMLieYh5NIL+Ym1u
5SlOUNGAcIoykHOObOypwHZt2zjRUiAfPp+QIIToWgJNB7JegOmNwr4cpsBimCX2+92IDwGTnDm2
EtO1PawIaMPH9wrqM75uMyRci05ZInYljjXrABDEk83cK/sG0S+LYEP+xoaymkT4ysXzfFsu3lxn
4uEahBZRsVrwgdNlQeQf83sBs07FpasSvb5bBM6vF7k8gMrqBEDo0SDZ2W+Mfv+vSUn8ilX2zH2w
ZOxN9nJfvTIG0C8fSr+Cjha/EB9YANw2I72g+CUJA/pfDt7jNoC8EO+GabjWJboKZdGVI32VxwQf
p7NI9FGcXDxZuI/PFQxJpWCLwRJnGFnvK2UMyujQ3cV3ZUgLI26DTUS2BCJrj3jOcSubJpoMBsxf
lOEW4ieZa92nIHMLL0VftBtiAfjjN1Ju5Ll+XH3GM+J8IB2lU0xBDJKNZPWglmS2vUiywEQoYacm
h5qVlYPazgoXie6R80IYoxnYkpYCU6MrHB61xIzUyP5dRA6NMTLfZ8R7KFcXXklqdimjWEqb5l4A
D/cPkjwsvMgxvVzk58UdJRr0PQWMbfbgWvwkDxh0SrMtVRhzCcYlOAfT/QcaSoB8kkS0Lx7qX3qY
y0iIe58CIGdS7NDVU4o94naKchI759w2MSi6hKvCo8jhIqQiPCCtY1GofONql5yL5FK7/M+0mwFx
vyCturpvRFvOeJbHnFtxqonGrd0h8POiQpUCVXOtu0SV+xlqCKilpcRCWLQiXWWUGs3O+WnnOBfE
BHtQiWZw17kxmNXLtp4WKfNQLYRbADwsBVf4Ecy9xZ1E4MKg+2iZot53EVxPyrNIagTOgruHIgFE
iT2ZO8JDEgkkQHhZo5evlrKTmTvAKN6IB86w1oIEz+oI7t8Dmtv/xKmv70Umi1zCzAUwmkjbZKKT
uPlUp5ZeyWlJ8F7PhoeiynRqnxTOnCFVjmraTdWu5QjWuPROboGlMJZeI6QWXER+m55Qtn9NospT
qgt837VwoIBkL3N8aspELcLl6W4khg2z4F6zs0BczWl5StXk6QeTvWDniyKtCe6TLwAUitlrwie4
hzHIARFQbTpTlkZxfIejKuy086w8bWjDQwQbQ8H7nCiDRiyyIMQYQybmXZogDL3G75d8/0HDjlQ9
2r3CkgSLKngfD2R5x2Qiq0v1/I3F4xVgcaTPFGU+Hyx0qMYOYq+cplvvv9Ave5z3funPTG75JiaK
p9GAEORv13BtpcATyLVQztEDd4ENwLdTreFBkrIkmBMG68ZXu14xRG1z4FASKXQ7oe5kKfKimQ7P
5N+u4mtRNU6da1fXI1oTne6V4KvC+pvOG613zuvUJGk/hZ/JIWv6H2e+aqQmyGUTRksOVvCL591p
6wUmnqNjOUluq2uAQctjg4B5gCBWodju/oLlPH0/1TBHg1d0Z1tgzP0e1Lx3QuXZsY3K5Zke36Tf
i1V7cK4bibbI955TTrMAnwij/SdIrWaydFJO6M2QXSVFjY8jRRUJG+6vFbkXfwWwR9nzzYxzjGV4
qAdNHcyKJTZgNXz8Z3Mf8/C2R1AHr6hhlfKnkHQCFW8/lim7/zvTiPjZGgEpl1u9qKN1a1jKZOyu
IDYBkKv96X5DDfbKh+1jELSUekhscAlUxfSt+nDRxtZCR/F2gQYXCndyRPkUrWuEXOPYEHjbAgeI
nFIL6emjMUIH0UgMmjM09+l1d/sG2OU1lktRfPJAGG6cbmAFUHMwPi8EILaxXpGUu2jkTl/SltHl
ppiKtKNs+KstX9Oyh4JU6jABPQCWS/fLnCMj46ni8IShNFC8AvO0pX3lKrknI1Vn+fG/G0NBPdJM
9kZ2OE3yUH4D7Am38WPBCnUiEhNySXTyyzesuubJrEJ9WEtSb5bQwKSAUaMeYOLES6NvRJC5yZPv
H83MC8eP17VLDtfjQReW8bLb/mcKXqowYnhLMUoEUuGKcCCyTcZ0ZeDy5gmOkF4saFTpHymAIWcv
wHeJpQcoN1+tI9vKQRAHppkUnIYsRtsqFoaytPJpEyQaNdSUvjVJnYOr50G4LGnRby8IRFZTeibE
MgBKHIMC/V+wQ8vUH3sXvMPBuvnjtAXa+oCanlC61oSeioWVA7LsJzRBzrOSn8qp2DdkPOyVZSzV
ZuFDqdKesSNw/3zIQSo6oN5c2Bc5SlGkthuhGs+YXXJ5D5PY8wk/7opzyclOZyLijJkjjjCmuBJN
q3dIcVuxNiB1LAhy+O2Q6ONgC4bjQNvGoJWUvpU9V3fUaukHaxBTamk8JC4sULfLwl23CaVR1Yq2
zlO5/Y0KOYLhwjm1BaHtBUVVjU3uhaHIxPUdJdc72ZpmPYwnb0ohH+Lf0mORWIjBwWX5nPpLsy0v
IiPx6XGB39o8nSKwSc9iEX6CX8F9ykUg+dv2oUKiCnpV/1sxosO+isnkeFL7GoWwV8Jt/viWQiQV
VdRPhhkPulxeiEIgXkE7ocOxj4MbRB+xIKvop4NvCF9WnsjewUrw/LigqEwGgQIne/l5vzYIwj2d
9M4U5ZISKm3CYdxrLsLbtMsz1c9F7tVZvci5uNN25oyvnaxa7YzBgjjFRz+1KS84jt5HjnJNKoCg
CqG0VIelujGoUQJoiaAtyCjZ7wvfv6oadhQupMFVAUVYwgtLrLeon76PJCYTdIfqigi/ThI7XXsf
u0SStJhKZwjCN2gvKVCHTlqzMQuzxls4rM7saKDmFBa7g8TYKdBOpNP+ZC/76Npjp/DsX1JosnE1
NJZkW83WJeOyIqom+u2q6KDQzP1kwHPog/2+8wcI+aPc0NwrynjRJZMvgn0i0p4rgQJKQp4itVWY
PZ/t/T9rwYuleVVpNkthCToVfPCnDEgawWc8isWyUPf0HF20GJbQGOGiIQ40FDMBRNwzEb23t3Qx
hoXEalOfeNGZxfFp6dgZyOHcS+ksJ/1120vLfxKOp0USl9YtZIHABWTbcUUVyQOJi++9yFvD1lAJ
1aeUZ0+eKp87kQHfSsLTAsLprRH0rwkRcjkN6noqrR/35rTMYqPRsia68IEJkCTxQby/9csI4lFk
XORJc2cMsttJaiLDLveofYBMDbCmQq/aYEzU6yoIkgOPKpAUqxbuGOantvzxRMSi1tZF4Y9Kg03W
jQ2VYNWj2RT/I4zY8W2dfK35ao/Qg4tKWUgfYUZd9xx52y6PLSptWyoOHSJn6MxAieh/xwO1h6ra
EpQrvSaJoBm8dvtSCKbpDmU8jH82o0rLfW3NZQR9QsfFtK/Gfws7Q+G1RHWOMtMRd/0zn/Jp25Ak
gcFycRN73fQTNMjlF5X/jTyoZSj6YtkT0gm2a9CFBar0xeC7Xngtp25uv6E5Pg2Sw2HRkeAloxha
x7o4pYVjRjc/WnTsH0zHRlLuq8vXd4FdoSSQym+yMLsS3F9JqsW1EdD9CMk9+f9hTUlHhoHByHOg
8wnhnHPOHxEGxR5gxQ9gSS1W6bFznGK2hx7LJ+HZoKjWIUNiHxm2sxzI65iRzn9Q8YfwjOYG7LZM
v/8Gqq/vFaTPuh9diDdSFre935g2vOSz0p1YS0ztaOZFyXmklNcGiTNZ5rDgzaN8AEZ1bKMGCEx5
oIvTXKNnZvBaAwZIEOpUA48ghE6eEgMU67YS3soLxetu1XLiAjHj1DIkJ8d7u/ETPc7KIDPveNSd
ZE/EQjoadQRG5h5Qr7XsNyIRSvLexc8zpytXPbFwsOylX5srGxq0naVNN41MuuIqrXl4GA8BPqVX
OOmWMH5FKb6wvDocnf+07NH5C2PwoYY6w0BTNgXAxIyQbxX5R2G6NMt8BkveyJxX3I9zA2vV0DEm
tEylRkQn53+cUmadPQlMXvbrH0QA6r7tlYGWqmy4odXOZ3VwhsohmxWtBGZd/gQ0B/B3YECc1OrI
9ylO3XiIn32yMGmDsh+g7uweVitXjou2x0qKmme4XT9jn82G1AKUmwgYR9TNsFP8t1vOGlG3aYvx
M9IH0KkD//QVN1VWKTxzJ+8ph/QAIpB5JOLW6MtoMPZfBQlJF5cIReo6vucPRFl3QmLJpyhYFlJ6
kcuLdlGnOIK1dI/zmbZ7CEG5wrPr64ohqxHo6od/q43lHfLq/1x8AqnAZQ/K9xfJMTPJoS+1ihp0
UjUejoXxy3Znb1omfuplvlZ3qBEMCIRCnUiVg708tz35xsg8pb1p00nWEnT8GfoR30DY5dZ6zKpH
LaAVShPmplkxUxeMY8646JBiFHEPIjjua1TlvQjc1lC8MmndYT+4ld9o/PUhllFL8PddB2UY4+iD
DhzBAwlvwiatJ97MpJ5h7U0Vqf9A1YI7giTVi8RLGVGsDzKl9f1f18k9fMwBX5OGSLO6d64/K3RP
thXve0+IIgj83vcJ2lz4OSL2UbrvxV4au3GwxkLYiFHIKJsSkHuZS8LrX43adiyc2Jknw0hfjA9f
Xanypq1YWBGDqIi7ugY1kwKcRu1HiY3MGGdhVas19bEoER7WpKznKL6mmj97jCw4g5zVIrbe75cD
c1tTPJh6DijSztsNZwY1vNA+8DHT/HE3a0YLLz74A3SeVZ/jqyv02xgTgIJTHIEcNZg6xzBMF/qE
12N3CL3m01ARHu6h2Rc+wKtSSi7fhchuYEIEkZFP4pRQM52axmEAf+CU1xBagDbKsvGOdHdgPfDu
Dw8KIAgr33xZxGr3wkOqvpYSsaOOKLC3i6DQFswjsRCETZ0mir59fHEmd8DSPEdXZ56/FIwVvylG
J2zufIT2q6NfF251mdjz49NebHGprdQdxkmTHuC/Pibdd9VpYYLVL9hjtnXrRqtQP4ekPHX7BhN7
+3U27D3Y+LmeenkILLF8/VtiXX61LCD7P7pFaTAuPb9/pPf3hpT3kEkpuC1isqWYHdL3U5fHjL7P
3RnMKpPanMPi03PokDK9ynj3JqKAiOcIpaA0dgCWN6IaUZbjYvc9817iag+xR9/7MFpOd1xEec1p
tJHnVRg35iOQwhoHL430Jt3g7z63wKbOnMDOpiBJ0LsIlR+4K/zSuK/DeHzS67k42UHBobfIRiCj
BOS9/sSpRlQmgQ1xhh9k1LPEjR8mM0ss5Ldg7+mjVmF529FiFJSRnSkIsh7g2wCITOMlbe0d7KPa
f1DLpE7hwt5FFFglLRuqrdJwPU1n71GuNWDs6D/GiGPZkKLq8QlnjFL/NINGQFfCpefBIiDKbFBK
RvzLyth4j3+uOAi2dAYVLd4WszBASzBB7LAYWXf/F7pEFt7CWTg4rq0NAcHke+2IQKRdYzvU1Vez
Nb95XtobQ97vZVD4Zc8LmP+gC0rZWYH/rGcMOjeaHh6AC6MXaCfik7UPpsgN0yM9bgkH318QGIsL
adw/vub8jV8rfVicUjWhK6VcL1dDZ5YKeoO/vLJIj7nytrb0cNNShvim08NX5YbdCEMvWfugE7vf
dPcgxnff/Dt3hkDXDZ/YLZiwkclhJ+PD77ROsi1GEopvhIJ3bkIdqC3jUEgPqpGgxm9xIctsQRo0
61xKFlzH3QDfJHUYhMF5/cf2ClxPUb0UyjBSHzXJaaUKhfFBRxXLuy/d6DtOg/veuCldLjF8Sl5o
hhfZddmYvkYRbKr56J9qPZbUa8l3rBIIlgZRsERaJ+/MLzDF2i7wHiRZYzIwPSuJOfQMC7MQ14Nt
S9UH3HZYpOTXPIeghjpT4lsKreYQwavT9s90wTt7FAzAruhQh2Us1Sgi9+j7sbOUUSajefX7Jr+8
Tcb4CMUX7i2aZ1zzSnTmRIDQKDzVH8/AcmYDVWYX+dBBxXvcF01dwpTxHU0MW/6wHsBJsDY1GjcW
k1ALPERXMmnpewFyMFdVfh1nP18yG0jBKWwVDvlBy5zbeK1FItTMrGBTJSwu7A99G86H0lKiPtrC
mhyR8nSOoxV1GBIz08Zdgy18l/V+/9KO1oMK/P9biEJO1s3QA1pHWbo6wprbnzje2OtmXHkNmqmR
LIl5OQSYj1p1aiQ1ISMVXaAtTjKbeeQpb056dM5wZuUgQp/nZdbdR3DcX1xiVdHuqVrh/gQLxChg
5cyc0a/aTe6iwUVAArzCMNfaV36LTP762K1fotJ3/ypGl4MVBTSDBv5P4lJ5BwXh1Q3wXxBXLIcW
AEr+KgMXruGZx+Fnd/P1tJ7VekE6eCTuWsLDV3L0LLnGqHHbZu0skYqbERUhTP8w+WMS1QqbfKSJ
2CyTx/vAM5PpYs5vz9Ux4Y2YNqitTHoiRwMb79/xOptHAl8Ntz6dICNiIo97cHJILTutudMcpw3w
G37x01SRthNbFLl7kdWM11cASGyLJWbLzWDOKD+Z7OZA9DA0a+OhKkDxtDfBgHxwQ3t5As2aSv7I
biTsaaGva8xPVCHeklPI9CvdZDQA8T0kVlA+BSBqDN0rQDQV5NwNwdqR5+6HXKN9ev69TxyZX8Mh
64Zb+zNs45sZlDly2g9MiMnRBbnVRNw7fWZV868X0x4uZRFmxvN45b+GDfX35HOlG/3sAxlkj7gp
Ok7Yd4+YNa/cCt9uk98yGABhRufAUe5NvgT3fsTu86YBUwC2TcIx9pDGf3nxYd60NE4C5D4pLvWO
uWSiTAcvcjXdNKKD85ReFLMUX2QUINCDwp9u7ljcJ6Gd6Z25uNJgIrzG2U/aKls3aX5Lx3qcH/zj
4p2UY5tUpTz65r1cVfngvRL6x78oCrYbUYD6mkgtr3XuFbgJmRhck2X7VJ/sXnfW0UtV40daCn28
GgupGFwoadlT5zopFcsxpq+SAQPnL3icf/ornyk27ZWLXbx0ZFbEas1v6h6KJ462IDqzUyJl4w/9
8CSEmPns8SdNW9Mw4KkMmSV2+xjRJ9vtVc0KUM1x9XAmRsUW3MPVHohdAJE+a8ZH8wtKeQAGZo+T
hp8QMyw4xBVYy5AkbJ4D4O94rYqzKLVtvP2kgXQKPFF+nPytY6X9zI5LkVJKzz8punNswxTyVEgb
oEJy51cdLY7NyoNUQBTw40OPHVRo71kPdQLugqNfMzrMO+yUcY1qFwqI2WWCHwLqg8xQmoGOkdFt
t6y1AxM6F1OcJpON9XTcwKng12v2MvYElBkgupuHlTEeoeoCqzA6vy0yciIPGMP0NA2w+8V08p3r
+HZtgOmRBDcM43Dclo3n28ffqgA0L3WOXOcSaQeIXw5rWGitTfZ5iApvcY6ionUT9bFCxxPHgz3O
uAgA8JMYuRErbx9M6lVOTDLJujewld9TVkdAH+ygOmv3CLvqMYuNPZozIu01I+DB5ey/8I4SDB/W
rNktr4dp+tE2jyFrCahU5dYMrNTWQ3FmlOXu7/YEuWqv94KNEU58rCmpAyABqheUL4WE4xC7XesA
BTr/uvyUMGkhJh7AAuFN/OFqw8+aaGCBCVJwps0dkP9yOrlVf912ePTO7546mCN4EGyDBwg3PmHX
QwotNTXk1uUjO7A0r3Fb26DpxeQ847fo+eAOoyrnpDNdG1M/dIHet98TqhQHvDcQ8LYwCKe/HNLX
DkqD4xGC7QFhjYfUoaWVsUrfhY3AGkHTtHSxhlf075q3cxd0Q0RbzWoDlQNuobq3HERQFq+ns7RF
OoKx95tEbZfb9m5zwZK4+rfP8oVqT2ct8Rq2WZYoUj7mrVKn3OAx59YPAcOtq7IABew/+pBwS1dx
Gc11Ko2sQpjy9jO3DNp01GhcRamL7dVm7rbAERAu51VlW1RZcp4m9yq0X0Cvoyo/WifPZluiQe2K
tPyfDqk34vZXJiaF4u3ZNgIJnY6lLVkzpilpRelll8cOFE82RER8z9iwK3v7GjnYPyO7hy+2Mcnf
YMms5TDgdbi9/0pUikliRNhEYZQ3O/XiRAoXU+jiQgZvLVl9OtxZbSqhGYu62AqJWMr65lCq4sXz
j87HPV1BVADWIvjk3NxRyK4+ydP0iuWSchtAVYYJjhadZwVdKb3tC8+Bdnf+TMM4vdEBn9punP9z
CyjwZXI7GX0h6xKl517yWyUO/ynAXVN9ziproNEGScEzzONrInEUBzVAfwCKep5eafpUeh4pryfi
+ZIDA1cKQEG2JF9BTzEbFIXfXQxhlnhCEatrFf+lwG8qqzsx09P8TbTqqtuXiD2/uUj7Ahas/K4x
9LoT7rDDu3+1H+pwhoKUTTVfmxYhy+w+tV4MW3/q5tZIw+0JKlZUKuLxtJo+TVf9uNm58y6Dza4Q
t5qZ31o6JAGKyjtU6T4BPXNr4nxf9MSjiBg7JhGmFWzip8sQa4tcqd0UPUtMGFac/o2ejY66xFVG
J5QJI+8E5wPGPUGiXzJkLQB1AFgDdJhsUSw0M2ZsKOh4y3ptUdnpQb0DCZ03J4ub70pwTcdaqA/4
ECIBT8EB7Lgnk8aCi6PM3JE0lmMt01UWscLvUjMI8Xe0TJnWXkQEB1cjm0DLjipYrIoaRTjzeFKW
+IJ/RsUxc1RoKdoKxrjXjDHjzznLaR9ADzuW9qjM08wBAKwV3G+W/4A2n4D58fq2WtF+t/CHKFRh
Ne+MUgVZS/9p6tEH8sFw7/CHFx6I9zEuXkzpe6CELBPXEcxPz0aiKCCBmvjrXeVxhAWpwm8YIFuc
f/anclG9iRVoOtO1TYp1XnKylzzBIO3yMxp8bKuqhcV3MQpdj+paH+vmi2IZay4sA4L55+5H71VD
d/xpXbT3UiGpKUp82bHgZgzc7U/tZqhI4TqEpeALqnaFBw+H+Lb4wpbA5N4nTp2rCJkawYLqFpiz
uLrcrIM/f7gdSNG+cpvzLcmsZOCaBFNKIj5j4D+5PFl+iHru+tMVidpoIEARrV02cWZBkRAJ8h5T
eQ7tx8xZ3sA39V+FMYRXUhSFePFSsa+D0eNKAppbbQfTjpopQKFc0dws5C3jDX1xKQIadGBQ1lKr
9Wh70clAZhs1s3UMy9BOmBHOrs6POB5sed/yhcWdl8Fs9ATUZW3lAgpM3yWkOLnjCl3NG6WrookB
eUldDzQroY3yDhfddsXb+iSGe/Jc4vkvd9t9nvd4el29bvDcLDINLWQu8F1CN9V7dZxjTpY7U8IQ
eRmbzdYLvaxfAai5DyXOC25oScjBOGAoPJrR+XqMJBz3V4AuJQw8+tyEMHhVjCy10D1/C0Um5jCz
/Vdpijbh8ixtdIncd5CeXyzMBdtbvH+CDs2wReIYMtiMS5jqdyiE69PRgVFTPRgw6cx7C38usdyl
jcm4Wq6CXSnu+kzCnXNnqMrpPImnnRteXBiDlULReTcTw6TyEdT09YweM+VEYnSlc2/uRgl6oWDF
jTk8AFgA/amadxUP6K52wvbFD7lLkD2MazzgeWnWRNlOu8uNM+08PJSVMejMjsm10UJivSssGok9
ftbYmLmK9l3KCY8YeLPQJm3tnTFl2Kz5oltE8i8G2zdBxjJiISBP60cztP4tTTPcQfVORK1ScTN9
tm97/oSpEO4Z5IYAAf4I3CpZDHS7wx/bOT9nQr8uNIKIB8c4i0vXCoClnSai7bfl1wY1CqHwkwDf
7imByh2tKX/lGAK5Fh89Di/Bxj1hcFtbf6MfCs1o2SwqiHDxBkJcf3Y2YaQnpPTdNG7VNwFcPapw
uAxJ/+AXwCUdmf5P5b1+DosRI74Krl05mUhziAde99GhwMCiI0ftV4YQcKWUhedsyv4wK/c1pnQj
vZaZkExsS1jF1vpmTs2LmxK3Cqv4q74zETierWYvSm3ozDGJoY6Up4y79dhAu4YTwfJsE/om4MbZ
raBOs2Qi8vBIFWkC0mZJB/KS96b8o98UVw9IPiwKyoMTCEsrAme2RKnNdOdbfzpN4JcZUwejQmPR
KeM6z1Ymt+B6Hbxo49LuS275woS7Lwc6JEYTBFHIRtYMxasmJ5vaYBe2BWsKBnIryV5CwcnZECSS
395F8VqK3eSfcFhd7UM0FE/dkV7HJKHbUQgDPWUQJZv854Ou/pQR6PHVfUj1AQTiuLPk1Qh+hTkN
UL5+Ytdf45kswjKr3oHzqRUdmkHfgYUD1jSyiAGmQZqw9ATDO3dJHcekFUERXP38CTa7hsssxYah
e31+/OAqQJ4xBt+BtycmGdAmqXjWtWkvlme5wi2R6WYiFuuDbJlOHfDwpvhrgfGP0YA6zsHglA/+
nL9+0HswtASItv95cXWhkzx2Kr/9Rk8OTvk19FmgqOxqKeky3TH2BMLDXKrBSUBz78i80LQ1Ioo7
DWVoJrn3wKm6B7CSETu6ht3bVkqzJw5rKo23xjmrZgj4BcbgdUVHXeWBB+2q/b0QZTggW/BfbVqw
8d5W7S374WsrS3mHyMjNiphMrmZQt51MRWjZcOAJUiH6pG2Hdyecs1PrQtDaMm39Dg0ryqaGxq2t
j8Aqhni5bp8yWLlZyyjkU0UgUg1arOL+PZLnZymQnc6bl2xmN4Pabcl5evyd3d6IWGT416dJwXmK
WtzHX+787kYtbnGR2Ekk7hxn2QkvcZnEvD6f9YTUwjBWfPNHkGFo+qfO2q6fTDF+GR4DypqU2Uod
TFNvSKLf5GMl+cNA2AnxH4cDHZzUYi3aIHBUVBbKxio8nY5npJZTNEGGz/fnd98iGyDTsKbGL6xy
I1ITjW5o3gqe6DQvb/9oEQ3zx3fHIrwgawywmByuRhPS79syM318tqaDExkIGGMBl2vN3W9ZpgCe
9Bwu2jqyMB5G4N/TR7CoKXnwvzbI7gIPxIKoQ3dTssmaDjQ8jCCpbavwVm6dFdHrK9OdfOeQo6lN
+l4Q7kxz0P7VK/b0GdxhNhFwP1eN7WHPzhHzS/16mbnr8yzJSmUdLSEQ+ik3HGG920wd8QiQJTR9
GfT/0mENZglbyr+eLHpoaeZYYZPFMDplVVztuLg1XzxXowqbhVSRXoh/2QYjgybhiVtrlXWXgKpW
sQFGiWJVi3i7I4xGygZTwdRwfvwpr8L2OFKekQ3JpE0GgPSFsDt32OJnGAmMdO8I7hNOMiOUvA0p
3iVYXjX6K2x1U/IAHDb2/3Z7yO7BzJQ91rn7n92KDOZ/2RI+VfWiu94OwS7fygM1e2O/mf1fXNSq
g4BUO8ZE9L4lAoUHM/+RgnRm0XKYybqTkMA4VkNsEBPXcfJMgaj0bf7q+uKT/TZo/+XhGQi03Ud2
GhnBWKCRIr7gb80+ApkGmwzzUWkdcy/8wPG2Ccjs1+3ZmiY1H6oe+4KFKT2z8S6SXyz+mUsXnfQ6
L3ZXRON1Co1L37GqzwTWGHjGNLeeMF2ZYYDzyB1exHQFvS25gDZi07d3ExIexmhan+1OTsYyy6jZ
qrTztAFvODEeOfeh4kV4yfLk6Z3kuSlqjDEZ/Amnj5UYolQykpR+1ow8lJdNbzo/8JQWndsRRw2Z
ltDnwlaikHH5tOCRsT3yTYtgeJeTH0gJsztT9MQt8q16mskiimzOEKZZeTmyiYCuxhFsMZ/tv+Hn
UUjHrRySk8jGrpofQdCH38brQ8XIG6vvBOaEU/7S+n7iWgckWVTyEsxIp95kDR5TieGhaNOfMhad
Uork9UeaD5wlGB55duB2BjKxEivF3tUfbgbC8LkcOWtgTTk009H9t31BeP+czZFOSRPM67NYDjVY
0uSCBXVCSTHgLqLwvfCqFW5RlpiC2EO3WnPzOWnmv4s+M0oVxbrIrdv5VaQbnQm2oUOMx0vdezxc
GORYv1TEDkvnrobWUuZcEldEgss/QDqvNo2Ke3cGsXVU9mMI3SI+/8YfpxrpD7MUTgsOYiJJdGVz
bQMwKYAu25jadBu4Yg1ItR5i14RUV2NtyYmymfRLko6LQY1gac2QmZFf8L0xL/ReQy2xpylwVhuV
f6OZ1QgHNXKzEdJcI1GgK2xFf0rDCC17q/Gji9yuaftsgDUwhtzMPFj0ppFRfzuewDdjepuFgOP4
wn+5pSa4RemswR9cCcB5ST4HIqMp1BENM8XxyV3nd3VwbMS9oPD/NfHlUF9t8pZcXysoImkphn7G
b4/fsIojVfJNIAaAGLDOEcgjrGXgjApTGjZMC3E5mTpwO+TgxUX+IP6eKQDQh0IM3moj0CqPDbur
j5nqyX9aumbuFuWEpoJ3Ii+JYvFXTgDDwFw6fWnAjWbYVTP+cnUfxE/IMHpKwSNRf6eH+9zaBCjO
1JWDu+GaRE3+EsxvFN3UtOspHlYKeUUFnyvDozhPNnY3HeIIdZsHnlyXypfaG8KSwHtb81muAO7k
fqJsx7vG0LOyAkussfSbOQfFAoXPKdafk2MNi1jNAIGpbhdKb5mkK97m6SGuOce8myzS93WtGz7Q
Sr46mHTOoexmYb9hp5QQ80YVMyDdwn8S95xEoSS8YrJkOsu16P7H/bcA7EuW3IKd3ib5iVcThebd
VA790pPF2FkLVCNj4+RfO2A7n/qASBvYX4m3fUvuQqSxLZHe2Xk7UYtXtSsrTSIpXdE8tsfBZZRh
XBwC3+cA/0C4W0Z1T3YBDQAsidQPeOKai5o5Wbt8TNGSrysTwATtsNBJHuBcgO+74EsLsAVX+9Yq
nG6aZingYDL92bkQ/rSsjCKcyqOJCy+Sm6xUFN20MAObZ/BYRv85VHkYzFu209Munu3zTD7Mgzho
Xe2edyj/yXzDQt/DNNlf8fQicIV/nabmPt/jjk6L5gwr0S0BBJ3/GcRGzEjBXMKFW8yJdxbTCDtL
mov6UCtqR1HVZdn1JH1zyg6WWMmijahEggEYo5fOsxzb8HHL2OqVtKTVn3nV+UoG188ch8TnukFk
wlDLHUglu1mNPvoZV6n+IwsJAmN4Z/32lQjfamDVH+Ge8zG2uaoD2aPyz+ZDuxES8LGpVroKcdYF
lNzDJ9FleI0au8QvDu9zZU73QSNI722hs8wOIKAWugvclFslA4l/fM00uVeNI1OtErNgYSWRbo0l
wFEonfiPvwYuOYvH+ignJhXDE0FyfJfTjBnQMPCO/BdYKXJlvfd3KfWhtVl8zvf4mUsTlo/IdhMC
pn5jBQx2+EP/vSENDJ3VghGAvemKSZhS0zkcBGf6cg2S2ecrSCz7jAArxTW2nVuriYxh9wxQ8yaL
J/Px78R3pfkzfDoBnb5J6Y8Kywncnbv86bpz1tBEqRAR8SL+YKT3F/cJHbg8bEODzXdJCiGZ+wwk
qSg33TZypNirMtZDPifA6Uk13MPzMBwRBlNbYoBKT6lKce/CxWtki8WZ0MgppySZV/C2JHn6/YBf
OJGQwUuAcbIB4xZNYMz3pwvX4vQeRd9Fkf6SkRDrvxfsQA10KrB9gljgSda0Id2Ts2neXidEArDZ
IqosrEU+iVAF/oVY5ztEhi/MnZT/pn+yDYfH+Lm79zGxXvgPeLxxExoa42Tobk9m0z7lz7A6qXgN
bndPp6pnw2wRwoPdUOez2FNYpSQwMISAhLf6H51eb1voOyKZg4nApFtIOyxAMfCHb8ZxF+mFmFFX
iwRuTjUmG5EkjHtBcL2Gl3rS35We2jWhOW+bZhRpLbsFuBD73/iJ8U8tCYYm1Wt2zAuqt2NVg/Zj
7F3bNLkqYHmSgIKs4jHznMn4HXPlE7lXOUxZTeq7munWqFT1cJ44gDFmQCLEaLrTP1Q5oFJmR7H7
zoGpPXqaI2HP4KzXVDiLucDMcBcFpns7Tifibhv8LzI+X+162wSbt5LWylz5EAnuoWEr2WTrrwP2
1+4xN+Yr53NZLg8EgG0oola8EgWvRTV7X4pduWM9SnFgUOEC63Z7//PxP6evJfOIv8nNU01CpJ5M
w7uQoimDU4S2QdrvaxqCn/D9pGlTq+m/vdYvrNcSvN3Xq5P4MEXwd9Pm3LJUv6lZKN6w0yArycEa
q5MhcjR2f8NotfqmUKj8GRSjw6Qk4GGaFxc5k10U3QWYbJKIa4QKWhic/NPAGydf23SV62FdKoW5
10iLHm3GQ7Dn0bHWwl1z0g/RERkU9SsO/ISwZCKLKzgJ17hWH6M87JJIMGsPZECdrgBoBPF2GLvu
e2MMmeJ0vxV9sRloa/LqlnPEVV1P6RB6jWY5zFq05svBYm4Xsmb0WSPUDbOFxFXZOv6txoxgk4v2
XWS/RwCVOD8NukWQ8gEitgP6F5NJcQBnVTkTSS5LatXabunDd5PGcNMl5E9v38SoF4RMjjEBjFyY
i2Xquz1HygUQtYD5KBplR5wNNAvNB8QANvFAk2FFmuAqOeHfNOxg3VmGiJ2XC4ZvqyXBhNphI52l
RJPsnv96Wj5SlK2P0F8Z6r4x5NMlVA5xdf0SPNcMPXaaua5kfY0DsA977hftTTkhtGZcIyptWn/1
8MAux/TyAEcOMaQHac094W83rwAl6mLkN3z2YKdADqodPTB4nOosmS9bmxteZXyzDI4MV3S7wF/d
3j5rdm076I4Tkl11LuV2cmfDHqIhTz71cN7IBr/KrK3NaZ2oo4HQalRfy+PegStWkNbCzuTuu/ER
YlceeXMCgLA3UlAMkre1osIm0viqyeAOa31+YKnjVAFfgMsp7NCwIdqEvlhH7DMW5FJVUemLg7wy
1KEjIGqOwCj5eWrqHF2f3X4nV4PGAu0GT+wzCD8nKAmPb4HE51RceDQbzU3Dxee0F8Wdo47nhVFZ
YgyGGhYvoheV/+WxqV3Ibv0WnNk1vRRUORWNyY1r4KZJTN4aea/GRZlZGaMdBFy4lcNFO0t9/g/7
o8C8p+JhYI1IXuUCn0VNkD4B+0XTPvWYwu2HvenHnMXjPMWit6fTp7FaA5bfPh9yZmKKfWUN3xTA
iny6n2XhhOfEhO1LPPpOADIq9tgD5bcpRAYwmYbVIpD5pQIjLssKpkT2IjgkXFkP1XRRnAbJL48L
ojsWNzco25R4volYjHjM/odbzWK6Gt8ERtzdLoqu2Wc8KIHJFM3o8D4esXe5YIKuKwcKTgxpUBS5
9xR+3gSIyfRrHV7V+VNcTe1jFleuctOq6wRZkSZY+u01mTUC5wcsmDUOcDKdatcOKmxueWdACnER
74TunsEXDHnZnj0Ar3gELHLPMSFHErNNebXF4AhdLqDLbXCR94mccwcCeBrVHCLTu7Y4Jf0WN5Ie
9oTGwiM+O6DMXjpADFEtD9uMLh/5vl53gr0kZ7Y5hWbLJp7oAPSUk2gLrgOkFsZv8yYckmfVu5s4
OtY7vWsFhmV/ozGrRQwnL+P/Gp1MF+iukT3JWsjzXg3blNX//MANFSu3Xa6GSCEnxAPh+z/RlCKs
ZCw0S8CfsDP9SUpF0FRlLPooJhLE4VnkQQcvrDYIbqIWDOZFYKIEO9EMqWJRKVqezdj+4cUbaf/F
A8HwXraiSK+HajMelqYcm8PuGi5vSd54wSLze64QA0klD5bOIxEK5WGo4q43dszP0fyCE3VP+Cu+
hsFnil2Z12LO2wRHuFue2QK3+yyqY30t3MZ1pO7KeLpTMh4dZ51O3Dnn35DHW+NjCiQm75R98Bnf
cUZOn1lzVUDmIYNiDUhY+agVIffb+j1xMFYJy7UOEdEPfRjay9DJa/ivTbPz8Q3sb9pDFG0fwk/S
ZRYwYxQKur8kieCL0g7VKtWwqttL7qjziIJDnsH+UUgV4aAMtBtyjDW3CZR+BNhfkZ5VW1aRRWk6
NpKPiojUyOD0QmOxxm9SPutTZVTfIn/lIpKdHcgCEDXvyI6LtXm1TnD7+PRtBPhGBBRWKW/Xx87o
2SizgmZwU4y3FtsBqmAqVZoYtrLfo4NbczK7lj1lc12ZOt5cRQerTys7QVh25wso7Q6aD2ADMtRI
//JzwfjN8t/yBsDbB3w3Sn2z3Sch/UmcN20lmA9eaNGu8YIqe4dwJxQ0iYxlZrsMCu1GQlD2Dtkq
bmYHDOeQPpsBRe2KZrQJD5l/Df/E6So0sbyLRqo1lYFg4i4HYRSvvfkA1LT4kP3KbK9bAppLlCgF
vw5EOVhCMvfGSnBAT64Qvv73gS4X/spyno47LG7aSkSojAaXu8lxv3xRdU+iyXuv7JYKHfhAW98L
qQ0JwPxVwRfzN0iGOhk4M5MEIOVe64DFZGj0n67LwxkEpSxrXlwTpF+kvjH4WdYxKpqU7ZcXyCsx
Ma7iy7G5miQDRoCaNfdQrRpx9AhmgQrKPt/GDLoxIgNt2vArExT+rTGtMFJQhq76OxT/UfoYSb4I
fA04mj3vEmPUOYYGCEd5qe2sAK4IiPiIQLEBYrpNA9nibUnpd1IVJRRO3LO9lChBaA3zikstmS48
CgJrjzj7pftUYFgx1iEp86bzz95JgROqfrlVlNuuiw7gv3rMq3faVBdy6cCS4v1kH8qUaLpXwGyr
CAL+nfsZhbKMX8vTlV8FPhPFS02z1noXy5KBVEuy/QvI/Rb+iTPi6WwZkgjBN8KZ9kcO9jh8qRyF
MbTw/Q48tSUWXqJ1yDEtmwn842oUhnGk8O9yfIuc83gRiHb173tFfkpQQTyJ8pmSu2X+OZXASpnK
tWv0Ewkg/zo8Z9BdPPrke4ufWbMmyQ8IJk+qHvM8XUhZrzki6KlGyy1TqrVU2Qh2accL3wVNHMlZ
kGBLltb1Db/LoyLMoiKKqD2uYlI+/Y9m4nElzWwnGqaONrlfLSVETaKGWvP+PYmLH/o/c+0TGG9l
TwdiXDh1SXh/PQ5vd0uMxtPZO61h3EIqraFwcGWJg/N2D1b3vS7Bdl4vqyRpT3SbaF3eqgB9Ngqb
hYDX0birygmuFdxRJ02VwqsNMCYCnDWeWEAxJcLyAjb0miMIzueXIigER+HABG/U7S8chn5GVnGS
NCE7AMSVqSDpeX16pK1lG5af+apR5hFnTO3y6hZNSgh1omVBiQSaIRZLqk0Alw6xFlobiEPzycco
V7K23whjNHjhjAbH7bdtFgaoP881WLvV1tEfekmTv781Sfavl8tSmbbYSt0LfrVE+Lzrr9ajCYCv
605lB+him4OPmZQgwAww6J344Wop43YoABBC54BDEi7W/aaDTAFSdFSGIOcyeNH5KVWoAAjaiWGG
NL0bpramJpjgaVEFf8ZNcIVScq6mpK5XGG102fVBNSR0vMoPznaZD8JwtC5ApIR0nr+vXHyE02G1
Jfj0r02pMDhk362wzsAb7rnJzlyLZEFvXAeW/rXr84QehPEZzVNE6sW3zx8wGRFzw2G9mL4cS42F
7aCgeeqzq47Om1aO78cdhBV99+nVf+an1YH6SMiBVzgDBxi31r60o6rMzobjbzmd4AHJhQd2RHro
BPqk7YM+i/5xu1cP9Z1NrCHWpzoMuGrqUDMS5zNnO5ezIOvckD8AF4/lI1X4/GzGJ/VAtAuag7HW
zVWiuMFjzzCwRcBe8gbJ3noArA0/1oC5cBvarGRlEdd8mS+ovmVmPO6V5sG7TGgAQNheZwcaR458
Oekm+Nhx287Bc2ub36qi9ZhaHp2zI31pqadra3wF4A/7cecda/cRQS3UPOia4CyeXySMhT2fl0j5
d1Fl83GJOrzexznUSmNAlEI+tq2kN3K88uF4MaJfYx8VNyubf6Anp0HLGXQNkKf1HUOFv/9WEDfi
So873wRbD242YkOAIhjRVq6hBLvKYFRsA5Rl5zBXoANrvKGg4tCOObnU0PGX4pj7zUy96unnoVUc
Igmx61inreoB5nGtnFNnnB06M4YGY0YSpzX78Qhkvr/zTUMEFK3oEWJNmOce2dPFxwxj8pxSimjf
gPokAHe1pSIjF/OwzdgyxKSgiZ7AfUuQbX0TQDhOppWfWwqoNS53xLpM3PvgYzh3/aqHVjMeE50d
uJXYKWr/UwZaNJsMsJhci6BR+iypvarHK5//yK1GnkIFY8SyW3BDHTXp3lTXh9kaZCa3uVunN0se
lnRMD3zCd8gE2jLFzYHSR+cMeX+1v0P+Ckh8kIKU+hfgOceRK0MAQsnplZhIOeo59bC5fgcP8/fK
teaaS0kKitboUlUbCr6EgV6Db8lrEASw7xi166vyaHMnD6Amj1O1S6X9jbiosGlvScrVnW1GPtZE
XWu7Rsr60z6s2TB3wGpAwvnpZMwHdYbKRJWzfSjJ03/QpZmQ/Ar4ROHeXD/iHK7+8iG7wfe+SOMi
QzOQHzvx6TyWbeph001+0alH5ISMz2PIkVU/GWYecJpXZtWTHnrqZvRhZ1IbjbDBuqTLsfhgoPmv
49NLZf2zy/KNcedQ54A3DCtmLup/8liJ9jn4HBYUHuaJeCxUroCcsnj3O4y1dOgDiOsaHeLgpS0v
5ioJiw5GsGhbHUpyA0Ov9tjwhZwZM1Beeu9t6x85XBfpJs0jCwV7z1ry0MMrRYGGfLZZiyohLfI0
M3SIYJbWFidsDxsdLJ2mXIs0ZjloqYKF17sDqJ70aNtobcf9/AJPl8Mr+YIQcUKhDhEgz84t3wKV
cpXZ4qqFK4rTBLJZAGRhJ3uKR+dbmYMs56TTYF+3hSub3CkbR6m39iMYw+BA+aUC2hMf+VA1WkQ8
UU5rNLPuoNj8zeKHcUk4DXJh0fjqbEV3LpIL0iMVHLJCRtLSN6xbm9FI3GpRP0En3tL/kMXhcIDk
pd9tBgMvOjC5KCs+qjcd0xmP7ZQtuVwibmEoaG/bZR8wxLeufX+SqO7vcwlLqSI6AydeSAqvSDnM
pI78lvg44mUNioJ5M2gUobSqbmZh4hQRFZrXpviuDAkVSrC77emo3BdTpSJqjoMHqqlwwe33JiJm
5TKcQMxtrcpS4bF5kyX3L2L7EWVJ+kO4xufHRe+ZoEImD9MNqJV57Lq4PVMSEJOuWsSy98gfa0vN
fruFLtYzgKmfl3ED/JMbfo728FQkTIPYO3xcvyaK8I+HWLJEa2anG36uyBxbhClf6Bc1KAy3J4Iu
wbY39dj9k+77hcaUmHHkyGquTGbQNIuY+KV3TQGFNTlPVc6gwdH6IOL65XkPcI7d8n6U6un0ef7p
sWdhSLYqjoHQld7pwZwmCCahNnGFcokw9eIThhQdM8nnueEGTG9UjcSqnz8fGhjwCo4wJnJAFgB5
TdREaXJEHCxOChy5BmF1PaQ6jdd3xL5fZuztl1Dk0NnDfUMDUyQFls6QCR+eBhueb3veZFCz6ft3
lppahJi6qAhCK3NBin3Wx0RKqthkgllv7W3d7kPGRP7AVbRyTc32i17F7YZP/ijyI7dxnqF2BsjT
9AkbFcUCQvY+HQWuXpOGKazNBWt1dIz77fENMk5WCctgVPrmBobXEvj1fwn7rFdwx/J+T2vPniSL
jfJAuCDUNPjzDj9BV2QV9hiP92MpTumsgrIxOTp6f8EiHjqzHdpffwz9SBgepTXI3kzppzJ0xWdx
mK/lo77pUPQLykfF2Hv1dF5EiUIG/IkO8JWR9ZewUaZ8PE8kT9aYu+yvbOVHFFanSkn9WZTHQwg8
T7yTiFq3lITCeP+Zsg20UmMJ230DXR3FYvSzOT/fRMRlOtdHuroIdtWUneWKnNmHGeNNxFqv/HPj
4uzI+V6GB1bimpzJmxm15wXxxc3Z+GlPqDvGDNRcgobqCDoliXFmikxXVAn+9stvO7aqNZnmdVQE
bcHm3iB0/+Zw389ZA+CT7WzROttLAm0g+O6ucwcsexQVPAtpN3rEq1BQHCmfQFusvnNbbduM3Ii2
EyOToDq+yvkJwF0kdJXoh3LWHaxKywmpe4J2c+jF9Hw3JH26yyBblDNJAFjfrBxCbNNPqpaBNtXX
SCSoSlTiMhZNHzvX9+pB10WF/X8a6jq/vL2PFVdSnIrZBoAsZgjJ31QGoSkcnp9U5wA51R4vaMS7
o3s1ADVmDNoWoS38oxFS7RfiBCPs1uupM3EQfNLqdhzj4lGIkVfJgLGqqiOlBFnNOQzz1RE5oOsI
EU0zWlzgxW1uzVMWYXHYcV1/iqbepKHCvvW3UBpmUnH82oJOALfq48H4ssIatU9vwHEINCQ+c1oO
+X8Eys69Z4h54hQG5yZeniZPNb7NXuGU3OY4N3iLkqApx4rdKWf6uB4TDpkyX1xHDBQ/Oj/P8PJy
V4ALvk5gO+i5Ev/FvDCB8OGYt+Ps4Ay+wlv4b/JUbYgeosf5MQPNtVXR02n9RgnoAcpjF0I2X1AG
5I213vYPxJIo+8WX/zwlwKRxqseRzfAUNkdUj81f3fg52isKTaer+Gw5BdQvsAxcaU7CgRahcaJ9
UoX+VgIadORPQmzcDEPuMijsaEh+MneniKeuz88+fnY61NTmHLR9yM+VuRsS8A/vAzUFAN5Vv1KE
ghBO/UltQteANW7uf/KmMwkMJIgHK9TI1TTsf7FI+OXXfQGoEi5+4FdbY5dS9FA7iGD+X1L6lm44
1kU86i0RLC1hJXYQbaUHz8PkEFl0igLEvwaz/+xNPlAFD19TH7TBbxNHFvGvU5H0DurEY0akBrUg
2f9Fe4QWB4XVhyF0Bs0gIZOHbh/cUPIFvtzDLKYNjLMElWQCdtTKrdubLahIeKKQLMGkVqChgXjk
lAXtUusoXYVZ4/nHP3TPuny4PYAexCKoaMxOAA3zPngJVJJXfR0gWqnBil5egLSbvBwIwvkNTE+X
wkt2DEDBpTqNBD67JfqBr1+z/F87NSJWvdVXfaUJNXx9XYGGw3iX/g+ytUND38wCJYEGGmPDYk3l
0jn6w2NJ14zxNHnRS4i9JkwixsVIOyPmVL3YWkEehl9M6BljhzmfW28aiy/gJ0vsEEOBE35Dny1b
jFdJ4KPaZ76+w5aw1GdcE4lFuwE7ax8Bx3Ca46Txt2Y9RUTiWGR3fyTV4PLPonmANTg83ZauCUTK
vGXyvVFZ4Ik6jVaCsiXb/VEKQXwKoYSI3g67O4u8i33xF9yb5Imi7gCipC1IOkYEE/undAaGIiai
Zk6mQBKOEBWbGPbOF52G/NWSMb6vY7LWOqAlBug0XJXcD/RAYKX1Ox7NDmAGOMeFZH2zsMnssTuF
E5f44UtVx26NPtpjURyimAJXcMoIacSXdjW0IwRvYWC+ynS6LlzSQtl2KX0GtFfCHaaq06ZkpL9V
XAM/ZmwHe0BSBX6CMLzsGGFAdyw1aPlqK2Wtbac7N6GzrDrtwvlh562WOYlvQylCLyvE7voW+3CB
jMYOPDD4tBNLPNDeJToIbWO6czX0twTGfXLD05ViJT/gueDK5v6d6hTm+BgbwZaMrk8ToADyJ30s
T1HkGNhF7S4zMFaY+2BkObg3W/eQarzLFu5yfGu5y1VJSilzNHOkahhtDxNoSi3jyIV5TviKqpb1
xwqbw+7MzOejmFYPBOcKgMxCjCC/a2d8txs6xbqRTKwT8HPaNf5LJuFX6Z8KmDOweCDOle+WmNwo
Hmv3paAzNoeU5DK31syugwdrLJD+HCZntvqcuf9S4DOU2AQ11jCaHfy20kBm9kkW365F13rn1FfK
yjB1rkYkS/5BaTazKoiMKuJ71OV3gysXy7ECLqy/RLKWGQ9HntCrqxvLu8hSizradTt9MAvgKahs
/ejPZgcVv5efBODvuxmhfJSLObAAxA9JfeyHeuTIFbbdLH+VlzKJh7qaBW5NhpnGF6meQPW7HzM/
b/MkWc4ExOmCMJQMa63BRIdt25iEyyEfifD4tGV2rm/U1EHVNHSD+j0e18xRkrHWgKWJYpoFoUaQ
MCR1Am7t8kc/E8gRD2y0F8cnvs2wlWern0s+k+gb0EyzSC+5GpAFiMy2yRLytZ1w5JhkdYVuIaLx
BiA8dpNzAkPBr+1s+67gcQKEuJ9wV4hU7bjkmpFVy4GWfux/IDx5JC5n1/5/mAhTIcq+wpxNxVOR
z8M3hNqwZmwoXphgA5+tgfpaLPBIOPbi4fjDnuwnbM//KUMzg4ibEqutyXePTr9Y+b0SsRBf37eb
1GiXqQTxP7c4BSNtKv+1QFjOBW0pX0Y6VHdUtYeFFlRXSj71eMy6oTIsWLAVFrj5UX4V9LzBCT1r
g83NdmcDiSaayFqmvVEY2/1K+JI+LZkCjf0VmHpeFywb45LX4rx1MuQJ6/BJIP4pMEX4DfMYm/md
TCuhxj71AS9gYzsB6F+CuIAgxlNXrtPFbyKiUioj4czmQvXoRb9kCN9M7Pfw+sKB4bzqyw38RJ3k
0ks6V7ohyMtiNmGTRmMGis72GByQ0XZfSoOYiK+R0dSfFWo0fXtAxs4Jkl/U4mQYD6q7794kvf+2
rDGDhTVNlJfn0qTC6CfB8wxgIeTr50bZfeOF/UeHMf284hEhJsSQfq2+PvhcdVcytnD5eIkETGt3
WxMaLufB44T+KAcN3OYXxZUzdXfQOGHDEiET2c5FXAYkxhjpayCkfUpBAAQc+1GnDBOF19WczWLs
zK1pxuNdAMn5nKpyiDGFZgI59wAmFbCtDkZ+wykqUHP4irTqi9lxVQKLZaAL4cWX0a2FEhEkSjds
SZNaVROSl6oHmpzigwDb1t8ad8VFOOs4cukK6XvrLDIVv3g2CTEEj+2ZI7NrhRayTY8kb0KiIWBN
XYexQXYJH2G9r4CD55aTpvdINK5Xrt7n/4pGsAvmue4b2RzqGAx4eC/hEp/kA7TQw3FKZQ1RhoSv
WCGYMVKxAo5RgtgNqANiEpOrKUiJAMw3zc6h3lNPcTAR56HhzTsD/mw3EaOT94PJScYXph84T3a+
Og+WCqqb4FcT0cul2WxFc+jD70fTAKtClN7AkO8fa5Ix+gY210Cm+LGCGMo7Bzo48mPYgw+4rYmq
O+Y5vyjBZh7s2ureOOx6pQMQW7y8qzCBTFE4f2D3mNJRpi9wTtHYolL8FBJPPFNg+4rwx1dhz4bs
ae82CNxVL+Qh1sNjS0Qra+e1kbyRGO1m4SsNTrRCA5e7VecfzyxomvIxEClXRRUWNC7Ig0D1tc+4
9BRtmWeKhaUSP3l8qTTpCWnfu5jBgUehs4fJ8u3SHfClYMGFzNXvewbzxTmtGPftBDAE0w7hCUlU
2IMKlwsRvcxULkmdsoOp5ObU+32C3NcRc5e55s7KKPLpL2QqXUqRARWqFeSuoKTRwjH9zvyhFueY
shpFGBPAM5J/dMDlUL3++6EYPt4RBP+PAeqPQALmNqO/luJLpfpwxrAj1pKjg5KgehHsVi6RMiOE
A2XuKsEdVSSwBu82j6LSd+g8u8ECUAjxP9g8u7tJL7N5CHeCTw3dwBowG580c608dRQCTJZx9LTu
Wh6DVsiie6Ftetd1YfuHvihsa5fbydcPnFS6NXfOzoJi8p6NkJ+KA36g4zKLGbxPJLGdxeoHxW5w
fHCeFld2vc1cgLLdxyQfEHbDpNDPyeuwdAxKEKyk16/jDcMqiorNRf4POLnyRUcbA0lIg3RrXxH8
VYCRbwB2Q+pyhkgY/r651QPyhvIGwvXyfuIRoMf0M+9fGMUKLDwhjVMNcJbO7hTWv1hfYbq+gwK0
+2i8B9CYvV4mdi4Zrj760DKaeBiR34vrSwIf8V0X9nTnxKkCl4nCeut2EhX/lS2/NBTECLqS1TP7
4c80FQddYi4iE0Hx2VZ1SKu1Za52PEGBzqjwfpuAjc723fn3SHKPLUWa/9vFFitYWX1pa4LyFGnH
eyJdSbVmaJnj2fMa/rbK+qdQym6tl6HpdHaNAQMosvPjvQDU4IiWP/Nhj39joQ8LmhF5vZsqcUzb
RT3AloxYLQ941/pVNUHt4FVLqELYWnsumFaKnuzc+vH0gUQF63p71t84YRrqhs+a9h/m4jpWyu3X
1cok51yDBpSFimMKmEXKTP9lunmtWrE89EW81dJq8esu933/RT9Npi12edBOfFvZeqQ1Sd5bsNgF
OqOd41tLkmqlqlf5PyMHKSuMp5E5O/n62ocUVzscl6uIklFPdgiiMEG9uyZ2bHPpj2ObLEF6d4Qf
7DliBxg35FSEpdsMNPsV3v9mOKWoRnWqMYyYlHEdILjGBG9vVOxuwX9RiWMiTqZKc/rZBeZcYsL3
j1wfPtiP7VJ/dFG1a/iw+Xn/0DVCEZ0r7irwztP2Dn1pGBON6cjxFgO5jWUI9mJ6P2ckFDjCCpJO
89rT0aquI1pyF6LR/I5ldkWhd2/dSjeN7g39DG1Zr+19AsICfEdosTpdqGv6ebK/DqFYhZHKw7kA
Q3kyLRLr3OMjjF5Ewrx19TnhLtcdJ97YxICAmY6mXX1vGIYCRLafpXtSoFcqqGHnzah6miRUMUfa
xG7GetWuCi9FZsoX77XosC/PB7Zj62RjkGLT9JJKrkeOJgFr3XG9v+Ug/GQ0VwJCaFyzYFxlgw7n
JpKATIT5tJ5C4+pGI9TNpUFlbiphMFQGqK6cCsSfgBIOAmX+LU7NzRuckVF1t79snrj1Zc3/2uS5
RAr83yjxfCmysb3MyR8ncvsyEpQUfRcuLL5xMQ38vahA7/5mMoSSTbgwKfvwTZwWlJhNnCS7RnNw
SceH8qUOHYyTuX/FwDi9aS8vHSVxB28rd6cF5yZ1I4Zv2b8YnVDwSx1jG4XoictSglzLWVBdcPPu
Nvq383SF4Ps+tYS7BdXwPyNqbCoowa8TB8deT/03YhAz8UWwzekfFZEwK+GH/L5juXig+2miCTI2
DRfZuxDhJyruC7ETW2C5E3zF0V4VxQYFP2B7f/t8hfl5BBUoRVISdHPtS94uZbiByHXs/FaU42aL
KgrNBHsxm3AZZXpnB3e9b8Rps1vrAsDFnSFRrLBr42fURxW/9X8vpq+HNRwxB/fVTbueD1wW8NQP
7gHrTqcTu19d9CrqZadRHor9DuOjomitLXmLxfuBj49/QLDjPkjD47yjXlbJR1bm78rQV7Dux9b+
h+zFGP2anG5SMriMCgjXEf19uP0gy++Nv003frseozgLqHPfTOc4Dhoth9CvFDVSHFf1Vkm6KPeL
dLCl8XwoXlh6snd1KBWwsa6EOTf0FjMMCaU3YwnmkAD/3nMrMWyUine46BaPwBPXVygznStqirsZ
2jNCK7g2xIglK0DDY9aDpb9HKcnl4Z3u94RbyBBZZCWqlXGuVAAR3rTn8XLu5K4PoOYTw0AS4Nxb
cbdHgWXnc5oR6Npu/3wq6YaHOcuLEqj9rCcIKF2FQOO7G1HWusYh28EzqJAcRa+0VmgpMqAKu93H
nokCE9khho+JDgdkDjGAODUSUb8KKA9AKBg1kFOrz9SJf5UyCQukUv8ElKeBIqMQsjnPvouzTT3V
dQsALaB24XrNQTWcPjqti6jJ/CT2bDQK6PWP2bRzfc+joRQJlepkCy2thZqlweku2Hk0Y1v0r1np
4Mi+ZXJ29219dPRp8yFmliEKfECClQKf+5zlLgbtDpgE/7CrJTRjh2IPV7H6SUrDiYB/2kG50lX7
flGvLaXdDEULBdV2mD2EPejqBFX31qaBTB6YraMXJU/Z3xfZkXJR/vIanD18GuA7xVjedP0m+Sy8
avV1oq0DJftdBxkPIxUN8xKsAitFGECZQg8baUtZ89UwSYM1NW8k4RVXL8Ai9isFDH8ah21NX5yw
2eK4u6IcQ9s8XodahGvItPy29mIwg+iksJgvDUPUrKT8RfpWWsvo3OD3kUaxhQTWqQ0DMNTBaUVv
C1pHiMb03Wz6Sy2yieN7i04lp5srO+IQtr4SHzaNvXU91BAmvTqZAQRaERl5s/73oeRp6AIZAUDM
G5qpEml4H7HYYspYwchgwGMqsHsZodPMAmYeAEs2urCw1laVD8rXS0wCZ00pQqmHwoXuECa95/OW
O1rMMX6dR15z4qVand86/svmFcfO1647c71QhxF83SFhZvvJGnudXQL7iy+1EVNDI4QgW/xL2IaG
XZ50isWjWHz5I1aLBwGAwRjhwyeJwtwwCRRuFA6kSHSPnq3Q6aECmFTidyNDl5ecVSBXUCohLp4f
tFdu+uQInAdzmkx3uga++ihVxWT37yIQLr87ON3rIC4HvtRS0IpX4DSKWSdtMW30p1bCnoDvPzzB
iueoh0gPBFqiZeGXmEODExBXv5rUF/DDjGqwPyanboISVNz6QzOJD8juZSj8h9sMzhlF2mi02+Ir
YMW7UNxIbNtzLnCERySvrPAbicaCapl5douWPsKiGjDZ9EejuDb0vJRLa2g9UuEI7zeZYvhhUP7i
foyxnwnAJp5rmU3OqrNcBFRQuYGjABJVrVAiDIO1w0V/ToU6/g5U+0LkJCrCnYpEOAUvzuwpe5pr
jz1tW/uMN1auqMcJir+sialq0e62SRYSF9bVLpTlTJJ69BrFdTiMyJlVbBAc5vEw4U8ZcZrucXy4
u9yd/RLcN1R02JGHWYU2EHOuX0rrIxa8FrRkHXLV61wcxXqIRlhvmOYXCCknDTHVUJ9/D+nunC1y
tvtoadMXgEM6sMCLgUJ0feW2DVOjr2iNtFxdFN+UCAOtxrQx2QucB0hiE2tdVfzvDPsfwFlLvRA0
5k7al4rGwGCjN0eEwllN5TFQ6LFYZ6CdK0n0TA4GBaONJC1IxbuRcjFmLu+HnUXa8BmDUn0/npi/
aZmHT2E3QW0a6DFFNVHgLuG0azqN/HiSJ4xXmGcyenL/vMU9tmPD7PySbsSb24280F6DL8K1Fsof
ACsHCkmiNgaoh1kBPtIL0CaQm4n5gKVWgOL19o7jLbKOWBos9Wt27oUMn8ZpYcbxCiaGYOdeEacd
FCNUu71oQ+zGNo90mkkgdr0xyUGRbdYf8nCH5PKmL7+nDA+4tCjbWKAc4uVLJOnQ94rYwow3ni/x
dHaSDvEsTMckyWoONvlPXSFfsNc8DQVjGOU+NRJaSxcN40UK9Z6rJZjnbKbNVN8jm/enHAi7qc4V
mHQvjVrTENtRWYa/BH4lcbcgHkmitwYvBEGucf1+pZRChNl7lE2aRd5Yh0xjSs6RMF2YDBEUrx4B
i0f0bAwV6ClLvdMS7EXp95zbUtFn8KKBBtAcl7OLN4DCVvheMdtQLuCMADixAL0aAmExDczQxl3c
VS6yrRqNW/ECvGbTU4ng5R89y6blTLKuC0i1eOpZGYTcnddjNja49dNKDQObEAXyP6W4SJnYed2R
6derJyKONSj8uxr0vTh8VjF3EBxv15ajM3Uy/UmiKbW0q2v7l3DQSPlWT1+pIpyKXCoGk/uDalbh
/e2MCUSu9fJY5Cb07CBanEMRNLSHe7LmDjPdfx2n7qibAJ4u17GJwpZndo8EnufFX63z7wXslD7H
9qBxVRfolNJXR3scQoGLuZ0RCYPrm5ZuXUaPOpByu8jJzX/h+ERsKwGhvNvEhUfJNcBg9NCiW/sV
D8+4i/L2WuNO5F9GqQ6pTbJEESZ52Yb7U7tudpeBPS57aF04/mrmvnCfFvcCYGe73f61uCeNhSG0
vEmGvEHPgrNf3KjEObgsFojJ68bjkX5mZ6X1yunp+VMjSYKzW38FpQQWQWJGc8dJ0sCdIDkyH9sx
l33ywSbB0VZ541VSagqWftPzaLmQvZ8MHQQC61SjYCoqR2mbIhBcKTF5NlCq+64D9nUh3bTPL3Jk
JdeeyxdF57piIDGdUkyzOCDI5bR8MQMA1OCbuZ+ZZRWJiYhoe9B1Mkhlegisv3W7Gl9bBvADy1nT
546lG0tAk3ogJ+4ASgnndur5+8baPZPdEd6x1Mq07ZmGKlveforXm6ERIO2XtgjRctGeIAznRzw1
bzZFLGgBo3SXyt00Qccj7JF6nyQCkdmN2pTqDXtq6411xswWHB/XvtktHWAXPYCrWfRp60I805En
QMjChJ2QbMKyffhtZMmvDcCCMIUd708yk3LsNOgLGvlh++WThTfSPoz7tIB2QvAdsAqw1u3Wieat
q3/2cw/v8516T2/bv0Aga4uZsIBlnzdNpyKldHRJgnuTz8q5cKbEoKeUhZkjusublKrnGOqiBmmb
NQgBi3Pfa2La+NnghFl7GU8yPrQFl5bSP5iMpvCh65GaUoGKyd5Lq09Vq+8pA37PuXcq+PWD/YaR
RvsR+Wh9ENwZzg9/BZGpDxtU2H5+md/QuDMGaHT2H0EnJyTyg0A9MyTzUXupg5ZDaD/QJgRf+MRp
EZVGalW6V/jesaMBioJeKQsyNXMINjltHlY1fgGqJvRu9d53wdwoQtN5eMgVeCgBhyU7aNS35TpO
I03NchqTfPWrKc/WIfhFDjJ3zhqYKHmJoV4r84XzAbeMkgScFoC2G0XEVfEcHlp3x0rRfcweJyJh
TeU+l4GF3i4spjjfRgE41OQhQxc5JGpY5vT0cCWrs8c7UX5Vfm/LKVQj/L98i5un4kOBXTcPqB+S
7Yririya4yrA+qek8vynIxT61nc/sBfKUTo3lmuoiNj9wgtKDLG5KzL1TCw+U6urnPKjhCrMSndp
yaosDbOCwOeengu4+NkhPWx4wfJAoTtPTjBpsVC719zppCcMAs5PzS9BrnXyqEvtjGO9czmVtMFJ
tHvEVYNFp+dhmg8ds2pb1jqjnSmGQbPfxGdQV8sX0w8+l8JGhvkwb4xo3iTT+Ora5Ppr1mvUh7fu
wSKsHd6BEHxt30p1mJlkusLU1m0EhWPq2MV3X5TPKUuOO6EvxClYmfisxOJE2dsKJQbRAuy9I6Vg
QD6Gd9jw9gEOydHtShe4pDt1e8Pw0J0tqz6JdD4j2omMaXHQNPYs+gQxIAmv1FFMSURyU66QMOt1
pIfLNDOZzGgvyDeSwBU652j6wNJGAqIZTVVPxtaaiTlTTEpbaxriIe511hoMtWQhPfzYoOaILFx+
P4tjNNuixNqzmJ+tKMaZRfrzCh5wXyCeryqMFQ2cWHhh+6Gj+c34YBCkEqlXOVkpLHLQAqhdXn8d
YVWyT4iAEYl3GmrQllj9Ar/HkaLcq0Onhliq4JLPY7+iZtx7xCHFlH7EcCzxu9VtelCvC+ngR/9z
2Z+1FTAW8a6qVqPnbVsZPdCdI6AYgisfPbRT/HyN/UDt30Hk76cP5UvVA5OIFZg+W+72Y3Qg0bE4
II8WGKqhTAbz72/u+cC+NL3Y1baxXwPst2lMFEsiOy+y8LUDsMEKaXc3QdHhZKWrJVtNZu3ce40o
TvpGKrMsAfU6HSN9QPwaqcKoen7ZWXecZCygBCUoqOQ4qqOwXT825W9vnAVy+y/UG4uanhvkeZum
8OrxDGlOodA/sNf2Ba1KlhMseB/GITe1KpRdaB3o5v2UGUr6du0SoysCfadu2lRpHO9KLUO2gR6z
/GLHnMkIVwoNiXgI1smLOnDXgBd84hgSX35FYToKpuCKrDMzVuzRVqCYDWKcDOXenELY1nMkWS9n
nQPExzFLnIoLlM+6HCEunWkmISNgxAcuW7730xz4sF9A81XdKPkF5VflqfMZMmQQ02nz2c3T9Fxj
Qbl3BUJkC/A4TkhSxPphxD4MZZEsV4W1zcspaLe28/7UQ8J80kH8a9rECGA4gqGb3x65TUdYQXum
0DzEwfW94sbLS2RepudO1QLoZU1ZD5OQ5khzfeFHfUD+4GUyBJxWPxH/bARLiCMn1QM7jO4JsxZ1
WkkhyeSCu1duM7Zt/QPYRcX4wotv8xs8hEkBZSti3qDEjOeQMzcJB9MkLy+PtlSbHSAumWUBrg9t
zJSwbfZC7NSNGhBRfsqyApQtpIzHRqb2uCncrGyt7y78ukCMBx0l7C29sAVYaG12cglHeACY55GD
3TGteeYTG2VDgDzRM+dQUxfv6kpGSHid60y12GulwBtj4cDjtKaJDr5qvUzO7Z03mKOOkhHQ4kXa
7d/+yM+k4L9w/YsYkjeCuPMbGXxp1mFvwHmZiGVYW9rwtDNhZM9Scu2NW1QcBL4jnmK1aAyed01j
TQUJv6+yM75Gwg+DgBfmxgVhskgNHPBHDCSQ3jhk/XCBz9i5tz2Kj69dBH49WhpJr89FiLJcTPA2
SmF1ha/MExurEyXubp4lHumBmaKKAA9aibp2tsg1nBT/oCRAjADuzYw95ImaPPavOZeeljH4MLaO
+rhkZhjSv6vQo/UkvG3+pq/u4RQq37MkhHOrLjctuvQ29uPw83dBUdc0xr7Gi5+mw44U3+yMqvFr
DSEn3ZS/1bDe53xIUJEWY5xffSMPs03AnC3DJq2LMKCG+oSnCm7mN5ucJ+mT/ZquDWDvqgAB/mw9
XiPzmSPT5SvQ/i9gxfxvVrVwU6HXiebMaSLo7UVyq5t9rq13A3qZcmYsS8uypS4d6io51Xyj25L3
adKn86z81UNpVltLMihiBukCoE1y1fnM0rRL7ZY8oouX1xSHz3CVGixyiMGHD9B6PC83CNlzfzca
FGUB/p5c1/TVp+UVDbYodEiRT2tMJ1XPZo/arLlkutj73eEuquFrPnLU7VrINieTrFUodXqpKZ0w
noK53+hgq/7ZWjlHwuCyZbZM0chllyJt6rmZrZkRvkR2TeTcnP3FolxXwWZhHGU8/qz4cm67jVcT
H6kMgnrTkDrl60M5MnT4H5PJSfaA7WiAmJILxK9dErxhMeTQZ/zlAvGe62cU936dwe7Su9osVP7X
K81OekQ7U/Jd5Fk0rB1HepfN10gZvKbh4ucyRMBTaVfSthKOHnT1eYwC7fwRwR6PCz7RewufMCOQ
ypsLZrHiICIJDn4+R3fRy4Ntx8gcr2XHF7CHoo+UcW3v1LOK3HpmxmJiEh6qcdN0BTWBLvmEAr3t
QMO/1hkPDOv7CxUsPd6AQKEofOLDrYmHac7eXqY5/zvRfbYKfsgfmAwySsOtUumc+3ox/77NM52d
4h0B22Mo+tKEd7mJs30LkYHcSp5pyLILtVMci8Exfd7viljTlQj9l6blNXM+jDm7YoGX3UWt4jOx
M46dreTx51UELaSfZuwtzPAQzt2Fx6wugHQqqaFU/y3/C/CkZo2Yc4/w6l2myFsJnhwDhMfUZr3Q
BrPFR8R9F3taXGFR2sP1Dr2kLOjos1NnAgeQO9AtzgztOT+vbBdKZPZNmTTbnXzfsZoqQo/KQlxy
dsg5sFzyhcSzJWs4cqNjv9ftY4xg0qL9tnvYaJh24HYoro/Zbv5wVlf7Kn01q6GjOCYWs9hBcNa6
GrcjMNtNLMUghvbx0/MUWotDMgynRD870DPTs0ZaodSRHQPZhapAHo19LEgNT/rKOKAfPwZg2rES
6IS94hQJsGa81TAMizDP7ZlV9sk2BXppy/X5JjlJsZKjcedl+eR918OwJcKF0h+MmOSfuUhZ2pK6
tvAgFD5eM8QdqvPKec6fvSHXSTTqsKP3lrbQI6XzDw0suwimzXfLEk4Zu3xW2KxyX4yoI0t2lO0L
UL5ZoTUrN8V0XlxFS2wZcu9YyH2YBRFFq6SrGMTCaQUbElH+gEYLGFpjUELKCeRLZ8TYmCMzcXwP
M1eEqL8vx2szWLemhW5pJrWVKr5gYYme8TQEdNLKyhZNJ0jkAW+uL/WGYwFHrxZ/NfK8zCzKERV9
EPijeVLx3B59vfMTJXyH2SioJYjySOqueOf6nguD22HD1d1SRPQSxf3uJ7Vw5qT8xgCpPVvA+nWP
FF/zwnXkuC7Qp60P+TnIgEhQWWbLXubHyWWAgqO5rJcSng6CE70Dxmrj7q0sQf1sidFoAr3rfBXG
hALUgyI7z0e93TOCGc5uOFco+TQ2WqARrE3/kGDl2cguCwTDqMJ9jPQOxzP6W2jcC9aBWGGFR5Aq
8xHVNB3JHFioQNZbgdAKFfr1CWoErcAqVa0X/hOJhlPNpSsGZgk+PE2ODIJPc3YITTVPgNgTrGQg
4V7WZ6SWBFteFyV2ooV5cSwsvrIbOisByk+CDLMt3ctOqJUEM9st7YgmE9E8BB2rl9966cwVDF3I
SWG9j5evSKdtME2jcXCQp/ck7zHo0RB4W7hwuNfldFTyUaX43epcbubisb911W8LqEJp0KmnBvHU
cHYPDVvFI7e+So6BnUjtfxuT8lWpC0M+W8GmuchQ2y8EWChZ6o0g0UWVVYoZJ41uLZy0mOc8Y8xS
k5yFmkqz0GVJFnBE9tlNHB0bfBxKnV8Lb92ZLXDLhSPVa8UFelnwy7zKcGqy4ukOxQaxZQYaNaBo
4JnF8ta/nuuwyL+2Jfhyckc0EtOhZ4gxa8+R7wlQxUJDhiTH/E2bn3CTdR6ntTYh6o0dNn77fep2
1uelt+p8CUqr1b/pdaxEpe6OujQBNYSnqNptmCggp2/wAcEE/aP3A4s4sW3I0KpOW/aCbBCImroT
m8fchfmLgLIycuNUrohCR1Gi0OR55WHIqGoW488Arahz/I9rC0YGxz1UowGMkC0jLQoVaIDTrW/d
raEtutm0XKhFv+jeTlAjeYdyIhZL+0EHnBMnkx/ATJxcVuTf1TYxG9O0KCT30OH4PA9yWxN5qnkE
cU23+DsfuPtj2ERc8+R3i9oSw+Zeu4xEHl1RoOtfB9w29fJsjv/qfOByt392QedG6NrREt1NDWZg
GvulutQRwCSO2VMBTD1TAQ20Hq3hbjsjdY2Db2AW4RrFZzHctZ155PW+qfbeyb0QExMIcuqfSe4F
/nbol1R2xxKfiTKq1Lz1YSRKzLa9YX76T/ljmO593Ez7mBOrKExDptSm7mS3umqFZngTC4nqQWKh
8G4qPeeNJ2VooMo4yM3ojzz3jyKzMgqEMKh/a+sxDnBjU9lgvoqKEFlA39KkndKT1LUaszc4I27V
qEZkMDlwNxkLJ78fbkYznOVCk2LD0IJfKqhrA//RQeEDq+V30gB/tnC6mjEFPslJ2cxwAwU4OUa4
lAWHULLAqVN5aDJus3qS+AYMturwV4W4a4gt73sva6TCrqKYg8UAxRkX2MqUgI8jXfKCZPSw/XqY
gOlG5a4MLVRfUvHAyPi33oZrv3eDn6y2wlSfhbJV87uOmpoL8UUu/v4qvdQvUbc9W7lr/xtLMjTi
a0viDx94GBFNCQZEW8GeIhDeO1L8esmO5pdlQVmAnzxPwYlfP35EDdS2RybagvdoF3BxsnO+58m7
CzFYHvOqhDxQQMxi9rZ5rhaZNYuNxrpNrIMol5FLjoazAzQqva66ggVGnauFFRS+XaexVV8b2FQM
AkA09GwKI3prpw5kqltH+k9ejMqz7GaOEpg1bIDONM4f2CLLKEw2vxo3vEtnLaIPDHtJpx5AcAh2
JlDeGrebBgs+mED5U84sXGzQ2Vt5xnENeQyhzSB2CM2oyp2wEiUa5A66QgVYIpZZJzoobFqI08/Q
0XfPZZybHVyZwcOroR22TE4+BOPybcxqArPbo2pDP7a5DLz3286dxYHqdRIUJxp91YifKl6T5OAI
Vu771cLhgNxo9rni3C4uSMe+JBtgEEojVz6lftouz9XnoI/pqCy9LLyHCP09H8U9z7MDHoswGj9d
glTXl+Y5PcGRqQJ467mWSnDMm1/lwKiIZSxZbLzzje0HbiveEbLhWnSVIqaffyJAfa9X3xAdLD6s
GJRKC/VXBkbiKWv3DCykcxrQYm2WXdN+XNJJII9R7XAYZpcvuY00u+RQvMJwIhTHZklYPKvN5pds
ubT7ukofXe66DGnatpvYmW/mMgh+9kU35maUAElDuFbNVnB/kD9W0FNQ1XaS61K2HY7iELYwed5Z
U8pzD7uBAzjx12HgoBLjIw3viPB5H6Ha8FCP5ZQySjayEcKJS7U5RmRTU4JqV0tQ8cx0eC7SC+Vu
sLggdQCf1UI/s9mckAGeMkqlR35lX5WaKy+DBJSXBhcYCmW+lTeIQG1ovqs219jQCclTcgZGgdwH
b38UpQgt4jstxptQmhuXd/4EV+ISR/JSrhQfwlUZhf3gn2dv2Vb5Wk+2ItAeu9O7y9CB0zFJva2K
74Yz7lfOfNUMyFTmRSLepRMcrKBFWpdFI3V/iL4nxcbr5RH1MoWhqxWD4W5gCvi/zpR3i8GW875u
1VAH9NIg24VE2h4Oox4qi6K5AOCz8HmEy/5+QR4E4b1NkKf/kAsa6936NRbkNmflflKV3puw3mpe
jvx4SJBJjVpHMQiWNyS/UN55/g15nkVMLgLUpFsP6x0gTvoy13mDIuSYNWrUaZKNqZT0UuT/RlYP
ycLCXWplVISu6MhlycdhBPF/t1dJdmXPIsq7/KONfdZ0Tb5xbGW9zSg+iYcBneC1VB5k4q/yXMzc
QXFG6WjI/Dr43NZVTTr3MY6XYCLfWdN2BpOQmMKvBsyyUcOvV4LXZ1Mg+aLlF4UfDkr6QrpMtlpF
9cBmO7zBWbAjNfbeYGPoXKRv+EdM7JnxvXG3yq7g5Z454I6Pd27rFtF/7XtyUz598drcQYjJ4y00
FeBcTq7+S4yZbj3ZdTICz2vcYmm3kIe3gID4eRJyr7hLoVbByii9U42bA3ReuzIgiN5ZWg1PgISc
uYGmst/UeN+VsS94BIkYSHfL0ppubokOOczeHMvMC53rAAgljyNm4FuIfxO7GbvlHTKDbIaxr1OY
8jX0bdL5bD9o0CREUtzgfwfZgf3KhZx6gsxwKjOZ0M59m0wEmtMw7ecVftHYL6SrWv6TWBZ6+Sx8
ptVKb7OnohNAoptsIliB4TyURMvdqYfS0UXxR6VL8EtboWqum0LnuDr843XEm45O4m3o6LcfJK2a
/6wbG7wxAz39R/K6F00ZvyVIhZxJhV4pvkX1l7mzLMZ2mhhz09By4r/xFlMEHlPoRapq7ZuksUzU
UFt7Bc/irRgXRsJ9tStrWR0NZzwrKpv+if+ScwLgyHbDZmvO2gstzRymDKuRwcXStM2RLxZj2h/I
IE8ZdpycNi+j+v0Fw3PNz4cOl+I3Fsk2cUuUNx5CS3ZDlCeKJsDlWB1cjeBNglmvvDaRfQoTU0N/
3Dv7ifXT6p26Uhq0IYz2vzW1AtlHlaaDx59QAVJne7xp2chguj8EAP+da2xJJNz3lk9C+N2CmLQz
TIPv0GqJFdp3YX1XYpY6eMYmI5kxMxUPI+tS3PM0xV+VIPYKeNV01ZoDycqD8YBJu5PHibUeLWg3
OLwMHzD4BpL8MOFvXae9Wk+ZJj8BpTtT784/kYyUyj/wNMdUoBdGrvFJpo6KbIRHSoKUN8RkvjJG
GhaJw06/BNmlRemsXAzrhceW1ekEJrjsQCYQryKHsicWeev1vbiqbxi1RCOyGZyID2AR9rRw152m
twkdApSCeFRzlm6coPivlnvZwBOo0RW8aKkEiHcCXKcU+PtLIsf4JCqXjqaL8W4qpTvEgWjCRA9c
7YsOlZPjFfa/7rQTrBlJlG1CKWMrDyUswWTYGKo6GSB+Eb2ievSru42Zb13DflrBWVdQPEv6vEql
ic/GxFxPucPRxx32hz6njGCOeuwz34Z1eefXWudRmvRz0erxZ5ZDodGeTt1nVkQjZd3V7RNykgXa
d1JrRhRehbrpGNCtV6MzrDk/PlJrY7KSZMqgwbpdLrgcxFUIsnR1suyZxkPj60dGqf8VhsqYDNdH
6i0mgEo2N70sZ8fkdCgjCo/Mwnd6Zb2bAPczWEGQOl0po70tWkvHZmOReED4zextMqbbymowMJLv
x30GAxyhKNs6Ngdek8JdXDoKC8uej3RQDzXF/ro6cj+OVpNylrHNxpXXq9+MSR/Be2CkumBytqOB
1AM5nu/1B53Qj4kx7O5AE74r8PgLToyazXkOU0nNJV29oc7XweHlCuh98zb9UQ5Pf4vFBb5wNKrn
3Ax0uXz8Dhza1JS6Hft0M3ejLKKERPmmiqvu2wYjO5JF0U3S8do/uO1QawPQBIbmTXGkOzPcWFpy
WJP/89t99GBSMckJmW4ilCyITjwQZbjCTl1YZGm9S3hGxOSZafw2FQhCCVaLFpV1uTHqUVk45pw7
U1BfBmrNUchV6CBeMYCzr/QiRHx4S9WgTvYEbXNxQShK2UzJoIdV5zYGZLVFdTIfob4BIO3SrrPV
7L1AUao/oxqhqApsXYLf0io8MjubdZJSRHMOjMCm1q7rUMWTPbJIQTHmNzorjSYRQSLEWdSz3eyE
GKAMwab8ZNpAncR2j3nQ5bEa7BAxJEj0eprmEUISccF3h3kLYdvs1w5qP3ymm2tjYDTFaHeQxPlc
7uZCVGyOO3sc7g722F6V32QlXHDzuUf2cKexwgxVP4AX3L/ZEWagj+6gltfEs1Nn7h7pAeNZM1sb
oJajeFyi6M9pfoVOvvNb4vymOmGovL8ODoC8zsu7QM8d8pbDMLXbdytFjhQ7GbW3523p6QGPZBav
gUl+6PhLmWGnsHALcTwR8nirtGcpI/Q3VpLgSkSTWCYn7dQiYCtGUpR9ybFA0QNDsDO3cpg6Q4V6
U35NOHJjPxiAA6oB/+ZC2lOUc97pe2BPtyE2E1tHqfn2Qs6dTUYqV9mKrphIcfQdtFxV+/302Uag
h1QzClxdKQczwmLj9o3I3amGBcuKkYmIBgvwSYhs5CMAcis9/q1hJ6YaPsQgb6TuzmtCUQlmGXNz
RZH5fx21u1YlsC6NROrDD457MJWOhwZVmCYNClH4QCk0NNLYyFKtBTHphegC0G3Y9/OyaQzA/0vl
OYoKOxJv3cXLPPtckCd7VG+KU7CfepU27Le/5Iwnru97L5dFn/iy9PZa9IIRDwIzVr7HzU0LbmKo
KwREw25D6iW6lMljzBgxW/Ydy5L50IN8LiVY6JuywsEQSpehEISHgCGE5XCPsUpH0QFZwB+CzAIg
fzphOoYIXBGIBWoIA4v/onUM/U3AwR4opeXwgZjRvvAlR96AcaEShyNi1VgjmMxiLqBP7eyZK+3C
oW74mJfoQ89VtCuz/tHzdPsTN6/BRe2CenRR9We3zOgO6Ks7Q5GeC5Ushl63Av2EYZSGx83YkjHj
LMrHfTzQTE4BZBnaf2YoG13JCtatyTVLXuc5MEkpIbWjZEFfhZdBhlSaGGkgseEazyxVTq2yqrV2
jsQXbmvwCn2EIEEoI9VKxXp3D+xuGzEieEs/IeMNHh4xTxZz9uF04xDbAsWABr079xfhaZRPkQDo
+jkDQL6kG8G2LnI20SdG+l5ckSIbYhyrSZMlQEEs5WZgCrXMEsnX2XKK3j1NLLsNmkttC7GOPA/M
5iBnVv4o5d6wZ93HBkaVBW3yx5HifbLdLD7qupznZwPj/mB/BuytHAEmYZd0SOOTNwJy2/w5aK/D
np1ZY3gWR8L0PlmLrYkxf2D4g9/Y8gUar/t82P8i/8y8BgH/Fvbf5QzA9uRI6zpFwXeorNqzxmH5
Mb07ZzjaCRkppL2QQtj9Gp68XIybOmVLvuzQU+Tg/lm2sa4xx/etJEETqTmBFP/4S+mNkWQEuNIW
2O3quaZvhS5SbJiEb+1VOneoT0sG1OD5V6yWPEs9AyBbFoJ6+uumz/fZBM4ENvyu4kCQ7KIyB5Zb
3ngocAsSrlg/zJ/2E1yr9ZXtEzmJP/QUt9pfRGK5pN/tFHCJEzQa1a6vOm3XPaMwvRZ7dY1wK6gt
OFC6m6j8eC4dKFFfhdKSiBCdRt2VKH25UHTkxDySDvga+wWBg6wQwI1Lq9lQ/vhdwrdvbouyF56a
Z+Ui030t72DqiLrgNzpBumA/V+ZUYDZJn6HA+AvkHA+sgFcFHW1W6wxcc0fmp4swSP85kDROJW5E
E8uPnu1v1d4VIP4Qb497QoKjQXJRXwWDpR5AiBzD3tCHAA27V4DhOUCtptCZxtYBzZK8q2hF9Fjd
xqS69GvQiFGHqg/WljTdV/yP9totwub0QdBLOcXeyezzk308/GbZDoacWTHwLjCjwndYgmnxvrIE
H5Pj81KTZAbnEeyzWi9rzipWteU89EXO2CxdaIfgFUD67RxICdryX3C9PKZP3tYF3KXP5suxVfFc
NW5lE86B9VYpw2YN+KMdue1Z3VZLeJE9KoK3SmMxPROAog2DNMJdvt1lIg55pVblzQ4epENk8b8N
8FcqcinqqJ9zL+QsEMwpaSpBT4+C13Ce5tdnQUXa8rvB+J9Tb4P+A/4WuatlWSFxXwYgzZ6K6rEh
z8n6+E8tCNjSRKH70VAEEj69BAttZSKjHENNq0x2WvuUm1TI3vU5JMpzDnxiu0EW4lB5ikH8e2bc
R47yOtL4kEqWthM8h0qB+xnINftop+vZ7/KkZT7s+7CIZsl94soBOUdIo4APb6TfCTYi5OPCP1Ym
DIh9ZmOghiHtZyooXJNm0SBDv2lL4fIF5AbZgCfEhvWqFENm3J37sSgrY7kUXKyhCNeygMDI2IV9
1OdiR1EtEeP6Nh+8F9+OI3fVOEY0Oq2yeKswaeN3oF6BEgiEnuf6JbGSnWdrGR1ZqLi7tW65qxwH
Ik7Z6areC0m2sZZAHAodfOGKGI3aXVSUY8p1qY+3itHginmLBAA29FlL4LYW8cbDsVgbT5VOlxsH
FICSCUzyRyP5eHwZRSgDn1WEgVG91XtD+y0LMpQJouMUeXQwshTjP1oTRKWQsSaDrWEzVueRmons
WBlPJExz+U1u04BX7Ak1AQttaQLwi3ZmJDTuhO+xu1t3WxKFZncvG/x/sNS20lMsf09WeuCa8oRo
b1RGkPmQWv2GMpJYy+3oQF04XnoyYq0/IFJP57ajJf23Qoane0HyriUQkq4OQ3kqvssSe8JgxdcE
LWp52w0rRsaIkjysPMFheh0rAp3DTgnbhIBHY81RIWXSuqWFTLB/IWBYpDFuL/CKUGKSzbSl9PzG
KZj1tXDwp5YxhsZGFb60xlNQ/ZYMYQhsDlaAOtjhF1p7GgiYk+6y+DjX1fSPIYIWbdQhR2H3C6KV
BtLtTPYYi2vJoPiN+pseUTEGFaMIGZINgKwxItNv6Kta6Flhd/JI3vnGzi9vWz+BAKuNU+uOb7am
E4IVq0PKmMH8s7YshdN9c8j9B2QnRlWvEB6LRVHr9pOo0zIFf0TMqHRwx5E5A5pVCI+/Fd2WKHIH
LP1+RvQqEGluxhtMRyqNjVx4ewGrKQDsPvqEmmPVLFrvQJmQCtZ7cXLc+KcufehAiNoe1MFzWLNk
F6PTGEhUWYPJ/RCbkAtUC1HOI3QtIS57RmdiRql8PKQD66toWD/Oi2anFx/jMDdDJn0n76akJcwo
g99ayLeWRTZCvQBofXm5KWX1OymYKZ6KbOfeCifPiMkcoNIGE6ux97+0Rm9YGLqgVf1DUxZ8xyLC
g4M9zBXr5jqEsUgVIavVeMpbXWnFqlQpKE50evCOyRwSp1YW2NNYA1UIspm/N4qv6ySOkgnK5xL2
fc82BrU5Xzv/ZTxyfO1GWADJbH4oIzLTkI/fDSvro8beo0OdiiSY064Jk5adRaofduATot2p38vk
9alzITHJVrGonQD3+TsfvjmIxgAPZXDB7F38SDndpteN7lL3mTplTVO0oUmy45etAC61J0OHtxMZ
IdSeciLoFqw7mr04CXT9SHOVB1hvvn+QXHfz1A8JUoxzdcU2B7d15FmMtsoBe6ktAbQD/YbHghmi
SzQPQOsMXnQu2SbiMKZtooClSjsiMKfJTuK/BRjw7zjAyjxC8kiTc/73l1wbckIcaZEY3YFGYehR
FmuW6oe6zvJtHNYlDlf02gydfRCVYYfl3YRQHCDAWbMSroKD075Naa7H+dSxzCeN7odSX7umtK3n
mtX2kdazCcc7WOOji4RBR7R/9n/IIub2nWnjTjXL+asSE6ksCa4o8J7J4ZJK9w1W897VdYyMAyig
dJyYhKHpPDazNz8m+fiyrG77HSot39Z5F60Br9mTsdWdCvXmC25EZdE68oMAVsRJtLIEiLpAKnFq
uG8po1L6FGDZAk8Mnv0zQKaV/6YnH8rkxaUzERb8Ep+L3CGP00EP4Yb11MbxUAL6787Md1m5ELa+
CbrJzlSybsKoOSfvFW0rYFJ8AHeWntKbF9EveJakk+G3587Lm4YlT4YnUdQ5ovflGbP9FDqhptm3
TfZVCJFtCpJd1RhqwyJurnDiEmDjSTZ18VmxyfAgiLPC/AIYJfAz0+NU48bFywbhg/hwYQcyCrbA
RiSpbiiciEC5+kT2sTQGjuvg4/HNOVmJp52aZBkB+ekKlWmp9RJo8uUS0qbWCpZm8oygLvDoe5/g
KtYSQqVgdSzhtwVYrSbL8xV4EoqnoGeMkshdCBTyAsqJNlicPxw/kTFfToMPN3CIAUaqJaeaz9N/
eg3hB88iimyR5dEcvt7c5Vnu2QaN61a9vTlh1OAu3TAhd2m+PSbjY0UglCBEKs8yPeefioNNrXsf
u9Jk9PlCNCvvIVUvC6UsPT8X+WW2d+sqK0WqvFhHlSZHLL/huoxEHDPRpo754+sfs2WgyhmuPmKI
KLSW7VPWa/B+6erXXZIsF2RncFmW024uI9y80CBe8I5jv7oclL6UVu9bT7UADA2SiyQjgmyPRDmY
IwQRMVT+HAk9kfgURRExLA1GzP0vFKYg0/oysgzsIs3HJJgLj/4Rk+W83mT8ZPfpHMKROicXJtuW
wPWrDnrQvVF5CmTlyNuxKVnUT+c7mS3yPmEkNcn2YOYdzW4N5eOsVOfuWTRlWOhio0be5SxZlDHt
UYEhjUys0X5GTti40J1bXJ+YO94Mbj/CdlSpFKKfF6ihhBGaSq/zA4DxFXzbjKPyUf7kB7El/V0/
RuV5WBYBK/6kxXWYZbToCMkSvffRX10dBZjvPZ7bDE/m8hsINgQwubYlIV7id9ynhnLefFQ1rnSW
6DzlCZp5fQIXSzceCCDMF3Q9RNapW8omI7WkZtHkyaoZsCojaVmXzomONCSANzDuA39AcmZcLX6b
UP6LJ47pwoCnKSLNO8ayNa3qS4vDgu3KIX1MlKXNYTzjEJncWNP3iQ9qJ3nPDW7JPvLRIHvhU30u
eA8lEhmTCv63xmnvEI+1/7fd7Sl01zn/cyvtoPXegaaeMyXZiA42d2+7yno7+Vnv7QbdeQQo3k9h
hb0MzcTvbrIMnFe8IMdaPdPu5u72b865rSJShBnARKSw1L0Ejk0jIrA0v/zQElJmIdKlFo1Zou2j
n3u7/Dlb0e3HYsXcMUyWRL+7nbfVP4zvs0+NOS3xq8Gg3n/rTDqrVTDWV+fzTYimWS7KvusNuYF2
QO5GWyh+VY51YcmFhgFvG94xSTIDCfI7azs2yG0LP2h+2/Qifcd56/etmCShHERs1zSahTlgc48C
vj6fnOJ1g/4qb2D4RT+m89mY2ag2tRPcQHE7rcs0NF2WUefyFl5uAtO+o3NXgoJh1oBBM9KGGkLC
/FwbsX92Czlm7aV8ly62/gtJNydk3Kb2Hmy5UVnCcuHjyF9It9FkiKgytM08pHLXAATizaC1gpCh
RfWnUE6yieJ1E+NzoAAD8AulKXlBrh3s/67CyPkwBlNDqpV7R20Bsfy3FChO1cDjWr4ANsWmWN+U
3O5GhN4nan7ElHmTN7/HriSlsrgUdY/IJBjYfkh1xf3Jtz2xkRahk4oyvNbLAzDZMLWR0ub0yl9G
PPwq9DYMaiJyJE96NFEfnprNm9mb8ej9BwnBOv5xoOZcr/xl/CspM47OHbDiEkD4bpW1rlfZsBBz
TPwVqU86JxQWcoMS2eKnfSIx6kDu0JkNb4kVlnJP7MW7EKbRkMt5c5DBxQieJu8/tjFW7+C+R6lj
qg7s+O7jdSnKoEWIb8giHfC3QZYnP3MpOQvynaIBVSJcBJe+CsBkDPZ7l58PehKr2gAH9Xx3IZs0
UjsMLqnZNvjE7amuQYZsX/rWIEE+WH019OXh60z22jGmg5zGH6lcmScD7L+5lnGWX7QZF3/NFUhJ
w7dLmIj4B+DGOaX8X+eDyagAJNsd1x0enfH2v1bgn+1op0Sa2rd+FyS1bnEPhdmtCK1jUM5H/fK7
ieorW7vVTy4Emp8U+WZXZY1bo7IDM3nDscBSG8uDeNQY0zernCRGAqVrYjzOFPD7YGJCfO/GIadX
3/Uc+hvyErdA161hA1oUfz1CGi6J8hwt1xozUEiKMPhzoP8Y6brTo/TFz3oilI7FVaS1qlga2vkR
j3yBhtOlCZBsH4qc4BKXHlTIoY8iOOzSuKCxWMBB9Man7OWVHG8LgA8bFS07zlbVZq+usb9el1Wj
bdT3kk3YCVygMUseIu1+aorvJ+t0kse//ZMSxFC4S3PyCrFwcNR4tJi5DFMNxeXXYwtp8OUjfmqk
ZBITkvurY8OCns7dHmt/GQrBvLQtEiFd2CvRjoTmN/3DAHDCeSEhxE1tWWH6ALzrdq0A5+X/ZKBF
SGuAVwzL1YqkKol2+GdXSbfZxGAKLMt4p4SJ5TzgvdNZ92MJ3cPWGOox0U5rz0AXUdT4QvdZN/Ru
O3qMTRfXAfEVSsKTi0CxY6uJY7e6kJIxRkq1kppIeY92SGg9AcGaN39VPUWxZD/noOwzz4gQfCg5
cxPtqqYVURwMu6B5woXifWYQI+qQysZSJbkjRjeN0WzCuPFR4ED0BrDV5srHCwbvD5EfU8iG19On
m/5LASorvvGInLvF+xxGQ1Rlq8Ifu1T34D1IoBXx3mTTLk0vhWJkGF7hX614RW5XuwFAy2qbh+v2
cQw1dOEr7Rg/kx7z3Ta7x6G0Tx7zXSD3CwLr78mqAJu00BmVBjeOWSrYxfrEGkve6oQQziqZUQBU
/dc7hqCGRKjldJKL7SZlUpIupo/chgUjEjzdQ+B4J120VkuVvYVP9QzROybZHi2xOP9B9EE/f0U+
rtT5e15mMh2qWm6y9RdcOCV1TkhUCTBbkIeNbY4NyQGhsdvcIRL3ypKfwVpsceFG8nsK2657eHn2
6fNQZLspbifwuy0z0F4I/gCCDJiRQ3r6dmtTyI6UwG50MiTgIFR4kRfmtWx/0dfOkM+lR6gNPN75
/O6y4ydWc5inG5VUTyNL/Bf8EybKmRn9eSW7HWt6asG3fYigDbE27BMEBxyqdg9kNKFD1i9lWmcD
TDeE8o/yHrnC9MOZoT439ueB8+ogSqfeRRhy+FjOX9GXvK2HFeGpH8yAuBXYZZwo7k+i9RHWhPPH
umkps1m4JIUk9PPWUhMy5qzWDCYjoYzMyOrlZWp0HJvGIkHBn8jAwB9iu9X2gPp4SUl3N3ie1CVo
lR6XmKK7OUvjyWjl2HJb/xnF1zVi340xOvoySXYhHfsBcmW6ugJ15wmHe/P/eLwbmGZHEI6Cbwsl
wZM1mGUXZgYgATfq+HjLNk4s5hzPIA6vZsJ4vl5KoBfSpLjfaEj3XCtj1izYKgxAL7C51FeYwIVM
NK0A0r8QKukABLPlXK//A0eI5FSpsYsJnCP9xwVGcfgUvkD5wwJZQL9RnAVFGwzgsW+ZPvH3K1fK
vYS/SdTl3P/oWu70buYkUJzthKD7SssjCs5+7k/RypU8CmKewLAicxqo/on2PTzwBM0gBLAuRwP5
ITnuUVmITHDt4hEwqN/HGoRqCeBC3eEauk493UzZdvoAUKS4iBKB6KY17bFEhdAJ4J8z80L+QONe
UDQkLB7sQVu6ed+Z3lH6HFZUC/E2snRf46UMhfyu82WXgha5ZULwjAwscpzd/xTgFK4odfzTg5KB
pHhL4rlp7g0NYGvr1TgjE2YF5Ws5QTT+c/yp9PJSvfEGi0NOglxpjvyPoAYmcFj26w0XoSxqnklv
qOnG6wBXhWO4VzgnVJhvu+NS0dJYLnapI7HvtKtB0fmmty1QyDHROwENKp7RuGEryAGMJAb8YmoP
hzCgpFJqPKo0EJANzPG/XvAI33UBpjdlQBiztXrsgbNDpGR2NspS4RCb8gNvY6v9CRzScnsyRbp2
zScjoDhsBuS80QhrM0tRW9rSpjooNlMov3VC6Uv7W1+KGurjE4brs/TkTsFdfR3XyYsfK3sV/54q
Hi5Ltko3K+zVmiXVKXho21zFtg2ph/Iiv2qJe1aCbCMtdcjnxAw4kQwTYqF2Cx+ZwzPOdGph2rNH
9qJehFnBdwzG6lTZSa0RmFmZfOHS/yLpacMFruumkFjDn7Prcjskuej2uu0xcbcr8O9UADNQLXVY
ntt9NZP/YOh8WxrVHiWF18ljDmYDOg1MvQL6xgRh4NohmYJyCCWeyvG9VYaQ1v+p7Wbq2VPkVZy5
eRHldW5CeCaI/HKObg3V7CDQZADT69IUKLLeysduNEzq0tFm+nf4xAKyIe/0ult6MKd7TuV9sIvD
Wr7PjtC6017iY+z2ivx+nzjCkM8sfF5MkQVEuXfJUxDhApKqvtKAgyM9k4XKQPP1JmHXipFvQv5G
ApVcDvIW3VAJR5ga/33FQ5v+WV/J5ST/Lz88y661XdAOZaKKjtgny3q5F9iG7Ogwu59Qj6d9rLwA
m1oaurL3zPPN4ca+rlLXJ+jH0AE4xdIypvoND/uO9P5m3JFhn47sEcF6KrgaoEamlo2TM24ocmDD
Ed0vMIOJOvr15aYnQb6a+9LKmr1lgTm8HCfIkyK3lolMzfsjqNK5rKLSrokSmqECWYVVnkoZ0SJS
FKEDwaO/DD1rb7mnu+m+naXulHfrLzWjfbM0vbxA3QnxWwWvrneqgEYLZs4lkhww2Cjx0CZT+jUr
HpbtsK9W1k0BHYXpvL9KcIuPtHZCOUqXqQ7YZBXbDtMe07Pzams5w0rHhZ4+7MGukzf8RR7WJEN1
VF+zKh0OrYwto5nmsAg8G6DiS6mnokxquUeqL+eY1v4WZwUUGI75il7xd4OL7O7TSmWjNMk6P9qC
CixOt0vqp06mdafARstBcw6eU+V9mEhCVo0w85SOsSbxuj1ZG3Ec0pECPSp7UZ4iSHzSjCL0A6jF
CGzx6b9fKqsFYljXcoqND+tuY1JHsRUcAoM778TDTdo8/ndYAh/Wwo8DBmvbxRXgwhV6PFfEy36G
1ik68b3bpVwaJhcFdOuGODqNtNBGcd+X0zEXOHDrgquwG3o5BwgpiYGfXuTgADh/Af7HV6nNnfAZ
tU5rF8B4LEErASx3xxpYX/0CfDiHWJMXElGNjFtU+OzGh1/rcWXWtLyNSCwj/gUSmkG7ta+D0JHZ
Hg2i4JMRCgOBBKDC0deN5KBFUwTpUa+UcmIUP3inJ7TkKnTPaexce3pNBI0bPAADprTTQ6RK2E0B
doM3+ipk1wI8edoX2NM70Azp9qGKFZvytsWY8lSg7c/HMNV3O8B9ouPa/7W8hxcbeyVqoO+pzhka
UqtI/3Rclf0rdBPp3uJNfRYz2HbHOlY81GcUnRVVh0GPr8q021LOM6NZbdBuSUdDxbt6JN1G0raK
VJpXnJxorx9J56/o+OGP03atwxFDyTNgdwTM7vkiVZbMf8mu4lwUL/2sjny7O7SqC3O2i5S2GNsX
Iv4ylvINuCvJ6SG2cY20PQbx2cb9wJldRmTGihZHsirM4UCh+8Prk/CXl7mtL0VqY5ewr3vZuGU2
cI61XZhxe0ilWCFtU/1qsg3akhFofapXX7rIei1nQxhzvh4E1FOdY8ZPXn9I0g4qzvOxGt6NoXSm
XtjJyd21I+m0JQSTOeg08288q4u3/o7oQ3gXdXB2v2NBZVs+G069eQegmDAzPR/HqgqhGf7FbgAg
oZaIsnXZSwllf6LvmNTA94cyUrbd6y/M9Ljs/MAXlV2EFzEEsEuI2rbDfx6zSsFhpReZacrv0/n8
kDh+bB7ihPIHTGW6wq+wV5SRKEvy2GvlHr4nrXHsMBV05laI/Or4Wm5+SftNz/PJmaZogdMu6rlG
+atQYcRT5iYsgf4xkLI5qeo5O4nUW0+j+gV4mtLNIt/u2PSIPZIkJmoACM0/oFB3j4m9PC+dFQ/4
Id4aVlNLRwwJBYMzfBLlD/E5T/yrgsPdQJEmVyaYgpI9N4DxLEBcdWIerKq7ezZx3cCKOH5gXv25
OWykbgJ1ukNp7KTybVeXXvkSxtajHnYjWnZn+Y2fA2YdN2oHfl70mIYRohDibWHSQuOc1uKvKkP2
RqOEjQLjuH7RO7A3liUPKTkP0l3YRm8e00PL+l7fPYHR1ltM40Qh2tzKBMsQsez+FN9U5yVJ0iot
Xe3FKeKWIkMITh5EJo7LzIB09hEqcRPCkprZXbdcPegFcd1VAlHPOlqG4ONFz9TOzGbBNhcUURoL
VsIJsXj6YlIdTqEhMFperaki6vdTkRuE0tQyiQ/tphSDFXGEp/H/RUEQmh48G2qMaNiXhX0SRwgF
3qTql1f/A+5E4PTE1KnY5/usePMWzKoUhs0UCY2qCQn6mzqMhNxkRDrWQb0Nifs1Di/zkmG5zmLH
YftNax/0NSE+qeBQ+hnzsZyZjOOE4/7TEhX9lipXo+2mpgJBcDNQJKZKxoZzn1QP9dGuKUDiqdQ5
+wXnGqxXW4zVzLAitJ57NtVpbqI2wo7IGNRbfZ//FqIB85Iaqy7FBTJus+o8+3zX/yzzHSkxVUms
gNj3iGXoi51ygZ78XJKLlo7Qu1R2vs5oauAXRsUnZkyXTD6s4aYMexdQvi0fz7adnJ9mw14cOLLZ
9ASMpTOLQcFnWaOvzXfNqKb0BTaM/uEi57KrRMORBUcivBAqBERTH6skqufhxdhHRk7NGw45tlNJ
uCzcytskwes9q7IJVsOlOxp6v3AgHh9f/EQGZ3AOAPsWiM6PQoxjbGEJGN/QumZpNYl4SBn8ndHr
XJI86JTY7620fcbsAW8zHJvL9+/xMKIKnBCXspmGyFbjO6Fhmup9ngXgBYAqI7tVGAhudlQ4BeOE
RoD2GeFtlzOf3hCkO4F9ge41BovmdzaOF8t/vWjMJpfmsWZGfr9/tMqP4BlAe8iakfljl1CzMtVD
VDJfd5xphaH2WiJpFJRjBSHwTN4knMgj3xHTh6YCTIsG9PCUqc9vCiUozi3cpmc66HbgF5DS5jol
YcDyp9jJ3DO6oc3eCbRnzAbSV0CAULqxqUmIwTTvgn29dMhEGLM0I4rm8oJGODoC39eAYYkENg6N
S6yZl72b0WAcfBeXSHpex+IIz+GqHDg+o81GuE9iqJ9wxIziW3ZrRwpYpSKi3Pvig6gMJg057elD
z2xvHym624fLOvGNXd1xnseQ1xhf2Yjxz91gGUL3lf5kqEKpl89psIHa91OdGyWUx0yd3UVKy8S/
OHqfyg0fzQ9LDbHU1BJMg0UDGDEJ4XMMshl6INiWh6uYhzhHOexJcJ701qdpOYZuRObRKtUMQ8ZB
Cfmnfm9z261Eo48utRh5DiJb0XtldnKply3WF0H6ehbMQsWC+SfGyixx7V7GRNXPRnDhzTrPRVZa
GnHoIkfrKCh56rvcyWzZgCWmUHhUEFEjgvW6Vn9IXyC5L67Cp8IwH5U9udGBktI9ybNZSjz3LnN2
5rzrNySBplzaNUCo+qQxF8C2IHdZcS6BmXeuHjB04/CMIw8XNbBmIsqq/cJ9Pz/rc+QhiCCfPybh
nAAAKWmeWOFHxh/1VBXURZTW0b9ZojqYrcHITraaNQdTRt/PFtxnwtldXXTsIv0dGf4UrOaApBCb
jTz3Gvymcbn1TYefw+L/oURlMvoS0uq4QTXHYT6N4fqmgJt2tijfVQZGM/4ikQ/em09NbOvMlW+q
gftlZTn/KCBO4qBFiHe+Wtn7GnZHsC5DPxS+pwcyi3Oa90No3V6op6Tcm0xhEUClGcLiyBNeJKJT
kiP8NqW/nidNF5GUUFxe4pp0IinjqYVRFOIrjyQWdx7xjaawARfdHPEHnK8KtiC/kw9F9lx+Duul
0T95hoK1uNBMLsPj/tRewOe+sXejt2yrF8vgLzUSz+qtGw8UBbBV8pPiaT+AEdYP2oJKpj/fzNlM
+zjBiH3VIhmK85sNrJyu7K3gu83wn5rhaL6XQBK/W/ArqqRYgWwBkzPAt6TdtCkeJ6r4x6i/0wOh
PAW9YnmZioHzjq3hBphe+nggmQBkeVv7iCubHhl8leC+wokIbnLsIVk4y9BMx+9yAPDv9UG+HWJy
5+YaacXtnRkm1mLacEW9p7jN1ftoMeFzFbLg4n2mSlWhuNsW3rn9CSccHvYms7xuYXKXTubnrBZU
j+/CWslF3jk2BaIVKw9m10c6/SaaXWVeeEYeAHU+9vfL0eA0KxBm0Lp7MQI0XIwxp47rm/M9t2Kb
dpdo+vBnsEEhJTQywvmMa+IL8LhCT6I8hDqgDvX+0yK7YhhtiSZX/xIOSC43DY8S8Cu9uQLCctLU
UpXKQVwo/pTlAfx68rNOn+l3DiRuTMx2rYKsCVVDlcQWFJ6Ya0R26xdBhQds6eqYYzQ66dcMLtnF
gaJkA/fZAY7w6Se3jOxUg5jzuwpothHDNIEivqy2FhWoOIYHIZtDQMk+3xPQ2ezP4KCmEi0A8o8c
0FUbNFEWGJCssqblv6r4ifianxzBNonUNAB6CGCKpFBzVZgTDCZWPVBWmUoGOKrmROD7p4z2ZJbv
tzle+XnkKpxNtZqtfwydLyPd6hQx/yBI22YdlOMgYVbColKbsIae6V9ZGCTkOKSkhJpl3u3r1OUN
fbxrOgePDRoevPA49hvnF9MOlwhXNS0jIuzE+wej/ZbbnAWi0MC64/B1g3soic5Cy9PgogBQfqTO
W2C6MQLvRsXQDL/shl355D86Br0SixYUdGI8n+Ih6/ayRhvnakgeAp6bPYN3qtZmMNvarpEiAa3B
9ys22jVZJB9OfFnOe6gKJ9FgsgxfMdcVP6OVSLNRexzy1uiqyqhrBF2xPLWPDIUdIf1WbgW6tOSL
OMIvIlR+aWQKWYg/QqzE5HUiExy3ZA6Ohynjn4aVSlw0omW0LURoNokXLKOniY0EYMxfhZnIgJXC
ifdb2D72upeNzBZlNe2Ura6tvU9Y3Zb4CObio/QpiGdpUyHK643ajsi4+H4A97x3kSdFLoHj5nms
75t2BLFwu69DEk914Ilj9VV5Bl4ZsefKEtrf0OgqHQ/HiOl91jVeJKTsrvY+BbzFzr+NRBBw22fB
A3jKqzHqlLiqmJaLb+WN62N0h1ifYTauCNWc7eMVRLiqHKAjNiVopIldsS9RlIhKt8BiR17EC3pD
8lGZ6Kl4C1nOEzgR2qM6dViE9lOkMa3AUWH8tanDbocFiu8olaA1sXV0QEGsRULkqXCsLo17KUrR
LyKj5ieVM062a2iE0CWYAqezAuJPgGXoYaFUpnU4sTDp+5EKimg0W4t3PCEvlTDdhLPC11FK6GiS
oKygJJuii3jUOK/Cq1x9MCKdYv+Lsguwdak8sEeYbyeLDYvHHAKb10UxlGOxYwKIj03qecvILlTb
PZbgxkTx2OZzrGjX4kqxkX9TE8BWPT4TMvjxf99vAmlwYf9a8BksW6mlD0RQvLIh4rVJFieN95Ik
q9g94NzXW7QBE5QQ8KeNkwFOMayej8BYXpCk8Q8qvSKJZrK5RDctYvebt+hCNU9px5yTs8FwyVpZ
wPjKF7XxoOChzyv+SoRciCq9bsm0C2g8uSTnxrV5WmF5eI8R70l344jgyy0TRD3QhCDaNqEemtrY
ucLPBjIdJZzlcUwvdw6HDfQ2bRQLFj1PoN4xxhh0RwTK652/2Ysgb2rKjAKQKWNBm2SKaPHH5x2p
BAImXT3oU563EYLTyre/ip1V7SGQV4sASwZ+J1B5Z79Duh9bMROY+VsXpDQJR9IyD5gjnO3ubtUK
lPzuaXw3urVxHnHWjSkMeTj9Cy+aGZe/w7w29VX5Tlj4b2IkvjmTDJ4kidey8qHqV8GK0Pq3fvqw
jfmaMSMV/ngVUwQSST2Z+MHc1s5QLaTHyLCqEniSU+jWoixynECrtPonZCswxtxeAw415yFkKHKp
4X6TRZn7an1fAZCkLdNOd+TtVAFaghS+/+Kpl9U8byRe92cO7etXGAUa+LrT2EQ0eHQXZtZyNYOR
8wqaunjfB3OTvajdAO3gCbMa4Ek8IPHkVC4+Zl75ta+a6F8FB/ztJHUhDcyMQ1B0pD1jMM9klseG
4RNdael/Ehjc8JS787dOeLIDzJrxTDDUOw+RGwXXa3FLmEJ2JuVJhUvYwF/0FanYff8tW8LW1PU/
Zco4vREO9OoIu19iVZAhch7F9uoSKcPra6YQqsS5X5YpIZNoKdhmsoH5zrQG9uYC9cpM2+I4Xwz/
uxqQL7NmdzbypSDxa1vtYHB4pCX0oaEDBl9nL/kf9L8BdkY2wZwSwfT07AfsBScAF1hzdEs8zn+7
ORxF+DdNYR2fPBbQqOuDqPBz5DjPHI8hYiXt4pA68ghA0p8O4JI90SMVax7z4ORR0qvJnffd+Nau
kV3eNesm2WVA1KpHG7DqKbumcaty3FBwdo/gTK+j3amtZ+RsyieiHWf+7QziE9qiy+Dzo/S2hBRJ
/Qamr7fRbYte7lax8KwZDa37fwYWvmR0atIry7N8zV1Fx708PesYpqoFMUl5KOudrBk1H9xpQztO
yXqB83hk0L5oytqmwHpi43d7Sopdow79YNjuG58inlvnMeVF6il3h14mmVsD5mE4U/SZR7vtD8hY
fz7Ii3WfpHZtVfeEbPqZ8HX3B1oXisPixpIXqL9EMm3ZC32M0uuaFJDAqjgSvumRBTQYXZ01I+ki
k652yFGkPFNt1SFabIyOlp/s/PSoVVYwknT/KS8/F2IFfhn67x7mR2W4GYZcidwQeKOS/gPArUCu
VyRPEet7k0uIfIA0s2DQ7v7hHfJiSnqV5AL19WWbNtoO6js/wrBaDsa3zINUonZv5iIqD625mlOu
upkBP5j0jXq5PIpbH+PSk5xyNSljoxI5i+uXK2fmxPJGA92O4sbqX4b/VbC80fkilNV3nE8uuxGp
4qRP6dqeE/fKobLp0B7j6a9M8n7Vfi7CRD8a9Qu+qoZJ2N6URWjxwpELKhfB5uB2RvZzxxIdQcty
U/deZGlLDI8/ALbNQrThxRiaPMQQj1WTgJorDs8g1mPOa+9zZbM12dKAJuFbA4JnDu88n+lJZrNV
CtlHxeTPIztwFBacavwwJJw/ztlSQnV42rJoXJXAb2ZgsbYL7pA7mqu7dtZYga5bfgi+2UT6VWuP
AomULyzFzyrxB5BTDG1ojyXPNgKDTXh3yZiAVEYV8pacXSYiqH28yKSscE7yPBKzsc1jmleDKK7u
es443UpUYd/pwpv7oPib1an7CunBW50Zi8F/nKCO789v4F3GSYeR5NvpHKFXAePzhRmPSk0TBrlr
RwdOEX7pCOY6AkJobGJsOFY1KeVn6rvh0Q/M/4iY+VjD7hBv4HKkw8QP1EYDwARL03Dqc5EOZU7w
DbwThKfhmuJ0xv9gOP1iiun0vg3Y/MwvfP2/ryB8iVoL2oMDpIEha66nRZnhczpi1aZLdQ8R928A
WRZEanAblf+LJETm8XIACOrWyl75wr0NHMDzADcK206ytglX3+RnhvTvRhde3+sP+8WV2oJ0LZIN
JfgvEdG3/dbVHB6DL748WyqW1OLOXuA4EVoZoipjQSiqz7ZSbrICcXTdtpJmy0Bnn058JUmb2bDe
v0f8XH50bbT38789f7HArmvUY+xL+YRy7j0WHEb30OQUw4cwYJajmyuKfQijxl/wD8ZG/00b0w4B
yfM3y2BQOFuW1SL+o6nY7qi7/FwMlYwrnGams16lY2Czm9q0En8NXan2hH9KPfMOn7LFlLVnoM0P
8pRUB1lUFHcJl9vIgpt9wHmlrazrbtYAhNF3Txtt6B9uW2aR5rscH8FAmZV0a3z6DbjsDd3HPZ5u
fXqkMkmT58UMAof0zhyzQwqQh8hNlsUAMaaHIPbE/9/ejgP7pFKckkwXAap1six+VxXUGETWF8RQ
CVkRjOYgR0c4egoCjKVXH2k8r13M/WtX7zz/qLYsRd6s6O35jgLg/a3uS+2qmB7Iy6DKVlzObWca
t4EBL8kEAaVzCVLK7EMW561yNXbg3Xo4x/AxL6Z6ypr/8lCADzqndodP+78P+8ZJ7zhIICuWh2qj
FY67qnnLbIbEnokI6QQ9VwgIVyNG2zU4II8AcyOrZTSJ60XrvbPVSJ0I+z3G+ndrqIBo0UIyPAs8
gFE3sG7KHRcKDIkEFV+EM+3rFQaPjbuDBFwCw1cyJiiT0BoiGmlja6XRlAwhMTg6S6l/uu7eLt4L
i1aDUtdQHhfFoq6vSCimj4Qk+19JuqRpjMF2wQW/GcIQY+1rjDFWtSOQ6KW68fQJ9Z9mspeuZRAk
Udcp9VjrokzQkFdv8IZuRqOpdmR5gTpFjDXtgewWF54my4Yt4W3ShFTmjDGv9HyVru/l6lxmpg2t
4uCxq2Rxnx9860D9KABokKGB8hWrYgYqEhoIDC5ysDB8G4cFJDabI+5AaukcxfXiam7qmT6Xsaw5
Mpeo8aQP78lvWdBDSX02WcLJm+inwBgobNF1RjxnYG4uBfC2B5mYPFSgVL/wrOVzqC7DEIJL08Lz
sEWVxJfaITiuYfnJNVAx5IfdgTPo/An5xfR9hV9BX0g8zgNpF9/75dtMA/KeQtO5EaZMHoAZmhlp
D//tEQrs9f7lstfwXr8WheQizShKAZ6XffP5SJogI9aWqhJGVVsZUwvFZXL2M65zQG9i2kmr0+Tl
pR97c91l+TOI+TKTTmFCanuQwhG3Ksgd7bam/GHF3+T6DLSXNKfk5OeGPDy5+pP87tCy7zP52GPA
HahahVn3I6Spdd5ueyg0p5C9vPj3elPUFPGCwCXN3EFjeANzfP6YYbaRSG0zOeCci6wE68hkpHJI
caKg4nhJCiCNl4D7Q383PC211Kaj7eZ1jK2rsRQzvOxTXxKUt93ZLkE7E+3+v4NhAliEdeuiXmAR
rT7td0aSI3HeXtkgYsjnr00DNmfn0yASb0TXA5ej4nPG1KAPD+HAIJTT9pKct8itg7UnNS/SS+vg
SsBaWc6Pcb7xXq0VvRmxzemB4UwEb9Z5jnYEZo8lMqSWilg6upbLxp3JDwrSAgBSH+eXjktkXQeW
jonxhVC+AsrBvi9sNCZ8HKuv3elicThqxm+x6IBm1K1hHjPI7s/f4i2gMvWP8nqyBzGAeltZpWxx
8QL6W1XwEtrNup1s67KF0CTHMxUTmveUbeU3CiGtTDQwxLtLtzovA8aaghRcrgpPBwxgwTD4alfH
1yqkLfVwx+t5HrU2WmGMNy7WZ0SH2hONo7BTloAuerLWajyZ5AESjRYSSFUVgB1m/WYiO6W0i7ld
P57M3XyMeUGB9Bq6GBN8Cy4l4HDsGPJx+8L4+4ye3F4+GRbdK5ReD6YrEGOQDRXavNVfL4Opy+Zl
Qh3DkUqEr90Pcs+hlATPQnIV5fkl8pPbsBZ1d4L6XblYh1WEoKTGevYyC0BpjoG2syl82gmlmdsh
GFVSNDE6wXLP5cU8WVsGL6Iv9nXNhtashujAEacWBggxfj+SP3u4XmWe9dLFHFhgSZQ51JT74TW6
3JF+q5hScHxHSG3Kk/RAVf1A2fl8JZ+vERloS1bHn/u905+xQ1u6B2TjbqjcRpLyEE+DzsETqD3+
n4Ikw2Yk2GSsdlPuraecod9knvC4rvolSrUfZgRnXDotsz2WrVYVcrHbeaXKTHITuZ9Q6EE7f5T5
jzxLdRrnwLviVwA7+z1NAfTIQQkYMxBOl9D1P2HGdWa6zwBOFDe27FjsdSrNvk923E/piAM7HUxa
Wh5zviKUXa5T6Vp7H7nzUZh9gR5hCaEc7Cr9gLdIdJjgmCxTQPzjPGTkuxUA5hCiynMrpgF3SNwS
CxB6/NJEWImwMRT7dt8DdQb+VRq2jsAb9nszyAZWBy1CHxOccsL5FNu4l7OGZSrD+41dpM0GtAib
RWvAH7iUWsy3W7TIOxBqZ3fkwmHlauoNwnzCtDiMvhl0INebRnIAr/d84y+8EwKFezPgJyqlQ1ak
JpFGezDJFCnn+L9R81tNUqB5zyh4m8KxAEAqX/9sMsUA/8IL4Ui42cyDcNyGubfhhyn+Fu3ZlL2A
e718he6rxXOnngwHzTTHxfavIZPfpBP/0WCMtSnA/PPemw+O9fRJqF+qNP2g1F1lZzKUpGf624m2
11oRY/3azbS1qLmZey8nyGDNk8RI1SKQAcRR0c/EvzNLO0H1mT6+uIrDlC7WjIu2yy64HRK0w9YQ
XfjPijnoKo6lzH7F7KwDMAYOEHosroyA5tyfEAoGd0/6yEAuGTur3cOhKuYoeF1CB4SsRTRMxBQi
2tgLsKndyjSqhk/qVthrX3V+YFwvTRVl1sEs//kjjMl9UPMjC41C1PVuzvY/7wQ4NDhtOlwrooSF
lKvtAMre1KVdtkW+T8Qfie7Vwo+KH5Oc6H4K1sNSLe/ti91u421joqmkYBNPTb8euXgRM8cwT+XI
zgFQK0TCBZAdnkTkIfTMJYBBAyS1XNLXGyX3jJUAs61LFURT08Ns35G6XlDiPwCWJtMdyk96FUcW
ML+H+3k4SJ0FHBIhSOsGC7WxmVfoMzcL5CYYy+T1WSqQ2orrHyVfZdvwh9zLhBXwzNJhtcwH78w6
bF6FB+tZybGV+uHl8Cz/FH7TEnwTIn+PWlNsc9wAmljSjUApPl9rXdvPeSnYLt709L52yqFrNNZG
8fxXBNq9SfjXf0r81aIAqGCff9U6PPfRlqgkc/N5FzdJb9LLBKQY16osgrxzfMqnOzTdaM7PHfa+
Z9nzXFH2ar68I9pxqawy1lSrHiHpPPU0ov1vQddMRpsqI3404LhCQFBHnLVELUUZ6LiGV40tQU62
NygASxtO85Uw9+GmNld5+Bb81BNBDl8j1shFDHB/rDVQupG60ANb09gtX3Y+XEFxmlmQGWPV6ja7
HPqfKhNFzNOm3GKyLd8+oo3ywOtr/99g0CXbvm1comuBUQYcwyLRGSVO/rjpMFj5iXq14gIieSBZ
zHhajeH08Nd+504+q/K+DZqRJ5p53ouJh+M2JLt+P+exgl5HC3cyasmUGdWJIILr8Ds6CEoIoymC
NzPfJatbHp3+DBFkcA6UmMV/kirI5ivZ9P3RxUXwjvJdwJMbrSzQZ2OGXXaaAa+O8SjHjDnIQRdO
Mk835uVJOX8PGjqw6jqNp3kcszCvuO6ia7sRFzB3PbiGmpYhvbhkh5hX8FQ4FDd+wRNR+eGgxXS7
eSzBXJxs/33cJiw1mK6Q56I+OhdBEogPyqvkP0VlJo5rRtKtqEaN0WKyfcDnYy//lgdjkZzMAiVM
DBegqpowb0vWs/3f32tRkLonHyamffD/WCrso84VoyCcBjidjZRwjYE+uZFQCoVo9n/mB4cG9uYA
7SdgPpQE8WpVNWCP5OBMXuAp9V+viooh4Nx6gyk/HBSA5b05VNVijywqfXs9kgmOPGalhzIu/Fz3
S805yptXkFWKJ5EUbjMkqVnaPZlvCExcHR1SZbE0xeLFwsk0Jxu2gp+mfyVZhE+7mJ3t6/YDrJaY
ln9eMLINojRPlqdRcPmVi/iC3SAf3dn2sU83QItCCaoMW1qA4adlKTFLXM6driuGkT2SSAvOmuMS
f1kqYpEaBEcjrcQSC7eWezGzs+p4bvHP3DPu3IYnfOSsPfgbsHAS7oVF6YjnfX8TGXrV+NOllcF4
inATAHvJ3eecYJb+p4e7znI+FROX2Wlx0PJpOB+xi+BUBo2jDKZVhJkpiwUM+QKpDNsS9MIOCkg4
xrUiJ3NtIW2x5443ZCfZ/kAu86mVIW9ggU9BUbf1pzD1eG2Htuq4TW+mu92/zAOomeXJWeMq56mf
zN/iQwEBNvB+WG6/eulbtAv8psfy9fwFhX+hjjw3X/yQLhiCS3CsPB5xfX1sQ51LmIXhWG3Sp9w1
KS66U9cBn4FnGNCAqh75wIEe1KDQpfuPpb3X8qc1vG0T4lbW54iRPJoNZZzVQXnqQ0JbrQMbhMq6
Ql05CmvpfmNZrHY+rsni6V0Qc7M2vKOdEkv/GxSn6oGpRnOtruP9F8d9EcS11lQK8yVDhsFGk3Jx
YqY8qqFj5pxtteYbRdFCUUa7jvtNAJa1e5GtD/V7tIgl+U8kr65/iJqIv8iKeEQPTkzG2moctC+P
UWN7wUlJlVe4YJmg8jtnqhlexsekh6D5NIxZUqXhKVgdTShuEynWoeRVTPCeqR7cA93gWnn9doJ+
Gexj/Ymb+CEBqn+Y7DTOd8SpXFyViAJel/MDSXn4uVXNpvZ6yMy5vf4sXFDGB7dfa58ldqzJkihJ
hZYyMXBfu6ASHfUBu1kYLnp12TCpkJ3kX+2pQik6qu36HlRsliKNpk8t828/aW1zbrlQIVci/2v/
Vedb99lMjfjS6+I5B3s+fKXDLqytOGRE6VNPWdHZsZqcr/D6cMyXEc12nOtijK9TCIyoznZZtl7o
TYwli97nUK9nv4bycTFwprhLynaVeHWqYGCAnkWBAzdd/o1xcDBr6eGHzFWqox59t5PQgfbT57x/
JrFUkF1eylMKG4Y9AKKsxtYhqp3kOVimo03GN2FDVIqnDon9MKo4bydKkLNhgwrh0qINotvr9H2b
daoDIB7X5kzSyt9nQbnMISfXfnexlHY77Z2D0MqxaO1+VPZMQYw9ecdEL+vHZCmWjIQTbx0TQIWC
Da9HOXKivtplewJ/FTimr9NcRnvUwjlk0OUlnRiFV8YAoPQ0EqEWoJADML5oz0cQ1BJ+a6ZDxl0I
4/6hz3O+BGB9kmatwktCRDHur+S6trcs7vJdXwaKrmvIObyknnx3Z/tNJVvnuOBRB47dx27bAW4O
TETaElUaLFtRQveBeNhUAwHwbpOTrZ8x/6gDq88Be621EoOc+IyfWkEMtFkGTIsjZ9149s8O0xn0
ig2kZccYZrij6yE5vrEr50PUd8QlR5FN8YZuo1g0ortOYyWQ7IU6LgqCsjszZAh2hLr97ragHvCx
EoXXlkm5KO+pSQR/lEnxF+dLihjS2qytn8+YlWd2A43ZMCpAPk8slZY4jd46v1Vsh/sH55WjhbbJ
jQPpMd0HM0PVLI7+ZlhssjsH1bT2BRvodrG+/flSUEJTg8povq0K0lRRBOTp4Ocvot4XXp1juZYT
7UUj8Z19/ZJ5Rjhz/e6G5oa/T0uEtUGOcAir2jCv6znAy82aN9SfLvruBIdp8oyhvnEMHlZT7pNy
3FtVvlaiBL1OIdMOVrXpa21iqEa9Uo7dwu/p77APgWYTIqsxj7MDcoOHLpzz0QeLLtwso25HZIQ8
93bTqVcDuKQP97HAPQDUiP3RdazWGIX/v/IaZXCf0+/t+H5uwAAiimjOuiel8fdlM/qZccW7Q3L+
SzAJHQ6Qi2lpQZHAlHtL69VyAMLgao1N84aLs4+4C5h07rfVE4peuNMOA16HAMg3b2joPHbV8ztJ
8XH/PD4J2cw4knbZ9h+JzIKFLzxCC18y0Ny/wgVOQNOANMglh64l43o//tN3nDkO2QonJtMfx5mc
xV+6UgDta0VS4MscWjnc6qXr6w49zqrMy8a61CP5hU1bllgLFDwkyf3zDM6bmqZInT1NRc2YlKgX
H1AfHkWVJ/ZKrpG0xozYsm+cSuD9Y0t8U9xIoYRQjjvyks7v9a5X+MuccxtDjvwzmfVZAF8ymHeO
hqtDglwVBBiVJ0623IqtduO0dx0Ad1ujwtfQUINHvw7bhfJSDTHKZqMU/MjYu86S7smy4juUsPkg
hmkbu3cYJETtU7emdZU6yvplRWwzAl3zL41sxJVXNFDwV4SUV8lY5PXlMtdOwjn5eHvXn9Cs0txc
WqepF+BqnnTkyQp3uLTDXjKaIm1W9fRgbfLs2nM0bzU89oGiOm6EY6CYiROwxzlFyMhKDxBuBWX4
akW9qYLJSXp4rD8e0aAHcoKH3qW9NXRu5f0IOh0XT6n7y1jmCuVi/0Sh3TW1lfbcFEW11eYZUZ+a
SB/ZhJsgPFQMF0d/X2wL7HvZl4W3Ny/Tkw4Y450yy9OeLP1x6DogKYn6zGoDFNjTHEqWp53XmURf
HOGria2CZqtBzcAfAYtsu0Xcj3bNwD3s9KZm3OQ8l0EaaaqHmv6XwXV62FrIy2j1RVtpJgb71RXG
QcJ8nZVXfZff6v0pbglOptUFI8RpVpHgUhJdIxw/zc9N5hZQh7UwE4kVVJ97dclsdS1N1nsPfCAQ
jTbMNbKDRImX5oAhoCsma0vdpssl0usmSNuytyM+ymbocyx3zVoGjVTyIXbVp+F3lkx8bLg2jyvK
pgJ8IXlqT4ifo+Vb+i1C3+A6mbBp1nGP2BZAyxP6Pr8KIKEr1HU3kTMpd+Hpn2g+JGR1YEWDFKk1
uVepbZ/GClw6IocMZ/anFhszUQMBVEp9azcY+dtYG7lZknEZQiLKNldlEo6yI7BEUh+pZ6mZ6kao
JzxhUCXtoGggf+yn3BTav/4ox2qrVOZFaDuDgrEeUtRuj+QgejmyKc/nvgfMx0N81MJIC1Jse6lM
ODJGzyMHyJ2YWvX01VtJGbGrQhjlGtQrSrkHaHsNPQHFB7i6J+D1VGyRRxFnROxz6t4qbuZWpS/F
7n14Ijuct5uQEL2i7FSxYoc8pykFyHQCkGHSyXCF/0Qnp3Ftn/t31MTu5YK1zjHqIREZWME8ZaH6
6QyLqwlfeQVnxFy21Z7YZ1fFCbWQ61eGfwXzzdHdo3aDAc3ttnaf8BEihviQEuZxijYGFmIGuU4A
764JUoj81KUt1TYKwuKF6XCIPd4Q6ZriWAZ36Hs0KsXrJJiTPAiDtOLB+A0ftAV0i5shOl/yOLfL
IBWjOR1VqxVEiVIOBpoW5wCpSHwEzOeXfSjzJwu4qo/IEmn/h013+IL+6WUtUDtEhXfKT12q7tRV
3mphHTCjU3vzz2KrF4uRgL/0pW7367EdlFE8btmplvV5uyw1AET3WJppJDwsikJd+NcsYIRzLbux
gjbXUcWEJflQ6gnuDrbzwKfvJpvA6Pbw+ts8c68ykap8p7GTKir4vtFyZlgnML5AZKK5eozEaemZ
MfAJ2CoHI54r+BMZCZBZ0LCDONAMoRUjnt4Yosv58LJX+dWFEssZHxcPlbAJKxSGwPDwszTOC6wB
gOJ6Wfqh2JDnZlIlPN9Hb8hF7w6pDYVs317AXSKts+85qBwNnjvIzybMBo7ChP6CeHXt85J7NEng
xXzwp3aHNLIHPbgdSHWyB/n3RhuHRbbsmofsckixWC/Fd2DVNjSRZI9R4prTINpRHDuOrDInZz9t
PUyF2rOXIeBtPLzR+rA0/bp57J1o1xIgI+jDLGNDNi/rpU96cm5fkzLeRDA2OughrPWv4b+NkhL8
5J96hXTZ5JQQnn00ras6suojI3OiaKyAdP2+MVOPK3IwWE5IkIVGIxp5bSOwKiF/SRbYDH/hNvmg
215CKpNFMrRzbKDSPs2boIxiDtMyCvbVlLOlE4p7jpGJ9KTQrNabmiJkjM9v3GvfGovfAdwwpR/C
CoNGLXtD75cN5oA8S7n3zfmnKmu973IHCxgOagRsyk5JRzCtz8KPcBLdQCzGrbnR/cUi565mMCtv
8KeauWuK1OgBycK701stDRg0CvA+aBQFuwCbVknONwpRjFJ9PFcKBS6l9bedf+1EmZFtboxEIvDu
LmgrOR0JrMsp+TgANsJiZgTovYNC2ksxBGieoSc9v1OmdYIMt0ydRXTkb1WhNrFmI2Z3GVw4bS77
XTg1oEo60KtZ7tEfohSXxnm8InROy1yuFRRpF5SsyYhRB6UqOwW9Jfm4WATowNw8VL51wLsjU3B4
g+QXsVEq+JJMDHXtQcUuCt/U/uF/vG/ZYWGbEMg5AWdOyub6+Xsp5m1jPCPlqBeZcLFxhnbCKWVj
5KrrxkBQMeaqIXhPQbFH+FnQqYiNpB1QDDhXN3FYO6gBEQpaWtM+HcnYV7OOGCFdPAdvr3TERvSg
4tFbiIFMrxVtsVxHvjhxqAxL0jDXWmfhrtTKBEqw+wk+3QYhr8tz1nOZtb+HJK5ubTXXZZCnQqyq
bkIEb3O49KvxGKWuDnIlWBIX0y3HIxRh3aDgRwzt4GsA3kzYfcyn8RNn4RDNnBkbIhdz2Z1s2/om
GFfSwc4rJGpOdDNDAb93knOuyy4K2ZHEZyKVgw0dwpaavnWokCEow/28uInB/YkCEmIm4UfJwbMF
patLldlluW6PUp/5oyFIYg0pARu+BdEwi0y10a3V1GsORCF6gkZAztqCUiGFT+avvN+xLX6C9p4H
nRuz+k0mMaL5dzf6tHdFUKQ6gdikJbfS6bsbgsLE4KMltqGMxjg8OOX/NAsdp8otIM7kcUZz36p/
NL1a9p1HS8ki80gJ8dXcU4+kFcSpOdgsNOLznqP4n3Flr5uKNi/qvceLb0JLNPOqXjXwhT2BUUns
ITEQSHn0QFYePrawJSmjNOro+FqEQ+aL9aVvyqvSniaNyTUburC3aVVFD7qiQAHfgQqVM/nAQn2U
Wq+Wzs9SwMdvJu4c36Zp2TWWFA1DFvtOYInMq7P2BE/XvYKgR9YqaDANT3KY+hHQYZvWZS4ZELNE
3ctwe6nhJCl6OgJQVfDhdE1FQb0Xf5QK2w9jhDFWFN48G0sFdmXfsqIzY1ktk8T7PmJ5S1zHGUUh
TEkPU8yOok+ivb0mKAAvcX6Quff7VUSuCBL7TWxQjnev9i4v2Mt1+AwoyyqHV+cahbCL4zBO4a0E
/8DEiTsrNb6XqvZ7lEAe4jd1z2yMPpYK5wvAVf+4zKFp/VBgnrBZW+WkJ+cXMYq9CYfYkcfPQusZ
8iSHqPuOwHgN3jpRIN81IPh7QMOFecBEExKtAuIDnBIlSi74EAIli9HtoemTbmJDgHctBxUAwG51
kJWpjUoUyztv2kPWQ2aIOo7EIxEF7B2bc1GQ/UmitfhpwvI+kNrUHkUXcuGbMHuSRmX0jlIK2HYq
KQqIkjWBDgnn/HelrzQvadsU+MrFOoAu63/VHs6KhubiXUDI9cvfZkpa0593IGKwArJ6JNoC5b3w
2Xo8QXdQGya9deJ2JjROmqjIZEuPQ3avUmrwYITezpYqZy3CQqOAW7Rw3sar+tfUO9RqzkeirajY
0EDksTvz4bpzWL5m9g3ryD8sLXKvxdxmyrXSJWaBmDA2CDJbxUlj9npJZ2t8TiISmKH/jSQT1yNZ
+Y11tyfMZ3F0f1YYPiD3H/bvFeMx/2q0xyAVIcROi2sS3R607KOpgJ83eT+qzzLY1hxnJpu5imOy
uLZckIgKeHiSGHxenpEl6IFMY7aRUVd1qjzcTcRf1UVbsQarm968UHKqX4FoW/88RZAVdZsEJFt4
IVGsGvMRP22x1o+FhUj5NeeL1ZBFhr3IUa8MoV73oZIqFKv9iXEtnYk5APQOajUD0DzjC4lA60n2
7fHKkGkxgvd4z7wkTEmnxS8bt/8erHsSKd3nRrbaa+TIMvqu3FCij6maruPYkYrZ8W/xOdT/QrUI
2jXg08akpoaqcgxsK+mwjcSQz7QU4hQvgf5+nhtrGECUS2TiLpmllLv/0w2GxeLjsUdl1QaZZx5v
ryW+d0eE/Bzh1i9DUE8/zrCfSWvaZ0Z0qeuhGCTPJQac+48J9bGRJq3rrovyBnbVnh2rbhTg0T86
c5PUlJfVSex9iox+W6lKZWd8S2/xbho57W1t1YOI7fM8FjhIXvEYHtPMsNeQycO0KEAxDnP/KLH7
TQ90cn9K4cDcRfiBNfJYHlQJ/+su2uPuB7hZc54AOoCiDU4eQJ34IbwxU6IdOEH2bui75ink5XLy
vdGtrkpKfKiWVliEJ1vZ7dX4uKZ6Tnlktokz+Tkx3iC3TrVttuUGaZ0A2noAdeYxCvDlBx6Xyc7P
6dzHUSSmR+9l4kNDvKhVWNXios8jywjq9z5xA3+KJ6zSvZC437rVpPZ8U1x26P7RXuxKWy6BU+he
ac1UEPvgLvy2h8Ak5b0yaC7OjEH184QzVLwbe0ndcrDTHgwFQd8CJZsmxkapHGMC1wbyqd4CjenE
FdmTLVZKcS/7thz4gXHO2mmUd84HpG4DB9tJHoiwuPqr8EtN7OI2kYz5Gors4J19rnOsLC1sW0MV
viV7rt3JY4hI0Kw6QVfbhMhf1FGkFIVAXUJUHQCljgRPC5mGr8w8ZoO2G2QgD/wMQ6LdbyvTZJxh
WCjgEJeYlgtASfRRmTWSTI83t4UarnHKImEkd2XmGa20jLTB/zzP0MctLDbYKdZ0YApkr1t3N58+
FeV+HsDapDRPeACqYDMGQl4sjzUY27STIDdPT2ymgGim3XCIXiyhxW6m6FGQ0XTRGiWYqcqeCTPK
VfEqD/Vy5Nh+CqX7DOMhBc0j3+2LO+aKjy537BV3kP+rPiIi6WNIBF19VPC/VPqYn0QQ4vsF7+h/
7UtuomkrJutv3zetAKSQB9FoCGvZOW+WXJGtM+dW9b6zTJOuFPsdRzogFJBysG1rY9MtkYrDk4Mz
bbYkolR7tHvSuWmhZ0nFUGMnJpOnOb4E8ygaMRIwXqC+g17TRjE1Yl2T+McSrZOgfdivEJTrITla
1h+X3g+DPu5aVYhr0AYUCWaC2rRLy+vAxoL6o/R6llwCNKN4aN23VT/iNRDSMt41kDJfRJtzZjuk
jYm4+BfnI5uS34JAcr6zm57Yfyq7iZHMmYwrkQKkoC0ohdTSRnR4mabIZUz6Os61gHhq1HtIxqPY
ZhRMUX4Hi71IpbLhnE9mOn49fGEuQG0O+jWo6r1gh08isiX+wedEhZJek4JQTqQxjcECuHxduuBk
fGnYzxJXhhrSiq3mA9AKuGzK+Orr6l06kqYTKiQTOJnRn1bwqoPRMEDFCdItryjfONzCWnsCpgrR
RNi00gapUPxOY4AHt7gKk6qUX5x1uYux+AigMmE40O1xjKGNy6Z/TLt0hXrwo6Alj/wXjCysY8c8
tmijY2p5PLnHUfWL3pFYg+byviBhhOTVfxRKzO8FzGOFKzlWLMabFJv2egM3lHswHli689NAjjw7
4CKde7sZKfEXj/ozZXszUyYLeXKwqL7ziIow2GcdxxRrKYcOQS19t+n8AlXojgWJLghOPvO3hVmb
u33Cz2iuXaAc3E88KljQPle57Vp7fdGVuida92qzmVmgUnCiHpvmUvLmB3ojMNLFWdtb+Hkd6kC/
N08BqL1fNy+sII6csUw+/RXxOMODk2RaUGJxZ58S1Eol/jqDH/vWygb8yiqORWSvlE9P++lxLJyD
I/114gtZdyU3SNdW0Vr60Uuf9fSAPvxJnkwgyCKmJXgrg6qn6Ay/KYPC5ntUx1XsXREgan/bMPWe
+2iL8XuQNMEwsUFvfnAUfNYCQK71o/LTaW4XCv3vA6I7WrWjfuIx2QL9BRueAvPsq8SoNo28bhCM
dbOFLZBGPzb6F7QgAH9LNbR2JtECXfIwycxWT6odINPzsg72lEvaRucz65a+am4udNQ+k2IeTzpQ
nD5wQ8QeH1NqZnU2deIQynYcx85UQePsS9nD7lyQJLcaty/yS8LM8+12OZQ7WlfNCix3W3GE9Nz1
W5/HLCcq3hMadrpy0e6Kn6cTnzZxdum2Ji7UHRG/zR8Xj3dn9gfSGi0kEms06lydGQKMkhxjleXR
3vOs9EPnzF7at9WSwuJbxDEgR1fb1yFkaP27Isca08TRFvYKzGEuyFoPPqML1hu88vG5XNirJ55q
1G2wDKNdIVv/H+kqNOnBW/CQNaV+oFrlYTtJ1N5oaEF9DbM5tqIvM48o8+bT3K5/ov+wbWP9pZI3
h7AWs7wggiwvLox525HDd7uQ9pdwFfjUttbuo8VFlmbDCBIXmk932DXT6fZh4tubYMlXuMlXosyF
otMQHgkUyNEVqYxnIw8MSXVLftKLBYCoL01miNJopX6HESFrIQy9o+yZWrYKcKgMbHKsKMuGpBlY
L6xp7rgsFJ9yIBL8zDRwntYDEAcnbXPrkSrR/MZ/q9fg4Ewq4nZo4CRaX1yQmlMlA1AFJq/5nGtT
GN0pismHNL5fksxhRHQeDAWUsS2i9CQA7zJbA5wqonNXb6iJ7565z4fZKJMuibDZFvCbtCmw9LXA
CetzraY0lIQ0aAkm6jt86gAcwYIGa98hfLwnQn3TYmswqP+raDITEeFyQeT3tHFirrcRrPq4MxFS
mb6oRK+cH9Abal8cz4K2NaldEUR9z3CA/1jzt4NPljSzQPPyWpaQwngbRI80xoAgxz6AO6yQA6lr
i2TJUpL3zILb7yYnp7YSe14GCl/ibW+If+lqKu92/nfmswUzGj+ZqtqIy+F7ffipeQP2DFREtCJw
mQChbVAU+ENLkuPxBBolgnSC9bkgl/F96EXfMC35OO0RhtkecAbcs00daEKb4J2S4V/GsbVKEWuF
6lvBXhe92w4IO3qcwRrnDJ0TtHepRap4Yoq0J6JaUMdz/1SEn6yAuRSe5Ng3Vk4Y1F77mldyOWNh
cQ+fO9c2soT+dJpgwSvHjR7jQgeEm9ibaGFfXeAKOUu2UKVlKXhvcC9v0NOMh2yZ2Xcquv6T5bjx
kkrZJMCEv6nSbmfB0V+oA1dukM1PHnUNrdS+Tjhdu6zkZ+X/M06QiN0+o9cVU6g2GB3zI2yzHzCi
D4huKFjjGTt90r8gL1QiX8U0ycTgIykIKgO/pQ3T5nHom89QgjLl2OUdSVWlc25VcW25fIVm9Pb8
W1V03juWUvBtFalxFdah707CpJRoBQJeCv2eLtHh+VCi7AQAA1RAgOxrs5YzG5t75NqgQKJ5HJXe
SxNMznKEyo2LdHWDrz6nZ6fXVHXwVJdaTzWAr9EGjev2GkSPilen6DaciGTxaDi7wKeWFpdiVAdp
ARSlWpmSiAL86SLO9zsNeskcCYveq9K2fEeOz+o0BQ1hacRP4TdfJaV5TORYfPSbbDb6gg/XpxqS
XMgUSX2AGPIw+SA9zA+2HjRpBPNIJHE8tDDFe9kJk49YJFyvd9AcbkdjtKdQNfwTt06S8AuzePcM
TrQy2YWfakoAJvuMWaijEfBtC37is4/auzGTddpmpzBY/79yRTOScILJo5wKtRkklOSBDDXSCIQK
GwYpbAnH4GvYI9XtDf8Vyw7SmgdrOaqV279hnfBmby9nAN/yjVU+XOklL+1l3jNAeKuqJ2vWmwF5
DgLeN+UJ7cWD65iFJ97/66hp3c4Ji8F6+55bR7DQK8pIcktJvpfrReYdoosUYTYqKkyi18EQqNMl
f9ivtvMO3cH6MF0hqtddg4PnP2ooX65+MMAX9EhxWUMGzUzBkJrnLQ4p1BBsVVj2R4+OAfQ+g/Sc
BQpC4DdCfnTq7ND908GJlHOxfKF5NIPKUkFshsgbyPuojSqS93+iW10bjNOq1bpLY+qr7r1RujhK
Pj26FyviN7OdgBPx2QkvUh68kruaCHWGbuwZZ2bskUa0eVLaBux3M37qIj4NYAgjmFzKS5qCceaE
d5mWLCNoXTqzP1MB4EYhr0L08oeDwVj0r7dRqCuvPoTlHgpb2Ddkf6JIgBuo5bzrNVvfKKSBxkJf
phV8EbWrioeyYB7qbTrvMbThSq/zVc1DZ0Pbw79xGzjd5TdIYtSUkWSTJ3nBsHDWQdUAzpeO+fuF
1TFeglT71CQulVVrqgl+7dd2nBme8GTuvHUiVL4g1mx8WtvqC/d65a0EsLVv8+AFykhYWDZ4W9YQ
cS0wpRXBO5HwKofEHJx1aH/1e1T2bWLGa+MVAbIPYri5So9jebLP+BQVdR2lpkC2Wk7i6MyudlGb
hy6IDCLf67PxSaZfnCOje5dMq14eZITO2vmi6vRAjuI1erQiFdl0kco2e0nYeD7AupoaN/iy+O19
rEvLO/0hwyLDDxtDGVRleBjukJ0GbiPsBrHCzDxUM+J+NRQcDYTZYv4T4yYwEcRvfF3g3oF0qKRI
6dPxPYja5nBNuf1UNujW/sHG7skSSrg5LTF6EBRm0ZEuQazcpJnNJykfu2wGZwcE0nEZn/Ve47Cu
QuSlppfEJDCYX0ZawOeYXjFl4MEjXEkNEDChZynMa2xP5cJ31NjqLS8PQcZYaO+U66VG6pVHwlWP
UIMmWAboeAlZD8GPD/cK0nP68KrzId3uKM+icnBoVSt2mGu0OlvAzD4ZvqEswF9Eb3LACoPozL5b
esUh0B9viq2xhX2VwzaeWzRQGRJwCiqzlnXJjfDJgaVRGgpmFOjbAeOefZVgSl7kcTRoSBjdm1kz
5S9goYRC0s79W2+sxCeR2qbyFACOsssb9UKXfDLny7QnuQdnoxGEBc9IU/WxgNnaVadvfdtlFZsa
WgxW0z4VErp+3Ue6r+xFATa9QPd96PcXRzsj8xNlTRLWTN3Ak5ESxFQZaW78AcJjXHTiACv9hXGZ
S2EmIZuS1g8ggrT5Z2R4fxdW43jeA7OYqCZ9NoT5Tv8W43N6FlEis4znBNmz6NuluqNqB8Bp8632
R+lmneJmpz6ZQaAH4TzZkUzjNYAg+AGprnpPnvai2jTCSRJAesIYfyhWwYgvwp+ni4bOKTmmRq0R
tXZjB5nCoHOrB05uZDKQsdyBHhfiJsl4uVAL6nvGsYIcdo97cCSTdG5y9yX36AtHCRSz5bZ1IL3X
K47t77QBLybJ+4BDm2TPcyqdc4ZTff/ktBDnkA7C0TeL8J177NzC7P8XZgvmqN8x/1Cmf1IUkbRn
N4Ks6yv79Qn7vLQLPDoHAtCukrjSWts1+7E8irgW8C+CmtHwWXvH+l5fzY1khjHbdTAOnpEStn+Y
uEq0Ccq0zusnuFi5evaEvunQekyehPsigxNUU2K3X5vFz6axuUjH249YEiKs2GFyVkDlHLyfCYwN
CSHNQUmz1BgnwuEQEARR4ZsoS6FlPNMnR7pdZehbkkITAH7heC9DhYP3BbGpU0E+VQXvFmwf+T5B
LiLG2W/O9RvY7PTOV6EASsia3jE3m+tEbRgnBdh2aR9IviLojf2yotfgOcmTQxRc6JDtewvJc0Lw
4OuhZ294heSyfKrqw16+Ol62fdYMM073z6roPLNr5VoMVievAI12Qf7k9qbUpP2D9N9sgBvbPZ2S
VkR+ZWH+v+MqXxPzrTmUcKgrBj55ZV3zM/fQ35oWBDklw4/7F6/zhkj/UM8R1GIn6mhCQa8BTqrI
Tt9aP9IBdhEC3BK8w1R4dzmf2KuAkmcqnVhr1Gquceuc7w1FpmisJhsmMEWHzmusRmsZ91yjFHN8
OFXwIwQDAksb+2vaaX1PfrdllVYRXVMPRw+fp1ltDgFoEUlb+gcF0zEPgTYo2rFpsaUDX1aQyG5f
BcGCBhE+XAfbjFYrK7Wr5ShlDA/FBSrSALCc0i2cPvximG/d0SXsAbVNNiMbn9Rr6QV8fGFLCOTs
lJomjxJ+is+GXjasUxOmMsg2YT1Hy60ErnqMAKNyfsC4VphNZ27cdbSI9K8oacxV3UbcejxYG12l
YVt3VhiMaZwToF2E0vZjAZVQlSEYojrZd4dPZLzA6pAQCAr1PRZMFe3VRxnJlobgj+f+nZLAw3EF
Bd3M1r+/wkeh1gUAcqSaIN5cf/p46Hmc3xkvmu18CZMpw+us/HIedO7Y1n6CLzh6MMm7MOxK/SMr
qJv+yJviJm0hcz6vzfU9klqTb9fYYvM7cpf1s5shpMohQK5vqKjJUmx0S5kQnpBqIjmR0f1NLdZ9
srmiU4dhT47qb25z2Yy4P5qudHE3NKKLk/rbJvUX+8Io1VSy7rlD+Vt/d7MvYn4Ac5v3I89KAb3O
3zqCPs14c5ERePEPRh9IcLvHGRybp0RnLc30SbYQWM46mpVfXZ7Z3qsL7Y1BtCJfhsBuEUucSYEq
/2kgcwozkDG/3/Pnsl3dk0TwdYvkoADeIKPbNa4xXUXW1tKrtafvJaRKLVEwVPuIbwo05vgj47oZ
Q4u42zDp97a16wc6BLevlineLlEGyzXeQeS9nm2GFw3qc82edRWiU6is8iVREx3DySm1jYUxnXaU
MF/aHGAHLmr5/NMIn+DqyblN6VpPKzz9ECPIaE2oH8MzHeuSY7Riuvg+eybxAJdbJrZhN1n19JuY
t6Czlq/DtS+Hxb1KRG3QZxdXm0taRyqb58g1JkLPPuyrU1Lz2CEA7xFZ0rBwI6n6CmuebbwF1YdF
pg/GyF5fJgA4DYSYTQ7FRBvBlcRPhBgMHH6veTslQKd5E3BjXeH4LgD+SUBsMzVqtbnbAX2ZFR5U
nvdybXaMuKZ34mj1WxK83XRCfEw6z7iLnlZPKrWUda1XUkzP5ITyTB46OXhvzgmMkchsOZWcs9fu
jofiZifU1XCCs/t3679NFo2BlpR0MPBcZJJoE0b1hg7BopBZjII97g8d1CzHdb5IJ/NUT1P/anEs
GNbe5z1yLbBbfBTy67J0WDQND2YIi2RsJbpBVOF2NFenLGOELSVL2sIaGbypSdWCF6iGXZD0h+18
5mAsxkXjjJT/DOesRmIPZoQ0bP9hJSAu6Bk2AF70Ufrt9L82t5HS//Vl+N/gVbR4diaaHGX2L9ad
wUPbwtJprBFCGPb/pSQ6A3XwMU630xlHfQdDrlhvmeGdgiXeW6a+Hbpi0pySwcTqbOelhMVUo0Xk
6DA4vDSqTVO4zNz1YGGx2+30ENXCs4ug7ovHAaqg0P/w7lJOSFC9Yf7R66852NNC5QKb7pE9sKkb
0X+bAeeyuGuopXbcv8w0gRtOfuXTTeIN7NeRn+vfBg86+lWOU7bEtFZXTRBV2NTfxmAi97PSZo7e
7bLMi7uHny884BzMji59SXaYx96SOKktHUoiSSrmKedNB1NF5h8rozp3SWkzjILOeMYeg2DkHYqC
jvxGaBX/kFAHGl6LcyJGDSiD5ZB297UR9uC7dgGUIhK5d5WIeuCtHl+O+Rh8XqojpkPi9y2ckqNN
rETTIz+WSXth50PUTposynEOUI3ZTKwYLrkvJoCohrLXKTWn8errd0BTNO0BjSKfFcTmot4Sb8Rz
+dZil18GOSQgNP2Ruwq9pR2HfeqiD+kiNFu0Avk0OTEC1jbMHmgOPAJuFgc08qEGbLIYdkyTa7cZ
9oXspyY9VubJVnNViT3g4ZM515cQK6axFpKauQSeF9fMxGiACAvT7vpoh8+aLp8fjrNc2vU6d4dk
wnHU7+qiMjHhrb1B6Rk98hERfTKzPPWU6Y8lsSCE7IRG8y3bft2OsQCphTguiKCn2ZGXWFk7/QdT
jBzXEiEoNeCv2zMRxH0Fki8nWn+C7UVhxqKUEfmbZ54elaE9IvVeGijj+L82wgvoJrWFMWKU4wTv
UZ2FnHt01lhY6ulAWj2eV4kbQaUL74eS7E+GwL/qXaeyC0hDsrzDzXcryrr6D/02glQb4kMilqGb
GLrfjJ54sj6UWGNk6jpaJc9xIUFHvWMO3h3p0htPjeaIilEtP7nNtloyycrmNV8UG/q/WOdxVBGR
OYMkCtOdGKYAy0uxb2A8GQZ9K0oc4q/o+6hTAiI9kz3VKhv00JzQ8qs2Eo3l3v79MMquTYdvGjJC
vHJlMxPjKkcA9X8h+iW9REtbiI2bnBrgPs1P2vDvXK2iNNA/sEkdUCJk4VMvgqBwnhOKn+VsvxEe
wT9q8i1CM3s/XMCg2E7jKGgF9ckz7XRMEXnt2kqW4NuLzMqoju0lk6aNyUCiP0/fAdnoBzR+hPg/
T3h5wtjfO/MMj0ji6DM/odEBePO+rLXDdyGASXu7jDrE7ynjiXCp9DTNhjAreap9Ztb5OhLQvH/c
9O9w5gJcc1iU/H3dhhCZUtVFfpcqhGsIewMjnIN8GODUt8doGCNdXfenV5dMuwAxEhHXEkt4M1U6
+jczBEluIebTC0GV9WjFUiggSn6Q4CZnfCgTnhMCHs0Z/2e4kOHCTW8vMtPaCg+JEEb2UpihxVYt
7xZJglr7E/AWjppUMUWEWip3shZ2VBw0N39i53WEiyVyRNy41b2u09KqsXB/My9J7iihfYoJGvd8
I4g76Tn22cXisstIBl2fODBjj0D3u/xiM0BlEQNUUJPdqgwve+smteH5BTeQWJMWZ7VzFM+ejiAR
2s3c48VUiIReE4o7ZBI7ZDspEDwP5A1yxDkW4Lv3pkiS8ln8IpVgcSzgNwkejwEWxUkoSyIJ46dx
ORvDZ71Ox1dAFbvga+X4A/W45AI3tCWUmtI0PBbJHsaRD0yEVIqeJczEv5VR5GScSYlICSvqCwQ1
5e5ffEKCCkibEjEwhcRbvAsz0MjxosNFjMLSqJDItnws0p4ZQxbxkqWaB5fUmNS0XhHH2fda+JGB
YWCtS4hstDOHTZz1m+BY3cggUafqkCStfPnJwWQiEIfRVykE6+oGY8lNwIkPSy7S6bjX80RuO4gc
BNBJOsMOq+8m16CF9oLgux26Tw7i0NKWEby6d/S+zv8gO8YWXvDYCHpDTk1wTID/WI2SbEYO5WiP
ijz2A9m3WOtjluNyWJoisAGn/mP5T12TpLK/pZa21cndMrC8rhoVGW1Y3jkKsmmliSv/SFvg8YBt
wZFcH7GhDp8qTz86BV6YexF8a2YeuNTrUrTg9tdn7a8SVtFz4y+54A3BXhnDrnopPnTWMTZZBbpW
6Hl8YT0lkQvQCnaCQijCnwBUxuZV3MR8T/+QPmwBSvqg+OxHAvUvmqWClIPRLx1XLdRjmTQRWdpO
67WcP1QcN7XhgkVSYWB4CkSbuMf86kH4LWKN/tRC+T3eqhmG1Vo2JH4PFPC2Z0NtJOxH8vMpo2VI
EJl4zwkyYok7C3AtMxjy5UO4bjPBADp/70CjsVmyIAw/WlZE4EsUri8+UXGWwT/IczOLu9M0qbLq
p0R3aiC8lRXcSIrn4uIpzU/4UDxU1dksUkgjAkaKNSxySs4Pyu7pjKqz5eNW2DATWcYtnoQHz5k1
ZnUyr5ONTZ5EtcjOY+c2nPVFTTk6zNH2jq4K0TsAjIvpdBpIFyTJNzXURjIcHgNpask8av2sVz0i
lOgPiC31TfTJZEUp+Q86haENPqo4VRM1+HJ5CXPpkd0BZM74w3V1DeJins70aG5uqUc34FbFTFpb
RofRnpsJDZLIKLttn7hspbE+33jAs3z82LUEyx573Ah4QuNHqlXHUHAmECrhaM1D4aCd0f1c++hs
218oS+v7DKEkIuegi9v1Vv3N0aPZk4hu/gNcc+CdToFvH3U6BAkZluEJ5jZxuhkRVsIUa5/5eOJ0
wI3nsfnH0VuodZJFwfAHoHfgtv8rJPTR7mddvuNeMrKUKMm18HdRT5Wxe9wMAl+GkFngzNWftsZS
dPQuwBYHdopMqHORqQ//HKevscPVnqweQc8OTclPb+xPEGi+zaRWM5lppYrujEFrzlL4LkNNdgCD
5ntgPBf6+hflgvn67KHphg5fQKeUNcFHDoQfpvAsvl1XzMURz+NXFIqhmH86hDXKtFTMcM0X7htd
HEfripKDmGRwXVDe5DFde0T1I5iMXzschjraXM7ba+WBkZJt4pwfneGKTS0qzh5cPmSnSesGBPRx
Y7qsYAR6mFjbDjnkSRq/2i7UIfc5ISBJQN5UNZPVj4x09UCqT6kfJNZGF57QFj6rZDNRCg4eH6fx
5oJKYRgRjGU10OQZoONBDU94OaDRgSWR66d26sznerelTbtHJEaFEKabRw5oFpbGyBt+AvGf/ee9
KifxvormyBh9AlVoYCCj4ZZOH2FoKpR5YtB15kSjzKPV3Fq3fD/uw3xkge6zB1zieuTlrfDK1k8h
5Xa9FhfBIYfVFLzSHJgnABkIHHrN1/Wpz5RGTbSUl3rvL/qmBf4eI9mbMR1JOVV6iVjuPpjOBG+5
iFjsaeELr77glVJ8LtYt2uYq8XlJ3TyfmbYAGD413uSdgBsMuWn7h/EnBMzCyz1UkR62y/LQKf57
zQNFfaO65wOlKbKFL+4ccPBxyiSZmJkam9QWCsyxDunBWxDeYk7bjVNkzIbckDRL7OTLHkuEgFt1
GWMReqULHhlHOxkSGxPmYo99BIQ/gXU/E8FrEAIBmJeZcGGMIe82urFI03EolJyzdTQxM9ED07PT
AnLw0VfVIo4QrfHjjWps2sY7xKY0eqiAPSQPSapI53UJLDFsjE4mVcwrjpyO5Mi6izUpsvgQMZUO
kXivRqIPMZ3c2/4+t+UDXo7WP2byOOad4Jibe6agiJTMDR/NnmE2MIoWkGoVZnI9edd9sN0U5F68
qo97xV0O4yN4CNGYdzObh0dQi05IppFIeWh4ZsahnQf4CIYeiyFN8DMTsj/1OCggp8TQKjNyzEP9
GPqQs0oSGwFlVXvRk3Ah2fjzdKW3AjvPVIz3df9/J74EXcmCxe56Kcyevy/3LTxuOigiLGe/MRY+
YUU1SoDdg9A1aTKOS/Oqj302PMqHvyE4C9/qFjBn3Y+aCB31k4SMnuzIuRPYQTUHkw60/dLUp8vB
da/4WOgBs5CftlMmqUQRcW7U2X6T2f+iyvwQ+q1SEmeCHXiQx3CyWAXUsEBiW8ysYpi/aPqzUEgq
9GQFv4bQukhTIeZ2yqMiEIPT6vCR13wAbEke5yP44z1v+hN3OBFJuUA6zNIuoU1dkzdEfSsu9HU7
St6TIFKyHGtl1kUfdfJaV5RTnPsRCpYU2v4TvQKhw6uoNBudZc3OmBFGXi5Ism228bNuEhO/SEjF
+Byk1b5K6vE5vQQjmnDlFwI+4Cr0XpAP3R3kv9IsGPwRsDXALeIUcs4GebrS35tjXrY5uA7SB6np
sePQGbSiiE89057qlPWkZNmTjxLZWS6MRfdjpwK16AJRj0KmgqIwO0dvHLryW6+DP8uP1EBN6I65
+gRuzOaD/O2TKcHIRKxxiVIIQrKBAFGfqrqqueNwtTMtmkwgxgrX5KriBKO1xnZWDWSuP7zP47d7
Xl1KXI/TRxrJPYymSSNdGCG4w4v/ij1fULkgHQge80nHt4RULhjfe308ZEAxsU9vqQY8TDJHvsho
PUxjsYPV/xs70YV2+JxYQRNBEgeH83AWfvwe5jEGbOLXWglmhyZZUG03lPWH6pdU1CRb3ZBic+BY
Y3XdXTDnzxg6QpvdgWeD9g2pImPgJCBGwaI2YDgkQd0B1g9hJXQsFCIXavyGShWuxLiGzRPHpK55
ix4+bqEjuFfrM4Jp55pcZbLAAaTJnXHPgKUEPfY8EbaPUGJ5hdt9Hw/Ypx2lTaLM3h/XX8JFv//p
C/RlbpIQSTuWsRgzyOrtXaI9YJS5t5GdzRdBbtudbDyxZAMALHzogAo+0TRQtL2SDgg6FQ7whiAO
5bHx4C+3pA2wjXI+yGwviVMZX1DHGzw9KT5P0jWMUA+ebu0TjSbgFvGPt3oq6ZHcz1Ko2eWUZIuz
K30+1DEIIlyfjegyhuVtEfcYQiKzjmykPLsdEyB11n1B/OXVopXRCcbF0XCLbq+Pl4+BvP9M423N
3j+wnm9JbYTaldG7+Rc7jTznT9X/GZXoenKc00L5JbKzjhHOHiqfMaRbFRZHmljZcZ7vDXAvDh1s
Yv//CwPhYKD+vQIVM+HW9P+TNWtwPb04csizYbOGZ8oeGD8vgmpFF/XY6JaPbAr5lmgY0zCRrmwq
M075Nm88njaXMXEXYmCK8wI7cu32gP7zW6oJWo5PhHeN+wkq8TOvG1pXk+x5WawSrTMIlOLbaBLm
UCCWnmbDge89cztgEXBty8jP/aLC3EPidxoNeTkMES2xG9MoCwUDXFVCmA6QsgxKlgqdcZ/0ptA1
BR6xEz2+Ay+sBsfQjDT9G90TWK/sOCASH26JaWn8iY8vRLaJEccP3UFK+nVf8LPsMkhsNQNBG9e2
x1Wsq0fwEWvu901bbRpqAIQ8XnkORNRffIbN38uT2YlutxojU9D6gmCgUthkkxyykxeZzmcctkw5
3VjsEKaqz46Nyq0KlQvFOOf7kvRpWExTEoaa70nVmlu78A7x719TllVmppoFZbNtn+SbXfYD0Ulg
lZRBcy16PdxSvT6Zd2RY0mCBG4yQbsNuySdhQy4w/gXarGDZayBGBT3ix5a+ZK81w9P0kKOBH/GM
7Bgs55olaCB55lt1BbLOM49S9XRTdKhFx9hbcbEtgwna5n8SPerTUjwRHM/bza+8qCosreVMyPQS
XnfXZn6DDuVd7v42NXQcZzpQ9qGFWnrM+K2HNTXR8oXhY6WbnBUaH36gE0kqXrhTiIxuynaeKYMD
q7h/1tv2qabpf1G4S+PJ/XjtSVmSylY+UgJ8DSxqXsR6I4TL9sHSd3cFzYcIZfD8lOWdy8mZRTO2
Oh0sXfAQusohwlZyUgvzwwgM7sCGiy3VBRInftBD7mI/ymfFK33z64AFnCsndXqMgwP03RY3CzPH
kLDtB/zWdvbB5kXUPs0mIaS1S+ySFYfgreDNprOhsC+0vwCrmUX6+chxMBP8RmWTaQj1LunAOExN
m98VmS8sBskgZpauSh9XNyNtvtRy8OIR9tR59FyNC3XNj4XCsdL+Y23J7PZd3ar/PIKCD+pS94aM
Y5TW2Dj+2M69boYauXFc1ne8lBUcSHsRpBc7uv+DU8zZIJXSEQY4ndNubm8JAkLuGEuul1VKvbhF
7x5uvWJAvEsHcL6tEN5+IaZIET7enYdbg94lvwmqtSISFRDCCjneH7oMO921uGLwkASK/5JIZcNK
IUhDcJj3Y7sFe8UEsYUt6XHYzCSmajTwDxyUzm7NRx9lsOGtddkiCWwsXXsNJMJ7A8tfl846L7DR
8CAfXRhHOGFg7AW8qm83OKSu+HBG8jHhJxJOXrpXLd7Kb5IlEL/NYcPZ4uSfwJlG/017KB+knps4
6tpizvpgGLPq7RyLl5ikdbvJHGLjX+ghtTdwQaLqeWzdZz9pUlE/20L6iOy0/mXa09vvuFwgKwVT
EgUML2fUX419xeM3cDr/l7BiKoyXjr4Si9YbZhZhNmY9yaBbklGQRZRdSsgcANHiMx/qqbg9UnIL
3dtRGko1sDyRjaoQ0hWV+3xW1/mqkoLkF1V0sj0pZFcqgUloj6ISFsxJIkdx4AroeEBZ+Jws/fYg
h6mpZndcqyH0VF84QR+wAK3e22LV1A9bNnp1mAvuya6WSspUWXLWRCtA1X8RMYsrYBouA05a2+s2
GpMqqS2DMraKGRA54KblQhzGOrjE4ber0Km6w3e2+OdINheyqazNQIAGi4Zd5CLMIPR1Mz6Vfs0k
JSg+r6TCGfh3NpS+56R0QSTNNo8Bz7saU0FfiMF/PSeHzTu9Q6kOJDUvcSUiveqpb9SiNk79fEJw
aq5+8S9Pkr5vKtYNCIIvfX5al56k4dGJlLAJ3fgfUpWH5McloH5d7+F51idOEa5cdduVQRiFfee2
jvrPn38BWycNPptkq5IAwtTbe+s1hS0fpcqr2OtFon51762rcJGGTDkIkPnUQiqWcr8lu4iyRV1Y
BwQAcdONv/ADRVKgZ8Aai2da1rSWz5U1rEAaxv4i32/0FBn6CiKa9aru7ALdIz970+t8H0D+palX
fQzvG3YlvvhCmMA4D2k+F1O5oIhNXcXRj+ZO7723redDaJYECg21n0TTItT9Xs0m4lnwiRyRhp1n
/hTnYHlGJo+XSaisNdvam3f2c+k6L59gNUVBk7NxJmzcP3vQENSbFGc7GC45CJlkV6PTJ4DID/J3
298u6tJmT1xPFGUKnz2TqUVNFb+dzS5fKvwxZMW+mCC/vH2Y8ardRoYIkD28MAul0MQYHwnLbFni
CiVUvaR8s3imo/XLNh/mZ7LnXfBvZexALZXgWomB3DCpO5czpmcCWzWr5kjRMBOVfJ4HlFHGwrL5
EnPVSuf31HwP1zOGrwF6Y3Zr6N83AIorArliCnA67WUfqz0yZadSX2/lqCbfFz4plOye8k/YMxD8
yfUM432NnccXreDi8eh4mOhZ41I3Km+YXA8tLT8iIfnQ290UU6Xv3bgoWma+IXzGoh2IpXyN9M7F
xK9fXxFBuuGIrO6xcdB4lNpQSHujQ7ZNfZpvEO9AvewjSqDsgbyvRAX5Aq/4eNVvGREIXum1KmG1
T91dm4YXtyEXpVO2GEO9SmlHQGFV5qSLj8jEF5o5WNlbdz7bPxuYNQOBjYt9gqHuGcaqUYe6RuIU
vmxEq+mrfk0C8fPqR6AHcqPHV5oeW0GRJ/xp6asXVIhGDYI9pwKyU3YTSRIEjdrOx79wvc+UzAzP
fV+dLSOzJVylloM6TIHoWTms0OmMEScHOrq5N5FniJDo/+JHQFHdYRni1HgCG2atEG2gR8rk/3/c
aQF3oEXvfb7gcIcrmSh+HDYCHnFfaMuzfChYFv2lj0t34qLJR48V3HF2+0naoO5lvhTvQUNiXEQO
u2CNpo6hsoppOfNT0RfROaEfo8s1E7sGQ/OtGSZzvqvOe+zbFRsurStm/AyDFXRR4a44lyUWKPTm
fEcwcUOv/z3hZCpsC5AhGJbLJgmOeLwEXh3MAVFszp7+WAN0dVhuuI2xretzSMYQlKyA23cHtG5h
rJmxVUNaUBkTtSUzSleNeMd38XjHinigHHs5pCezxscqhmtmy1eYcdzbBfBIj4r6vIy6LNib2LXb
NS+zycz/o917UgHW6YygYvAp7d+26oOtYs1MKOgXKCzhiOnCEAY9xmgw/pcXFs7ASqVPxbe6jx9m
rlnotIN7dqJ6Z/VPc5mFDT6SIpoq7y268ZYyPDm/oAWFNhUIgGj09OrUF2qBwIXMEX+8wQJh5gxg
nU2B1iD+y5pUO8mvjtZq7MHYFfp6xC90K5AOMBSmH11w9Md+SGx9r/d8GtRAyjlzF8B/t+PP1nX2
YU74xJ/65uCZ75X0Sw4k3SwGJR+FbAGYj7L5do88FqvS00eCZbtrP4K7a2ZUPYl4X94M09ikEzV9
rqFywccREnn8yVXJjX/3rZR4C8SNoKzPDJ0kvRtSCin20yPTxVMKGChLqYG3qcAaENQbUC27i5iC
JnmBSy5SNBooxTEdNZb4QKVhefFW3/I6Y1rn+z6ly1MrvpnJHzOgQMS1Ang3+ZPPMlknyL6opPQ7
zlOTcQO5Egh3tD6Lb7MhJqxT/LL8JLMhe9dm95P9yooXsbT0FkZ1M7UMDR+g2VYhe6HCV3LrvEpm
RYAT9zfwXBrtZZAcmVbUh2+lhymhpT0DOJOFKRTpDc0TnJwo9TJmUC9fvE0UHz02G2yht9/r7CCw
QtKgYYAXPizHyITbNMvDhFqwBV4wjQYR9cYMaxTegg80LvQjz5lU5GNG1o0PNoZI2qjyRbUp0cDx
zwjS9d7vtlrnp0qe68YJ3mWIglElQb8Rtbx2CXy8y6sn/v7FeKwasNmEkaNrHkwTq+zaYV4YS9N5
IC6dYqgntoPgfxBNBsLJQhg/5QqmZ7GflnhepAnWV2zQUINDN7vkgyj+v67xFWiTffwUme4/obhX
AIR0ZgGbvTd0MBgHxzP+mjiUR/LVWl+VwWIdc7cdxhfCp+/cZrKuFH+KspxPYuT+5T8pzaTYOGpS
DeNUbfdCXNwqjl3zoJvrrTVqqWMTCHbyxXjfwRhVF+60namPilcMdM4pRSKiBMD1Y17foWpvYDi/
jxSyRWsxc+Tjt5ZLkquHFZ/LmiXt7T8dlwLLdYDpyxZohlW6Q/3x2gA/pOShZbXaK/e1GS1X4yDR
bnQlDHyuKGUGN3x1MXEH1NArExd7GBuEpS2SWZXJ6Z+SzTy6xeza4Llur59s1QybBLdQS6DnvU4V
RfDkX9072AIFOX3l2M/9g/XMHLFMr4qK0w7gSXhyTi/VqZMHmd/V7XourlPZp90tl1/Qve7exTT1
YFvrvRbgRLcBQ7WSdKmBuG04boX3ej8LQW1C7zkSZ5mYdg5koj68GdnX07iiqCdUa6YL6ZwRFqgk
RFVyXxw8inGZe/QHYneX+7L+AaCwJMor6P60sr6+BE4Wtx4Djk2jou5KHsxFzlpTNMFi4K2Md13D
vDhvhuz6mRJ3C97EXORe3+zQkpH9AUbQi6yNq/Or827J6hnx865VQuKGHx3mrIEBSI4oPZZtutFB
9ABLsPo8wJwWjPfdKSj3wZyM517xC3oeQzqjsRh6cQFYE7B0PBt835e9ycRrVBHD58o9ci5hfWxX
SMtVD03p9zi511IZrMRpfv8E4nAGsvlVpDnOfknFtk0v30/xv3agY03NWd3WgvbvPa7fEco5PZ8X
7CTTY3ZOTjnhMKfzUfYHiYPHKqo22QY1RfDFFLl6kQCqx+s9KwzogbC67m+rrE6V7cvRyE3MEyKL
lzoNVfV553xWropstrWpCiZkldRHSDUEmeTZw7muUXxLvs5Sv9orc7IfH8RRWZh0hdXGKFZWPAJj
HUqlfEiA4QYGgTOaNQiQL6QCIe25pu1YPekB9URiWVBDQG6AnK/SBMRc68Os35fD92LoZyR8vnZW
PwmlzkzEjVKflTznV22r1BrZtZ8Uh3giUXiGw3qUm/Sp4wTD0KN3rs5C58xkC8gCCsZTlB/wTyUG
3p9Vsl94q+G/PTPKShKcBmFN/VVhDglrcvoIZYDjf60r7k6NYAMb5YrzqgftlQyyNT1h3NKlt6Vl
1PDE56uh4gAQK/eUFweb/Hx21OoBC1fbaPngpoeKrmWszlbSLbMra61bjMeuZ/btY7w5PaKWiUs9
GOzXz93xVmxA5Tmf6u0ubSTRrijjfdvEcbHY7d+GzlJgQ0GSnXh/yswJlmg3OfqjEHvCRElf/kUA
lJObYzttWpBWobjLJOyjzCN53n/z8sTstkCOy/0xd49UXUEoIQ8q902vVu+6BR/f2lGb89OBTsGg
asv3ZkLhsYt1ZL2CL1twJPAsT7tMjOwa5qgWrhy/cV3x5rfoZW5UBdt5B57KaBBk8N1WTkCHYO+p
nzQl57OcvTqdvoe3SG3US4WFyqnZinoBWPU3Zjg8dJt3RNmdFMFim1OAqguVfcgZB6SZEiu1Py3N
sAkIFJDoLFqhR2jqM0CQgPUFohv06fraO5lsNoMMi+Df+qSqZFfhPELLux64ui2ibMwwOPQzNJP6
r4rnRVs5vYpBk3BlZ06iXgrj4qYQVRs0kca/vg+b1C3OW/45cwCNvDCmW//afrN8REXksTvO1LGg
kuHmilWefrSJgmvPCGY0dyFkTk2GXNaHC4gTlZVA//3HuIOiikq23xKsoUOPgY33D2ssvYMZ3uXW
cwMqUMY+F5MltbPFt9fFc+QebJXTDPnSIfwL7gTwwW2+NYEJ/nMYzfyGwqMc0WBQ1oTLE4wG9JGO
ZNMjTVjVF8Xu+gcjZDHGqrRczULQio+eYodYOHW6bPvd1L+C+ku8Q5iKDua2x3U0ko4ueowgMV7m
E6JV70+SDwR+FifTWv6CCmRq4btmstDtllR34izNNosK8ErpGogse4+qgOobU3t3MzGZLRbcoQNF
YieZmVSTQtmYQ+E2WaNUUgl9BOrohtrZ2lAyhLylfT6XqRqLwTsu6wdTzcmcqGmx4YxIhMxVwg1F
CxxdzkMvISctYpTYI2SMWbm2iOjiKY5SSBzp2m+4y5Q8qRgVd878CzFgYtri7K8JdEXTJPz9oK1B
/tiTlH9g6Jt+21aCxqBzyTM8fW0raOeXGJy4RcYbB1JCCBXdeXGy+D2sSHGygcJU2ngR0WchtTbO
I9qyqMMcCwkO953xNO88XJYDn5LjLvbih5pqDvcYL3XAMi5lwSQ5HFiD0zHB1kumHdmkSGMSCDT4
BZNGOvrjA1t9bg4tQ6bJ32yDUYMVHxfUhFcc67IZIa62oeSbKybUboylvXLmtih/JdIzvQ1tGaiN
NlIv3ICSOLEzb/kftNmck4NoD4QGJhvznVjC9d0HjriK910R4iVutNckDj+do/GQYvuZAojhFApv
EsrjOWQkvCdR03OXIGynMFd6hyob3Nwh4lfLXpx9dEPFLVzu+V+hhTt2qeu86n6DzLXeOfL+g3JK
jMmocNantD093uiCp5avm08o7U7FxoJtyCqNjRa0RSwo3MhpHp1AxE0/+qkHES4eHV49Fnf4XkhB
75vGbhQSMyuILn1SMXnPbOGJcc/pvUaiCWJ3yY9GQk3Vwb1lcMHsRIeBhrVriXTGuq6LAaRMiGSZ
yGJ59tj86OOHfTIoBqizAjzG439ouWDLQynqsvChIDEGr4A3gVnXlA6VhKXjFPaXwmJAHa0SNyCp
llGZFxN0298udfDY2WKquHrVNrNV4PyM/1Qkqy/AQLY3ioQi5jWFrMLaky8lfyCljG8oQxmTqsv6
amrvzgEJKJ/mQoIHm8GR4EerrEtgp7HIZ+6oaa79141FQS6rfbZY/qb04TNyucnk6dSiZIUzxGHf
FWrN1XGgsWozdpsEInKYWIx4qVki+WRBJ3PY0w8Enrt/PEaQqBO+FCBe5UCik3i7dtoYWonx6lto
ssCeS7/ru051sq5HNMpU9v3CO2A8FoZwSGYfrXVFUdvtCDhIpUlqLnDtq3iSpOPZ19UK/zdIyukq
wReQLmE4fC5BNUnGuU/i+5jH4UZvWAv2U0uVAWoQ0O8hJrKfXEjK3x2t3/vH9jbP0Mv1vfsgZn+U
mUm+khhSi0TmfKH07Rglarh09x1Nv0NXAZo7frPVmqPsopPdS1Jv/miPlZ06V+3bSFbK7SJ0ANe5
qHbkTmqN4G4E4agZqK+oFiEM8XUoKsvzRH+N5c9g/3JkRpNkVA+pCh1WBrmPvD4wVYEujopvBDvI
78NV0VfqpL9TorM0OPNSDMdWRZHpUor+L7Xtqp1UDkFJB0NsPQRraiE4OzIsTtesqN/Dp/vxLj8n
4wYGJF9OEb0qoqpDE7de0jkVVXVphSfNzKYf11KKXmKISMQcJ9Ch76OxdpXjbo9cvUhO9T59lPl6
yde52kZ+/I2hW706dylkQhbrW8i0FPuFdMCKYjtIhSMXODA1sCyAol1zxm6QQYgwHUcsivRLDkwu
jj2IF8Hq7ZzWQ2+Qo0n1Z9sIEqa90/wrCePv4sbQYenwe81j35tRZFy5ICfMwEDjew4K8+KWZu7L
r/EKuHEE1PybCcHWuqpZRQczMCv0Fo0thYsKKNRlGqsOAE4+GumbhltfD+2CEWFleq7Qr9cU5Imm
bSjx630vksDShxavv5iJxChZcpV+OQTN/2zZyHbTxjfTi7sdG5J2WA4zu/0Inb0AV2CZpg6ZppXO
fga91i6xRjA6w/PuzjSW9UBFrkPmPUWI7lDARBCGAVr4ju8pWMATOx3CTMa4ePmrdYLRN1hSMJRP
U7aw8Q98UOCP/y1noL19aFNSlVXST5FHWIerYLrC7c8yFelPVBFrcxL2Xg2OTSCBdiWVBM4U35bF
sJeiCyct0/DAf1puGlcwcWy5SH0qvjiJDxgtw5CHCIxxoGXDMaplYRiTHWlvj6ZIcnHMp0AzwqTC
5TLqobhIEypQ8nq0HtkRBEi3yxPnXt1tKYKGRLgQ/S3KLt/2GXMrw0qVKBUUy0hCJuNi7zF47M2X
VRqZK7a2pBKv0r7Xpvk5XOX4EWcEXgZ+sc/K/sJVcBtLdmgq7Pz6kAlHfrW9b1hXL1EdeoSOkqzw
bIai72dr+GBk5sduCzKj0sQCT0thai0vJbu0rix/e+epeyD/gpQkuBk7fxXm0E4guRzXPgU2wShK
uS4khz4NAerxE2iX8JUggLsNV4iTTxmlvttt1nz1MreLFt7+FZggYLiGtDHi34eA99ok1v++YnDU
tc+grkJIz5vR8o1s8Hp7N0Mjdddg2d5ELLkUFb/CE97RVsGbmoWLgkjJmokiqAjvBR1K4cpW6PX2
02ONN9oO/nTkRzM3IzheSEz1ahFyXvNGrxBgC6yoD+5YabS5hDrtINtHJH5b5nv8tj5PCRaT3JzK
ASkvoUUm3arp6MCBAtdrvP4Fsm1qo4GZDpZ8M22561jZ9g43D4Qi4TYwJpePPkApmtSm4ZUykpi6
qnkn7RKnAVUZQI+ZwYRYPA/FQ8sIj7R9nRfGWZYM9t2VFT/3h0yVLYcHussGT22hEwthYgPYwQik
HnivRJqcWqshZ0QW4jZShuehvS0e8tU/i/AvVpgiWc9MfbSYmrVOz4og+Vvt8f+8dz06C+rMUEFW
ryVKOGjIMp7SXzmfW6+w0p8jNr7pG+jn3jDXdfS46mawsiKCTvvXiVZLZPn0w27Whc9J0RWNkzct
U4Obyl0gKSCCrX6bzwfNKr1lB9QdtbcJ56KPEpqzVxnE5uLm1VgSeH82tI1Q9sUcv2y4NpHod8F8
M8naixE92plnatrcZDRaJzAyFhxrBMtmpVgJsFZiWmlZZEipOTCRcdp6Bdu7XZD7KVr3I5ch7+80
JeQkIGAikfg4KEhuyH9FBFtM6LGv+w1mRRB5OI2oYrXWx/prhqq2Te2heygIOQBP0O05rIYgW3uU
oglAObv1o0VNvgt6qT9hhVQP5QSkWvX5BdON3knetyC59xTg0EJ4hit8Qxy8BrJTc2IAI8pKoDXX
xT5N9c8agop3kK+59sw8JV0cvMhA20jjZE4io65DXpDYzo8k6uEp9jTutzJHjid5bbvw/fw4y6lg
UOkFSeHOxgPG94B7Ak+LmbmoeR2PYU+3hZURwnVmRHOXF6OZKpgQBcnrsjpmF+R9ii1DGXMpBtSS
MdNZY8L3fRNNrfpP7eYApifGIp4hwRv3F/iS3bhi2kQAkwuyNhAN/RK44nSqDJAFueHqlYt6+LXx
jW6kRXepr68NtdgNdga2ZYIwP2WXQBs3VJujzqxY+Wvt1ImiBnsZkZrIam8Jef5+Go2HjhEFQB9Y
7nbrTTlmGEn36xgzAGGHmXlb7t6WgoZMC8MBvyxYcXrFnSz54W3PpuuJxyprgKuyUskZSOzOHKfT
xcngFJ+D40OzyP0Lv+cxloKqy6UJSDvCjv2gHygLFYcOZzy175E+MEPZ07bxKmfYTbjmcfvq9hmd
qB2vhJSa7OMgqC9mCmD/xCEw8b76RC8v0gcRs6zB1YVrh9RnA63/xyOBQqk57xz9mEFewBtfkIo+
hZivMGDujJeau4YKdVQkrygHbhdqNqpMEoj4bL5VFyDgS34Ny3n2g3K/5QvYKPD2bKJtDvJNUCyh
3xOSuiDKlo3/eqtWYbNHHPI2tXUAC6HlObuT4tnttHYi4e1B+UW1VsH6UFpR4ZmxVbUBBvOT9hkR
z6wR0DIcvr9EYzBdvxrC79mymH4wbBZfMe4gUIMOe49nmRV/gznR5P094ncYb+fjbrp+VM+KTem9
uuj4wn4imomllULOJ5M0yLF+G/HaNjKJNm2//mSA5+Aa8P+Y2hVwO36HTidxd5iUJL5CecHafMog
6PBiXD7NSEE+Uelm/4OwvOSq5KJOgbfUhkTRzlVIRpHxi0euXQVbawc/vIBzA61tmjnj73c+tpsX
qhU06EXdV+pM6JilCFnvB44cvwL9NdV/YWhemvyHcwZH/Q05Iay8bta+j023jp77Lp7JtKstFiO2
w3G1EOJqajTIUwc+TaPjGwHqWpTMWRoEIAxriWrdw8JdEKw8bzubvE+Dk1WzeUPoDaEzrXQCC3Yo
dLGEchGVsuoWWdh3SfKYM1u+w45Zmh4jF6lwc7YHsjV7LaHVF2WMdXmQv9yMZfeXlA8xzvjXlFNs
giEC/e26reDa/+KZhDhQKIDJx/FdLv8ttRPEd99q6XhpnLztUclRb7TbI0xMtvljZ6RWL71bJbXN
3J8G2mRH+L2tiwIiv4RJqFWmah3SxNVrjVj0uyA/imwPDuR9iS98jbLnX9FREohU+tGY9Xs1qdVz
PXn/3fWzCrDDPzhrCyppetPt9reFewcbQQpJYug3gop4z8+gkWdt2bEhrYb3bNbZdlUSYSe93z4n
ElrTuJEoIaEDR8WDre+u9qUSngLQIw7M2AGmuHH6lztXg8Cg94Ls8mKmWBaz6iiO/aeJ2GdEezH+
h9kWNEShuJvIEm9sDvm0uStEILvNoo6etLn6GW/2nFrDn/Ot0SDizDMs1Lblyj4i8cYOT/MBbAAX
r3uwYOXJJDyi2FY7YaPgoYBb7qaUMDus3bRZREcz9fLu1l6hUtlXfAWY0J2dDvfqNUYUmQ9vuBOX
pnTU6RF5rFCdPD1tWny3b/l/GkASn2+UsdNUX1eYyRTulgjFHSbraZbhkbNo+BGIa3yb1D6IqNnv
TNL02uFAbezW2HFQtHExqRTNFD3QBjOgG2imv2+OVCjBu1l6km/CPU9xLrt4foB+/2o1O7W9eiY7
7+C6X+QUKFp6nKcO0X9OFrBEGuzkRQOxxAAmWTIJqxPt9fYK9kr9cpbksRjWglJ9yCM3sqOoGEPA
ZLRHKAbK2s9Zdv1QHXDokR5q5iaq+y8JnaewxD/T3youCDA/mPM+NAhePn2ulBmxgZ0u1RmrbOnH
DmHJoXIZ+5EQOT+Sd3c+y/o2M4Z4+D9FXAuH4+r4jf7oyieenYA5ryjLdl9KmjLUexPjJNFwmc12
qCO4lshxw0Uk+jp2KgF6CmGp+ehxlNJDifEoOdgAArcireh4hwie33ZsD1YbPDa/CRGlbPDuk2Zc
ss7PtiS8M+OSBHAWg6dvNX5WRrSTrUTISidHVxN+PD7nYliskmkVVAl9uYcEuk4d31FazQY3SY5d
u8997UdHW9EdV0qW29vRsneNCmu+xS2u7nPmIBYntkXxd5xukBVPOWFY5UhgD1Z3qMbfE+QOMM0C
cdmC04ZsJ+B9rMML2d9pelVm4x5Y1pIbnJ5LLb9Chxgh0ryvEZlXcx+EcE1YGkROMUIPHU+7udtf
HElugncdpKJfCFnviKiImjkCfN7pVxI1xv3hKJ455WWnmvK1h2rktJbzqG6nK+V1nZbtMmeOTHJD
XCuAa0ysxsBL6EqpaeEchz2R5aWEyJDhHo2+RdPCJJH9+76gf4COZezRA+njV1tQod/RURCDy15O
HtlkGkLg42q2QLBDf1bV7zWyNFUrXGGGFS5fCnsL3fyr0rj36uv8SpSr9nPTbXgwB5KREcK7o3mi
rcFL6jNwhjBc87M6dr9ct+sKBuP6NiEpjqZfE9XWGKdgQClYdL0pVaPjFA7slXDTs6AQQuLrKnkn
tF6hMPnKWffwP+5fUez7te5URydeamoWN3mO8CVUYXx1bil1FRPgOkin0kmAcJd7hXoS23Cba1VP
q92IRpKhoakmU6fhZ5ACZsq2kyrkZqjH1HvLH12jCF+pRxYU57E5S4cHyvyqj7ZikDSHliBDMLBH
ndDvoYGGI05RHtDDlbVIaULYKt/9FS8r+mqhrMpsh3U6Ut8OSKruFESPVPh7F/0zJ+l+T88bU5Wb
RXn/Wk/nXF9+ttsI+4HdRH6ub2jqc676B4s5eShcbpCqUxO1CqTF6koEolzs5OD8Id6d2sujj8c8
DzRqMiuyg+bJZZb8P43y9Yq/t1XWxbziT9Kc86fV6pO5SSucZjXMue697Fxkg5lBYkpk+tNeaqzV
TDRtjmQoh5figYgb+LwhI9lKFJi+8+9owBop+XUVq4jhpOn6LICm6VShMGL6TBnKbWB+Smgr3E7X
NPxtn/79Z0m6ENUv0Ng8Tk4P6i6ITFCmf5551qZgju2OKRkveksMTNpWsRQIlK3AwzdJbcu7qGD+
dyJkqS3Q6AHNXrC0vO/cnpttH64cM9xk6kGf417QcbZ8+bEfnxiKhiBLGYBsp7UQ2fH3G/mcv0Rx
4Q5WOBXIYHkdNzLR2SlOsYLTNJNNu3aDbQY2CPPtx+qQZDANUCI9n1bNzdBHpJYx7ST9kCPOrWIf
ogtwSl/JOaPAdkXJq21fO4+vrcQJcNSKHMWtV4jqaamwUGEcOmWRHB1eNvh+m/CkxXUdXNoIbOJR
oWMUGoxeE8yZA2FzV7yP8GU5CvYiPgqlnjjNefAuQ0virtWDR3mF6+zuj0q38uFnSlcCdfcSnmjI
IehitiDadXcqyfKCpXGrfpLObZcdXgG3/q9sT7yGBCHp31DyskIoQ0enFxihtHkcc2ZhodDEjKeX
hdENBhboqpDjj8nCKI1b2TjiTnieOa1WOoX5rrv7LwIzBrIMNtD0UngnRyPXj5zPB+puZgygE7jQ
+4IzUF02P8jIaPJauVwNEXWU3OrzavKmK6ON0DewxAoijBVIeF77ijUwVRA11xzUOZ0MbSpcS3JM
xfExqElBAWGYYFxhb/s4GFNrNNbsU5wtdvVTQF/Zx4RUzCbgV6wxp5i9nb4IpQFLTXxmI/iwsULr
0juUotLXwPC0pLE6FAOQe0nbcm9+FQYZ2BXPwF0iIkSl3KSR2hfbB8x2dIHM0Re2RLUvAFS7oWXa
1dNeIzD5FuRnoP8zGqAkIRWDvMIB77pcsYcAu70kx5n/hQx+B6JUuVKBW7Og6syODOp5po/Nava1
9FvOyYaNkPQntetEYnz2KV+pbtYVZAZdwAOx+i44tArETGTmJVxxt0lE4txwanygof64zyWMurPV
gDs0Zae/PPhN+8+IlvBT7F9ZHydWFBkcf5tdpksoeByRrxARINM5TTFkcUkTtBPmv67yNOs1OKnX
LYw6ODMpQiJI6S2JWSRYQBEl2ydAwAiOq5tvQrI7976Pv1cT4kQ/wHdqQXPoLp0C0CrPBXh0gUyI
9xitL2/zD/5ZpbcRmcgXOMOjzpWe14Kqe8U1Qt/G8g4xt2wOkjkEOY9kyYRZsOT7gHJKau8EHnaU
bJFhF7FiHGaZ4ycfV0WAiImg1p2jYLzMse9WMQ5P7sOfrwz0JGFPQ6NvJQPb8UIOy8F62wfDVap8
5EW6rxLPcL4TJ9OW83SYx80XYytnCDo30Pm7d4b+YHrCRSCiRTL+75Ruj7+bS60jDFj29MqWrnla
nI4eIms8VLDk+mDhbc3DhOW/R0nFcPYgSdoDrfyXoHcQlskEqiI7nT6JTXgwps6f2v3wvjTs873P
v/r96WiWG0Bo2ea+jZLBYKWlPNRx4Q9mogwNBbCvIuGjIOjOgxoKbFzTon/+XfjghxV3keapip7E
zkRSWB2UaR5e8OBQcNMAwpFGQhyn+GelWZ1lXGujo3zSMKbTCCEcHE96x+Dxl+M2q1FUeTFxc/cG
ohPMNNwKlT+pdu2AeP2xVSPcVYsUWrYSYAU64iQ65T0fuQUZaNtTwQWdu2igRRtEMhDesQqIV7GZ
1lMVNZTqjbAm0lXfnFBkB1wiE4UUusOP2FTewks9EREZVjHTWwT5fNgui09ITCJnnJtbpKPOvG1H
K8vkQs7O8CRV9ugcCac3PziZAsN+y+4OC6QYaKnkEa6wE4sS+IdLNG9xAeptk71wySDiI3SwEsaz
sO+nFQ3L7ZqDexJGgryA3Kl/P2gE+ushDgJ+zLmOM//XsfcaHXhJRmmXciOM8BGGs3eB5WarRbgP
WyO+JkqjTYTdrkcbviJ/ewYtrfpvAzYqbifBwUVfu0wjL71eumU8pSYflL5l5kHbBWVormVnoz2a
etfGbkeq0T48VTOvZkEn0562VlFb7dCd+gIycwh4MxMhDjRrTt7RzGF3dvwflMOVoCoXV+rVCwpb
Gn2Y3hx8nCUhspdZ5ze9SBUJrr+BZ2ZaO6Sf1UeA26WfM+Ts4/2xDwXI9VYCQBwdQWFEnZQbTImy
K1WsSPpHQsjI3UOkzqeio/XSq6fIxNyWgHPJXb4760CCPd/+SpvSfigYi0M92uev2ylAn6PD7ziH
1AWjyGz4yQ7h0w6hGiARQ8kG5PF9TkwlJctrLOqiOWJ6nkCyvq3FuZ8czPhOUSCH59iBRP18UkA3
1RAapCW66tGsqgLUo/vhpQL9PNDoWkQKeoYC/QN3o4w2szWndKzbHFJEkUEhaKUR6Nt9ia47RS5c
/pJLk45yj+CCf/RgDUe1tV6F0+qnBN82LLu6p6K9gB9IBjTt6bmZgWqd66S65Yasu0ioVGR7WuYC
owwRIXc6bhcrD3cWljGwqlZNxbR5QzTFdsxLPBs2AivBxHS567P5LZBrZjamBdKpEK5s3FxCzPgQ
VhfogG+43kfMXCz3XDxnP55f3C84kLoHq/FMky579Q/8DLty20ChDlgAmjaarChWoq6w9DkzTHpt
22u8lqQ92FZGLYkHlnA3e8zP/5jtIITJlP3pae7Qie6blBukZnphp47u1j6UNb5xqYTSn3qk5nvB
2YhFSUem/y6Xg9BXE8D/myWa2/KPxPfl5cfdjhYtaquG4k9yreKGqasrm0CGYRYEMQYycC/newG0
4co8UWd2D24y63cz7XaC8+xgjqDJXmAdoZ6GZnGDsVStBemlC2f5GHPR/lfsLCZyXkKse180dbIa
NAlcjUyl9yj0MyFzAutrFoVEyGW2DgcZQCWWEbom3fSrXXuCGISLJNxN2vzRrmFHXtbWIMOsHpgF
mVA6p8hXbPrzzc9ZpDs8OJS4RZi5oIesofHvvSc/Mb3zrG8bwmH8j4ivOIBfLfrvvc+qPG7j0hWI
5Blzq+ops3ipspR2ZgteoZjn4q+yFzjwbC7PJugtB5Ob2cNBMuAedkdxeOrHFDtPn7M/GlOFa6+N
TOwaRyqxuheUb3u6Rim51Q95b+yPIrqkxejOWavvdVvJPwGIyRhGPsytXL+MHbyq5kcYzPkGx/O3
iyXEmZFYxo60S/ejiWlNrITrkBbsbMgP7O8XU5cSgKevobv9TLmsQLeSs7gPl95DJTnNAbItcv8D
hPF115ZRe94R+Ro4xYgx1Ya198tMlZ97y8CePaERU+q4KgAYKx9PZ09f15MaeFLuO2NgJtpNAt+Y
RKiVSnBYpBaoNDPoqIN/rL7s269nR1apGWFnh4sW9reoRNl8U9zW/PNModytBNSLJCGOzMxT7Jww
fo68RqIHcz6ZPMdawjFCpoo+Va680RAGZ+6sMOTUIF9fR7xT/TImwqNozdqSMJMRxzHs11Tw/Efa
xIfmgY1HDaPjatzR4J1i9qw8NTZwmb8MDoAva1JRKCmuAU6TmcQ6ZzSZuH8A+DLPG9uzfbBTmtjP
sxUDbtVhQ0FTqqXwXwsqvBrzPSwZWQN7qr8D044uNfk5mnLhsALc1khDbrfJCSZE7jz2NjBVnggT
DiBb8mwIzdq4Ugw8p4Vzk5AzI6Z9Dfjda8KgoFWa9X6RxWjO524bjFgcuxZu+zDB88kDh0sKCXog
SCtE8MGJHiNQObTVZMLPs5U3LFbZ97orXhFc93T/vhxnMqNahq3+edzeg3AwOJBx70pSTnqO4C8P
V4P4TwNuwI614y9S4OfQn7WHhvL80IP3JZnqYV8Ib+TjD7GLrMhAbALVxCHgvyOeTaBK/t1WlWQy
4iuWX0puh6v5fkXizYP7oUu6oi6iwbeSoZ/K22OwBifNHGuKnqPU00KVOfbhBGFzf2nV/SC0BbFd
NjHfJgwiMdnNTDalKUTkAx29hmUfwpxjHSgT5aA5lTzZTjbfwpRhX/1J+z9bSQOrrsoKqLZSjhPD
P5jMsYOGMZ6HuPUjVwIAaz4mTp28hTO6cTX2V6o9jqTfWrXB9Z8ZigObLVW3z5XY9Jg5eIs13D7o
UzW6q8lkfhMJz0QnKDl44lTdEqU6DYh6SIWV/zTdSa820hqkbk7/ckim7KETA+Rtgm1QMG7Ur6XB
hrj2x6WetJFAzjMT16e3BPMNhwwo4nLKw6yd8WRCfarWp41rneAjvSL+gMiJWhx7YOlPcIy2131T
SVPzIb4zHop3zzSK9MGDYgTU/BKrvlEWGLeAYKsXREcvTRPvh7RSkeRtXONQ0AGIX4Jd0gh7SH38
3ZKgx9VVa0P3+Xtt3molJFDmXPcfQgIOOoV4CKULituNZ/JVXnfNbtQ5WpVwZmS+xJg94so9wuhg
yeMX7z8/rOx8lrWSNm0LE8c/saq+gmraNhUa1crVLrd12uG4MYIGBzE+aH6jRpaCVWCnMdpEDyNu
ZF46W369Iiv2DlWCK6XiMoQGIgUY5GF6HO1HkvBbvyPW1MR3J49aMGehl5BPClUedQAMKDK1PktJ
mgWyg8RuBVxtvrkE+ePKDIPxEWWbygn0ff3nTIVmRlNUW5rr8DKd9ta77yTa+KsmVKQJ+RPiyMfB
pCJFFvOG9NhJ4SHro3QOQqQvKCFGRLuYevBQTN7ujDnhyNriRCHjXI38ZrywdB8MGoE+GnZu+IhU
42dYFCAzDvVmBDe5R3ApeLbq86YzGrdoZ87u8E2UUjWpJREqZ6FZxBfZFSm4e02dra73dyv6O2CO
ZweRiJR9JZvvxNvuDNx+OniRDHUedcrs9te5WEwKSSiB/pGoAKmKNOpl+gpLRX6SzGV2/ZzoTMWZ
cMHJzqs0gDahJLIOM2ORFGt+2c11eCzr71VdKLcnG57sbHYt0khBAKrnPwxi87XB+ef543Cv5GfS
EV663C1JpsRn2so9lbfnOCglMqenSSuCwDfilOp64xnP2gBrHzZzHf9WEaeE8nL9mShC1b9Sr3ly
mHFxVyHceTtON0EaCX1XfDpFjD6Jj41NAWBnO46HnmbdKSBCjg4zVfomhKXaaQiPxyoY39y7IUP7
oyVfT2bc3u4MK4Cq/rzLFPLw4vFffOc6SIH42prKTwqUxmEdQxgpwaH99/bV38Vrj4/gxefQD9pt
UzwNQbZP9zgaIrPPHscUxiAAKdSiWdqcXD8zf32rBayPA7ibnpavU7u4bWRYxHwENmLvGoFl3yJd
EWeTtgclXPaEqPclz4yHOAuiuuXYGQ519TPJRQdKnMYuceZQNTxzRKIyoUZgNXjy3RbSAatvP2Nz
i1CkqlABiAabGg7iUvlNx3mTJdoUJfbNjljLTgQEzsIGromILZbQFeOYxQePwTplKn/W9V4Zki7d
P8q0AgjB5WTHi8RIUITAvfcqJpM/e1loUuBRJDPqe7QcGRJiKsWMv3Qx23ptJLQ9XhSb8b8BdVmA
o16bIQL/jjAA7hDO72FD06Sw3wGcbTKitYORb3ZFk0dnplG8S7+Eozam9UD8gcb/JP/aQflxdn1L
N4ua3XX8wtIcEyHhv4AHx6v9CJabjoIrKUsIcq7RAWNWUjcGohSQo0gONT2tsRwktq/7/2F4s8m3
TjMeL2DyQOSQXA73SIFerRZFsVoZRGau+nZhqSykVIbt+RT7smPN7NcnKTzVnG80pA1jc5TRhchb
/+YfaFy0uhmEg/WcWvKr49hjBHga8iM22qcy7ByjjIGJrQlUv/WJv04w7tBdyOd5o+VqfmEFEdR/
4nBHmcePiKjbYYpprFfmPGzrFmFZ2VJjleUKyqAYAEcUBKfiOVVDv7chYjUhfAKxYPgjEHjDhxaQ
pAIww+8qhUIUu0rk5cvsuTe5wdtOX/1/80Tj62MYvDFe3TO+nVG1egPbN4YsrA19xedlWzHo4S70
KNNotmzmj/QZ1ljhGmQ2sac+9LFzOC1b3OGhCt/8mssiB89D0VV7aNKXnxyXrFHl1ZgGZOiYO1y6
u4ftEx7WvS2yMV+fK55vROzP0F0Jp05N23qCqF5VljuUxlBzNXxf7JzaBl2ACUS8WWqjglnEJcqq
EBu+I7CtfwYv1P7GFqxeBwA0VX6czbMDPdd7D6+Lzy8K2n26YpnmgtrDrJsvu4yHKn5E10M7aLfa
wJ4ubq+NpWYco96dlvLcSt7Q6XQ4nZeNHOsu7cUPn89rcNpeonsuc7zAUNUWxmVtkMJH5dQENG8v
NLm+btnA4sPqZBVUbzo2zrwK2WM2Tqhaqg+LwYP3r+RfjDlWtlKPuV3s17TmnA7qhW+FZ3uIoujm
QdgYgjEhWJkyuqAQTwD+VPGjzLS7fTsa3dL5Y3cRwPrT1IriBbyyssGDxEdo8D/pmMLAdUMOKp3H
pcwu3TZ8YYI7IwinJNLKmMT2weEHYABaanTJvyrny3OEh9gRO7wt91ijTf1TJ+cWsQmW2QtX516l
EapZt0aiBJedWDp02KsjCCXuTl994gh3W6aBORtJVKD3yhA4p80U8xBUcsNfP30+FP28xj6acPjf
A5+kPvZuenzZCHMtqQrBOkkPUVT3LhYNj9msDZYTLSLmS3ICrezHELFDKGs30K9OVWbtQfau35UZ
0Cpdq+CK22LcPQjr4qRYXWaljEOVwQbwZBDJFP7F5Z0DpKw9Ob8YzXOUiVLpR6TzqxwV+YegUdfz
CIrnFuHhsbWtnODL6CjZqIPHyNi6egdXwRpbN4qs1Mr2ELvHD1bgxISK829r/9GV9OC/ZIzhdYQ/
xDedddbH7YOHLK9KtruLCqMO4b6FYCZTmtaCOvRt/SSPvFNsdFwO24bQiRliyGvb/SIHJi/7vwXF
K6VnwJJZr6gPFtpmg0kFuO0M3bFbv2s19SnrVqLmLPzJk6DEY4YeUO6U88C7ytHmjOSTDKvcXRE2
ZbHi9cdZhdO5Pm/N04GzrPsQ+jCMYCzwreSuKcGe0ly+BW8pHT4yuI/CYbOCGdieoXA0gW9O5U9d
2tT+/IpsOZ77deNdXII+Gbzewajpw+2Q102iwzW28jkC+I+9WT2bNImyYtuEnMpEGlOtmNJ3gGQr
JHOkvudvJKC4EXLN7TnBwJGgr7kGYwsjsn7L5RyJJNDktPBMcfHi/8V/QfgaOL9aVXLl2y654KvX
B7vnGtEXX5a3wW9ssc/Ya1Qcj0R85ikcO00afV3k3rk8S37XrVaKxog6BhbFb6p7CZB7oJ1Fyv3s
f6zEOwyjdcMcd5HOWlCXOorIiAbamRoTLmMRfSqxKS6V49t18SIY4T4EWhHVTaWFM85ecZFxzaq6
AoOV8tIWMp2HrLCEyq2d/LE5K+vZ9XR2EKPr/xy75plkVE+dkAnZjV4lReCpXDITbhSKkTkykkaH
fV0PxbK0OqeOsItnD5dc9zGH6cbPuGjnzQkMeMbvPhnT/s4u/MurJUrm9J7uVLHL7Xo37/HlUI5i
1ULJ4xJe+XGa1iqJ4EZ5dWUbrKFW1A5XYrwKz7/bf0OsdLQTQ6CrROj4VtBv0AKOkCGvSQtaQkcl
ZBFIe3K5Z2rT33OVzY5yhvYlL7Ctot0/LVzNvGAwlEkiCFjYaIZlN85hndG4LlpJV80CGQYwQnQk
cN6pCtCt2zqwBobZUiR/7k02+gYPq1om6n4KthAwk0W1jkxTUlKVbSf7ysH7TBBZfFX+eY0F9I24
1EddjJ42LqScHpGZGQ7lWf+7bh3rZuEghEsaQHxJG+Ph3XQLwsPqR1Fg/3TjIhRhALZR6ZiRkZ72
0yFnWV2ZanCzDwa6XtYcFWkEzwCiiyndU/q/lOIdqGnLCiMNF34qXFZQZ3v88LfZuuWtEqa4yNEG
0ToJdEB4PwQw7RtpSQaN1vQ0V2qNvYzErMXFdGko7KEpwflPpHfPQbNYYYHmjjGz5SoqSNSnGclQ
JRKyRnzvZIGqthmNAW4bj/q9Nk7GmLuSZtxKBMkyQjoToPPIFKiE3iTLROyYWCRC/KF0bDxUHVmK
XqgR+fNorW5GecyQLaBEoPJdHbcwZCEBSD5VuXrJC6lwzA3YyJOezfgQrCuGhCJLsDrUy//St619
1Q3+vooPTKIUMhp+/UncIcPZton6wJKyoyazcrVA7NR8ObM5mqAkg3NmyeXWG0QDXyFxB33DDvrh
XsBk2gaHBJkEKNejWrMpMi1pKi3/8Ot+1JQjJSplV1xn2bHeNRp1KA+1/LzF4mgfiSeRjwkCwGyx
0okVW4o2FRjeQ6vhBnrIps7AaT06mh8tOSlwSSNfl6hzf5B8XV6LN5osmnihcItZEl2iQuAK4xKz
crbrZBZo+WowOXHkbg8T2PaQj2OsK0SvXurMuIfVMLpFhszXHOX4Whsw40Bw/NCKQSfk8fv5zAzN
wR7UkyKK0A+FNACw2ICcxiojNUXghPvCLwi1bSyDFfK4wAL6D4oxTo3u3/+jobNlsO+YjfBhJGN3
lOsJt+ZfoUu63DuXrVC7LbOjwrJnimHTtJAcQ0w5jbTLHcQ6i6XWm+YUjXWk9Ytz9kIj/3o5ABQ7
g/8hgsn/i/z0UBYPJ8XxWlQ/jTU4aeRXR1ZSiEA/JAL29Rxt0pDa164mTsCwT+qjq6qF2PTwkJAa
qgSLznkWKjuQHJI1MzZz1TLDnKruKEr7YrpvI2mxlqda3kKqaaw1rXBxNQ/t5W5lSKm0kS9qorjv
3BK4OVAydd2nElA2pZ8DC+qKzOLC8bEt4Vv+uZA2KK8BMcVaQ9RFFA2qxAG5Oe1NPMsqClIcVTuN
fQvJr8ftyiE3bepmWmco1V47X+vQ4upzp8qrD1S5j5hD4x7m49y4YBhu9/mErU1b9THOWEfFMqyg
O049vT+AiBvHQZELcq1Xd+eP6aVcSwakXqhPvV5YgHftNlZdlXg2VPH2CaeIY1SbG/G9L5ykGLif
dEAcscic4oIeHQCeC1PYo3c4I9mod0o/XF7a0s37aSpkSX1/GuaaZewdzq4USZf6GHd6JfMU5UyK
q45i0KDMYi8nC5UumETVB2IO4GBoxxHtQse2zT8YsX6FFllGLou5beRxeMaLFmzgopUW11Eik5/O
WIkas3WR1pOywDxFlbpm2nc8i/wdghvd6Achia4Ym69vOeL5Ozf1cx/zX9andg2nzI3SDPB29DAX
VQ0YsNKThrUmOKixzU14BE4rRLdrnaEu6lc2BiF7sI8tIEybeye0o0GDuThcluWTMQdX7SqrOK02
8QKTrYth4Ain6ysuvoLkZJNW4HdxwcX5K5mM5ygMQCHxtdwpB5I5op1IHG/XdB6ewgwGOmUiK27D
amqkrdecZqc/88SRN+pwG9GDTop6wJtfU2CJTjXI01kaqOIAZyaswAIzNZzFKsvr9hxDKx5Ni4Wl
3Pj4t9rxsXP16C5kMnmnQQlJnidzfa4fju+XymVAm1uS/lTBuR9OC+gfLQWNOlQLEt63x+JTnPzU
FEBTc+7xwBxBKxApzbYLCZbePR0fa4vxB5hiavhP0wX3NuUahX7/L9lriIIVYHM9ID9ETS9MNOCk
tKjUm1Tvs8S6auXwpuYQje/a31NiijUEvzj6GH6mfnpFiG7d37Rqv732HlIh56K4U3QhWKr1NcjR
+VBLV3iuEb6og32vqOr3Ch2K465TO50VNQC+nJEZR0VnjbyEEq9aTDxmUuycB+nFCZeZrqv570Ha
dChBG62dUP0q9vOWawVDXefz3ncy3hy3NopK4J/sOS8is+e8e+HAWdZqpusc6HZTicjhaJD9Vx7K
eOXCZD5KOMwuwveE2YiPP0JdRDY9Ct98/HiGbyYnawfGpwChtw9r8p4134ZTTtZYskl6D/HJzD86
QJ3CXwHBnbVPt8sQLdG3T56XSUzb4wYV0EImGxUmGZoh428zToxfvb9IBlbxsHLUkPUwaM2J8EHh
uD8IJAmvRjLHab3tYzByVSRheH6XV7v7OJkvarYT2nQfWSav1l/ZbUK0UjfmLsr9RkvM1V2HKl7Q
XiFSK5cwklNhDHLSCSIKPPafopAJ8Vz5Td2Hdl0HPy7m3q9ZjGD/yilBe4/6DeDNEDXHSenFENML
LwI3VkxICQxlib5ZddVkndE+/KdG31XLMLR3riRqmVMRp2InhvdppyUmibc8xg5JKObNJBS5wYLr
785sQnjA5Dum3TOteUP03j7qlOM4EZ9xA5N3mbzNWxwIiRwvjoGUV8AfOV4N9MxgRJ98wkD2fEug
cUc7OB5pCZ1uyHV9nO43i92Aq0QL/ZJs+PPu79ZNJguaoTL3st4/Ojf26U9xYcgpWEUn+rNa+o6d
GHW8aRLJ9BOEDzU29rJIEIPF4zgdazAmo8aqSpv0HsnaA8MPln+tBw5C5+RWfHCLIV2T4C8I0WXT
HEd75X9U4AavG8sGKPorxW1yLClysDfJDDYrjg3y8eNLLhV0Q/OOiHf1FubbBNqNiaWcHFzNIM7O
Cfy9fkcUhDkQhj7FdcEekYBCBZInE2FBwLDGOgBSPmjbJ3XT6chbpgK11Asv4IO3aTbWBV4ysSVo
n316DpWHk2RkzmcjaPQJc59Fr6FeU0u08lnhxQFbyirHy9JiULQMIi65qlkNbzXHjujSGAw7KN8N
pVSGQAheTru9Xp1hrTbIPurvOqv6S2iL0no/BGCLU9WJYOTny9nID/fXQtNkv7KcgFhoj1ll5aY7
7jbTxals6/otwDOVqajRdpQ3cY2mW6pVi92ytZuq+Jt6qOaDFw7vJ3QBaP9VMLdeuiQMUdhoiU0r
IFcCLhxFS6I/OB19PuyGN1kAaNrNYUzsGhbLGrVpaWHwL09nOerDhEAqusrdroAZfNNyjrPunUmq
d4d5FGvEMIucI6c7Lk2ozZBJ3HlM7A/An7s9XVj5WdxQhZBPqODpuJk3fkXryZXwoCcq8RdCAa1C
/YCCMb1BsLqIc3PFrvfs+CCbzYyUzJmFOEnbxvqgPNSFl1Pd8M5m/N7zTivxC6Md7ErXbeRorGm8
LZzkwSxlto3QfhZwOoir6ABqPm1CYAsVzpQEnknFp9YSxEMVf/t84w3CCVx+7Z78HRb0i/5SOQfy
q60InAYdYG8kZhTKlk3qPOtwE9zSjEBlc2uvV8KrBf5MxKyGUXCFeLxyTUhoZmuvzUDyjj6RITms
IBOuM8N/bZ260EBkuAqjDZZEHr0es2h2nDwOR6UC+quVwLDiiDQkbZl95eJLDmYSmanoH8S9FWkf
BNauVHPShz+HeHpt+MzgMRbuSgV1FU4ZkY/AhNN1vR6h+Xr0gtPPtG8eVvPdWYlpHXLpIwzeoiMB
mUzbikPyKMkwgYl5NZiL/CGcP/wuytbhOSRCAdGqHCG0BjQ1XahVhkufvpXCezjCwsNr0TR2bNkn
XaU3eqhgGSXerqkZlOyaaXJE1K+4M6UCLrkCsQVnsODNTI/Y9rjg8IiJrBuh6hpIOVQIegVPcqNO
aEisHPcy1o8rBDu2AuDpSR01ql5umEDclxI1h7mNxchU6S53Qm/tjAXfLhowChE68IiNiSCd+MKi
lNaXyxURgsvDJbupYs3sT4DOfq/upwoES7DUalMU5TxIHqc7JfxG61h6Z5v28p8qv28xe7Ykv3IY
mrdTEoLSLgAHXqGdwccqMCsXhYfO0onWm8hSlw7oZbzixcB7CLnRjFjtef5mdU/+MqkWmAGijxIk
fxInXFmolknuqo522jpJpWsemxOuRv753Wgf2HrUbMPAeTHpt1CIKkW0PvDFvO5gyzYmJAs0Edqt
c77uYJw8HcLGk9Et32XdQL2nC85Q7LwkMwFYgPq8msmq91j5Xw3DoHp84Rs1IbtaOIlaU982N2Xn
rD+ujuOkUW9NnRgf9r1K+9948k6UmHUBWOAPoBX2ZhrZm9KKbNOCANyDEC2Mvmv55pzNcNpDolJC
jCJ6yn0Q3ZdreseCuJ39j4+TSWcjbW40cop2gfdABYN/97rLlyLSQHR0E5AxR5SNgHQ8Jy696Rdq
MOOW5LdPIEHbNvPCfSrpZ+7AQe3eW7Lqj90WCPuheImdR2LF+f32QJcxk+8Thcc4M/D3kYzdbGHQ
u2FvJec7OldKnIKADNGiNuTxKUA+CMznijWOYL5uE6uvtB5GhCQL1Kt3/KQ9XEiJlcDdtVAzEu82
r9zJPSTXi4cKmC/ajS1/47HxpcsonYBIVw6fZnVh71vwJEMAj6TOam3ips6QPUotAXxqt2MHYj+K
xHWR1CWxW8THX2o724psM4mxUh45kQdrmRCEJvs2MTZD+DFOm71OO9++sHpxopR2XB85zdAJX47Z
AhLl61tR9WhH4DbgnmlTyTYGxQhk7x85CZGsJ26C7AGxoS6OwsbECbhAbmnQ2m8EGiKZsA8+85vV
RJ7T7XFdB13ERKBINUy8mOIs2JdxkXVjktrATs+0fm6l9Bfv0fEGIQHnrkVqdV24dptKMLtZAcXT
gUAFOei3OJBZKbkDXZr8RDOUzzChfC1+cBh+79z5wsH/Teil/KwFFxte688vHZtC90unc14UM/8w
zR0jmtcsU288HH/EOqWwZQSeRcYwEx0MzjO+YRhdZVtkOK4qB0+yQ/u2wpO83ugxvsfrA/HDJTit
GDHs6aDSNOoz/9TdC35Sm3f9PQ1Iepsee4QCoHM38stfgwBJpkFeVeMTyEV4Q27/ekU0eC5tUAzj
EGP5cR/F1QYAonwDUbc3HMSj/LzCtQlsLmHFP0Lxm9n0Dcv3kQJzvVdvON0Grp07C//5xO8IJiRI
hO2Dd5gke5ojmlUTORvIqdQ1PP6G5ZKeC2D6UQ/HLSnORTdatE0dZCmWWjFybjJb7oq4JCDboPiw
MCidEFZ6y+oy9XtYrAuigJgFpWw9rTUokmnZ9D696F6irMsbwm4opUEi/X7x9LXWMhWnczdr58iT
7pHNCdmebwFblUfTj8E4/RYhnQszEdbke7D/Z5ecO0EVW3sQvyr75kHr+Wl4FFsWyUGJLtHABnSs
zyiMr9k7XL3BP13s7KTk13Tft5eJn/dzbYqIJJ8jObZkOz/qswqyqwrU6CdzVZyeTiZgkb/QOHuq
20Uje9pdvXX+AJWjRn49fvsrAfCdNd4PLfJP8RykMMgQDNIZw5KGu7cIcRYqjFfBRRgIa2agdjBU
0SrHvI79vcXbQjjBRZepcfkgGWBeLN1bpIpmDJIyXugciE81qUj8lj6lrPXWABtmTImJQZB+XQ+o
MqwiH9gN6Pqvf+537w5EqjHOxDCWgQg9tkkLVGo8mwVrin6e7oOLLhLnR+zIgXW0lJ8GaZGv4NHY
3GaAW1OtOBQOy5au5qLA1C6dufL8KoC/+e7ScXQDQawSJl0F5TEbAiPjV8x9QxZwwEXN73+cpbTd
cgMYTYJ1e9aHmRFWqtO+6KSa0Ac56xzAbfufmckVgnkgc6oHqLtUb+pJbX9lWhuv/pJNRksbchNU
HtfI5e1K/ldc197Y/AZGTnuIsrg4JtMUSS3+1q6cbX82wRXfzRQKUEKb6VMQG57xQ2kKqEfzdMCz
lH14SdrtVVlJjK5a9RlyXBMzq2Jx4p/UicsK7MvC2ik6PFDm7YmAY8ye1PaXtEkcPcDuPTDwB8Bn
wDgOYobTzqSTELwRQhv0hH7vxb8AGOhFoeNdmrxI0waBvFQ0XWzssVL7Qp1Lo+RcosD8LJMZHSOe
gXSRD9g0/ELX6BC1IJxwYBGG0sTMlb1sqzrEQ65PunKNpVUQBHtzPzvZkATyN7wIq4P30dj5J1ld
YqGeFH043tKqOziWYz89p8Dw15q6YEmNVlATPWHHeLUBMCIyF+on6SikbiPuRtVDiBUhAw7jHJ3Q
UnDb6G173gFeepWDXewGgAh8E0HcwInJpprU6smqfOYzvZpYIl5uPfFllign6V9+DHP35JPMAZyc
iQRBH3oSTY5csf5A241RigH3q4SWTwrWp0cAClgS6r2yz2Ffp7XWanaqL70QB2hCBAndt93FdZo8
/qTV7wCwI+EzLZUAamCey0WdMuH7p8i5f94zcpBS5dV00Nix2vsrRUf4t6ioRtVemPC53KHe2DRn
GXWry/ScsPxgUNcOKsrkJWQo5k8nK3fpOnYSGlBfJHnfuHb1HTjw20kCaYriKCBS2PuhRR98neNE
tl06k0KyPSPw+8GycwwazbkxY79xfOTWf9dG/eGTKU7rxXpMycmtyRAocdkzsNhfEQQt3UfPB8lt
2A1wn0TrVGrFxIJ6BVBSEne/8uCsASspCnNetz0e2jP6/YfMUqrO4hsjBjZiU9rB2GYJpcVHBm7h
6EocVsZOMyvKZKQMoEYhgb2562Z/8+zmBE+X2L8GPHMyE4n5e6fw+DYm8Uwtn+mbG2SZ6jzpiCLz
eLxRDskPD9fEzHW0suEWuQLHIZfID08cx4KTJ7myEClFQg76m5OBztncUHJxMmJSoKHM8wHgs0gY
7H5XGZiigbY9fZOx6wmTPq59gLEu6vv7AGanV815YSk04zxPdO13c4IwU0SbI7TMCL4YX0+eNc4c
KAiqPI28gBPiU+e8u7CKJkqt5r6j8Q+rXQ+PP5TO7GeSXnHhAGPqMta2ue5GRk+S3oUSBCN6Ccav
oaRJZieuzrU2Mm+FJr4d2YwptPS33Z5UaW5wELciaJLuVlffA7fcMTKrnLW01yCQxmGU9o1zogTQ
tj56YSMAt7gu6psXflXKPu21N0yPa60q2iYDg0K5ZHkMucSpZxCY7KnnoD2Ke7ampUJ96wsnl/AA
UNVblI5i3svG/FCm9OeMUyzyzDFdmPsnxionijqQK0u1SBCuuW07bRqLHFSr5Ih8os0eQ9Plfzna
VJc1QKEi86NmCi8vW4LDjU+7puGxqocioRnYW6tP3UlBEd/adjpDuwywVt806EwdavsVGcWepTuj
uxr2yS+HGxwvmkzoXxD7VgMJf32OUSqbbmv453viAsmovAz+ggBlJ+2zfFPtI/Qnh331TVMr9EO8
htUqV1mxaiUcOfhfCVTHIKF4inbmUnKOKgMjv9XwqybhjsWJ5xFdfscd43Yp9ln+/MqhvEhtVGt9
nKuYsM9+ozO0AyLNwM2n+OkfaVnMJQIKjbJsGJTLyDbA6lW+mo2Bxm7eCNjgLZ/IqhnZ4xTUnvlF
kdjkF3SDgXIbLxroenXDt6S1YWBqWc9ekA3dUCMzM+RgQIFep9ZyL+YiaoB+HP+Gjzwx2LuY3no/
cLri1pOm69JmcnEbgkCr1v6n2zttqzV1OTrcnQYhoIy6d5nz2Wyca8RK9tcyjeZM5AfTFOQl1aRj
BaWoqVTHOTgWUZnM+Vfnvv2PuAouHux1z1xgMOwCPPCEEd9uR8l1Y66n950rtKl9/6CdLpqjm90t
dTa8qUGGBprFwbzeUDgpGVl0r6W3UjRPmZWTtZ5qEWDhABKKau1YtwId0x4CG3Bkcnf1RsjU/Utc
qBsqOGOBL1a2wxlJ9RBhIMqQv8QUBHKxjRcM9mxCidELsy2qhv9+EbHZ9A5PgxfwL1B8NZkdGP3o
DP2jnWB4TLzga/+7Tdh2dChtslgLhDhUXoRGNvumaaZzaJvkDv1hEBg+xfOJ2F3lzDb2ecagDmyj
BDzqYH81cN2FA5utmIQbbKmUfI0TX29RFkYeuIiZK+bo6swv/MG4MDxUHav7PHZb2Cw3ldOe9ni0
B5PyQfpsPzRMo3H3VTSYw6ac1eNyW7vQKujQFOfS0BVPsz9TKi0Chk2rGxkS/wvX+G9LY3DCtnSj
m21V+PPFg12prRkfWIhhU2iPG06KgJxf+NqQ0sDZ2960+vuCbronGXxVljy1e4kdjbUvLIogeHrV
Gb5TGH0NewWyZTitalGJMZlE5qdNkx0i6XEQ6NFDvKM45f5d/SdvyEnKuMfq9jHDgqbbnbY9EfQj
QYKvnvhZikctcI461YBRD0wc8ke3E0CAFGSGKsid8d8rI4vgPQmUyFJTklTdzB/nEUFeGgg1tmFO
Up4ra4+Mv/Awp1oYH90VEipRPCeQUedYjU/6ctZ7CzigegAaCf94qoAGh9Zft0bf9RgJfLiNg76R
Rm3/ak5FXIQSp2sZKm2zeQmPbG583hOyC6Y6/EvvMXLqDD3TyLkyOZ0PmpOrwzkpYbH4DLKotXAP
/6OV5VXt0p+M/7xB6eVdxN2pGJipTikkQ5jTmxq9CVTbOlrhDI0M9MUlvEQNaRw9DF6v4uXPPPS1
bDe5UBmwUsfV00r7Aam6nCIInaZV4b/qvD2C2/AjYPgorvS6g+WezbNan0OTHAqAMLeEM93ay9l7
X0vbDHA5Asro4Ni0wxJD1qjOWlP88xwwg1rQqLecDsF74fHfKG0oK3WLpklKeznS9lr+gLMLd6AN
R143lY+CO03QLfbOWZlzhz2Qzz/rKlplDalo4VW16VDXVJW86mbl9Uu8sJKhyiIrc1XmS8m6bqlM
pKhxVIwH2XJn7jfIs2/20LlwdeRTV6C1krNeLcktAMKXj/s5U2IxdiCm5zIhBMAhExaiKEk8mwxq
CQqiwVNGJwHxrgVOB6JUgvhze7dCyS5Hl00WMBnlfBOLQjUj+YAkexX/q2X9M5K8/dy0aXnWlfFP
+3w9cizHKiTNqy/oDnFcix+360jqeWupGhyjZJrrj2i7JBrfHvooV7no3uIQLKg448F0yBFKcTHk
a7jmtywDpiiX+d6upqKZ59MxxdqwC1lwt7H44m+DXFFGa6eJ2tTnM9+eKuGq+yNBXZwi5jCj5azO
rhci18Z0+eWBUlAyy34bW/3etMeP5AdvOT5usN0/XvcL2NVeFFRHUnEKp6LSvqpMnEApOW1ea4fr
rD1NlTFp0gp6JJyLw7qKgiqUCDXwouxuYytDw9H6If2qmLHbBDdsBuo81j7fTR/Mmpi+dbPIA5Oe
7PXeCEMod37C98Tb+8OJiL+v4BIyZGqav976fsOmyY3lXviHWnQrembciLd9WkKzQL2r4jLx0zof
yxLkEtndSf2mhPzfuH1YrFCVAxQ9fldoXAAIckIXJ4HcrbDmuMaIlJwqkrkhTgC/ER3DWuymQaGC
qFZeE2gVDF/8w9AfYEtb7a9OGSiWyGQZlAUmY4oUTyTvZ4tGM/Bb8reBMWeedUEg2aG/RDgLB34Q
ak5nq6E1mhdJ/tMtjZUcKGW4WySiuoipF/Wvn2t/W2pI7i7p+/gvzjEYjRNFbeCTsebsB9KnjDzx
Gh0CqDpHzH/cNKurPAmCY4G/JBpJQ4fQ0UsJEq6RusU0PDWyTFMQRzT4gdVkc7e3l/pIPXPlzemm
k8sSl51tTDEDGQxEER89IVqEU0NU3VbM4fUNd1+B9c7pJ4jcUdvOXovg3mbuPsHHjROcuv1ch32V
vyz4j3pbxpth74Le8aAa1dNz1QOJCzNQ47SSpQB07SdlIE3wCPE9dTsNhBZp31DHffnucVBwviTW
8ZrVQI4Qh5eV+G1Qil9VO+Y7MeEBKSQGhO+3gSBIk5n83AbFIJFQ+ZGd6q7ltyLN2HGAnI6NYY2P
RXDseijgYa4yJlTjd+Fns2LSnDgCdZHPRToq3+TQpxevQ1CkJIUGmSqLNISJ2+IDK4In7h2wRtAO
gVaOZjftTQ/Ja7uK9ccpF0/x9u2AlXscgzoMRq5BC3z2GEZFyN0ovO/yLIAAKm+naCrtBNWQmpco
CSQOTWN00Ij/F2SxuAph6uSy+uuWGVknDyWocNBQQJLwB+r/OdDn6KUDrgyk98c3HJ1A05T0tuFS
maxz+r0eMhRCj1ugsaaIOHm6qsHTHTWdtw4/iDBVsCIndD9hhe6LCF8JjZrXZG3XlVnKr2Pu+Dyl
xCvkvl8YeFFGDyav7RvWkYSAp63qWWkxsN/D3YZUrGBpaFyKZsel8Z09fUnGgICPKp9CewShQKqJ
e7LtmL8m+V3G8Q6h7h5AyjGv9PMluBEGJ//B+FPSFu4VFG6c/aDiapRVLI6tCLI3JFTH7nQkahBo
M7aXnsxmXib/WmSYqw4QwBr4/gS5kPimapdRbmboDdeMRz376hAeR0tHxHlO8hnQxAhsM+828381
cX+YwgDQut0UF/hVYSpML1+Phacq+t2WZxhbV2t54jr4nRLebyUJcDYgISZ+0nweoeJRUhciwEwT
Ys5/HSeSHQmJA0ScgZ3Q9rCiZan1HhDC8sDdGgD+b7CBpL4qf9YscRQPxDdHgaEY7KXz409Rrz9D
blSZVh2mE46id32bi9MD4A/PYEcCuPa87J2kak48iBCNDlb5ECCPLoW9pkuZQZjkGyv0PejUt/XW
oXC+tCzIbnMez3dGLlu8ndSbTeyV5OzGiKHE8EDp4sWj0qtDjuoFp6mlPLqHvM0cplOVf55mpOe9
3urNudNpFyF5iDAYCQLQoPD20yy7qTvW0PzlWA/icfffxgI3qaIqEMjjeQThol5BMEG+kYyisKZY
6NQfeAA8lgtgH+R/68MN8VWzys0NF+28MCoLuDS25Jegfu3q5rsIyTzKwTsE0vC03polZpabtR4z
5kJkx6HklJXnX7b5fdRhHCPE4go8tU0OsNw/v6Ndaw8Pn99n2LminTVZEDpjAZ4At4+crmvT1DWb
u8xTCCldisv/S4ecS78BkMQGhOBnUiWxA2SIm1rKHBGs3NnLk0q7IzwF7bGxQb2GK2S6mOAzWxTa
w5hCLMbeKi1U0pdlq5YkyPtQ8rV+QXRl+6Ba2Km+ycT/soJkenbTU5psC76srwhP2816eZRF+Ym7
7lsKLSUcm0AdDe8s/J3qFVTAGNL2xMxG5U29xd13BCsRdD/8iQUoPPsIzBwW2RtavWpjY5MzheqF
ZU884+DgWKbUj3c46rg7rW6ZFajOx+eOwp2LiFSIjpk4pwAWHXwDyBNreV0GoIRZs+efafPRqnNq
rOVeo8OE3YC6BSTE6tuapcdqjtm5vVCDvgVCr8rL6hODWmlducCU3MqgvWzSyXZaJDPnCnnSmKk2
69f/lOgRJV1DTw+v8uPTRWcMe3cecvBZAx14P4HEw3z574GSlQY2aOmkFPmr/07gXbYiH50lbo7v
4++5tyJHM7D6gBHYBrBGQPQr0phS1ssazBGxrfLoLhCvnJ9LQGQR6pKFwt2pcF8BukoEVQ0CC7Pk
DBLx28+TM+y6Yx76XWgSjhNi2XkJpYDwSdF0J2svfm6ShnDFE2rf3oNfJAk/WOdVeuxPOeOuTh6m
Owg3/CeexTzR8oiCQkpZFxa4O3dPiOACV8nCQAByIttb7DytFltpjjQHvmkYd40yg6K5XuelK6TT
OzXxOeIejhpxylcoXew+pA0icLjCPjGF9Pj4JifBKJdvyKgco0hIed+XO+cn1EXsQjiGY0xC3lEn
fRgy0RSreTXaPj+HJ9FHHlfJl4Qkl5ApAChmGCVhPC985QPTfqFl5+0qmn5dQljY2/4jDCHx/1eG
mDgAHt0WnwnrqH9O0s5UTcY4FaRSc59UqQyohHPPOl6myxEDtQjE/u/9KB7LY20+aLNq7xMmPTlp
54moCksl6SRuVrAYFduliw+2SzgJOkWlJpz75+loOF1rZL9655Xfwj3LZnraQ46TIU9FGNDt8o7L
kJzakdXr3Vvnb6UMYAQyqmK/LI7lI/gTogUcea4Vb3YXKCmb746NU/Rkp+sj0Ws+EKl64Yc3KX+k
q9bmDuSEQoAfxJmh7PjBlMQzfXWd9LBuZUJqwwt2V2m9JN2wKjUXKJDajYLieLtiZZrjred5cBAd
AVjjCq8E14DnayS8IIiCxwWkDvYm/oZixzJ2vhQX5loBW1EjhdnnkqZjZbhZgFKLO0R3Eb69tdZK
GoEWBKg30KrkJufzRWXdAOu1MrR/L+bBILNAYlUIo9t9rtaiYbtO+VACsufFma6/oWzaXVoddCru
t+ipgry26jrwAjJWapA7of9S3iyeoCA2G4O3R8FI17wTdw4OT1ZwHSJNB9cdBe3fbQgGvzYVy/bN
XA9QvDpStTYNHeNPT0DyztjhQV+Fo1BRx3ddrP3txhgDjAOyhheZ+24yXRokcMWuC0LwDSTt64Y9
0xZkdoOyxlyeFUstu981ajSBDcSZjBRfN5xHeADLY/AxS+8iZAR1sj8VvsOFjT3pswaa0Ta/twky
2U9fvG8CPG4E2KERS2tVDzMhRuywhDc6UMms6RNjUNokEmapFTxJr5eAMR88lWfvJZ0OEvtVfnBC
TtBlZH9/3dsP10D4VsYt5k5/6Xvqa64cbRmj1sw90E0LxtSzpW7OCcq+p7kRXv/xY21sNdN5gsAf
Fh2nefu1oVZ62wp5nJhlDmgtviandVGq5ES7wozlkb/KQT9K2CfwyKgqK7SN1zTN3jNv75udm2Dx
HyqEq6yEzeIS2623ZG4Cen3+ib/GDKnWC9Vwne1NhlUZDAiZs77SIESNviZomAygtJOrUcPhkZZ3
w064F8e9sL5zBwWFykzGkO71XWlC/yNrl3aN5GU9O25R4+cFCTj73Tka+7Ce5nKqQq8Uub39V3pd
LZ/PQt9DHjQ5WrmIVgd+DzEFjdmIYD4d+mJv0aHw1onZ3frwqu3gLYXW3NDJ2W3H8x5IzRmx2+px
FHiIWFJIwsGZg7N7LFqvcFNsHJbje22vOzJ9714ZF263PkYjNuZBivaUsBwL6WAWTLLsCgOjPkvk
eNe4lwBClFRL6JXPG3UWThq8FywUb4E2gKQcSuOX8K0DV+LWFf2hFMmxoQA1R6IpL2N1GnnJsrT8
89ZGDeascsqf996FKHWJ/LqyOKYgbCr5vPrq5i0X6orLJryZBFJhdLffDUX+bEBYkQsfWhvCPyBY
xZC9dman+golMW7ZSejz1GdXjRTBWAUQCTNEOIA4ex650A/lU9cXKzfq66lcQ//JRKBsJQAz37O+
y2ccO979V+ShSi9d9mPq+W7yBt5pnPWtDc7XEOwEwUAeIR2mOuGRr3NJx7XjNTN/yGxI+edK/Ezc
9zQ2ruFuzIqGK89K5blFR6fg/RDZy0kCtLMojgWlgkFiM8zrWhB9kgnllDoO9kYaeXp3nWwMze1v
46z3acgOh+Jof+3FOsXVQTtYeHG/CFHWK6YeqOBW7cgplmAvzMEUS0XXWZyNIdNqmCi71s128L23
VM7H8hcZVuNU6O36/fZOIEfx0XTyJ8EvANBWCQcN/kWa/OUXVsuZj3UUwoBE4Fw2SNtIQrCiDmNl
ACebJgeiSkHWmJaqjJYlTDWG8/irTxJUXG2wF0vEvjiQj+gYiNQgzeAMYfViScFZHCKXlXqqI5Ij
9Cm0wF9jOpV3FnRoZajPJeZWQUOCCg2aijMUoIDr+yvWTPzw9YW8bTA3GuGmGSoEFLBGeBYcdOl7
nlqtb1k7iOuoHDxaOd8U1FNSN7mAR0ZeFSVeYWQ5EIaWbQk0/JJygtByfKuVq0AIQUHiszY2OCkA
DYr3kCv49b/ItZxSfpphCQ6UI0PLLPrQFuzVLFeD2XdYXbghlTelBVeSDnm2HocLqPH6BaknBHKK
0nyw/nfKos427wKh+f1NN1bSvfpmMr8q6FSak43TM/9CWXMa4pyZGkwERXvJyp60y2ndApplwCAb
lZbTkBcDAX7wSERloq6EmHrU1q2fSxC+4Y9oOAEW65PiC6+0uDEq4ywqrXUSBLKoyeqDCTffSQHP
YcVFnz/F1m+M3JlVfx9Uhkj14hzk+HjEMgxutkMq1epxlzqF0D+XgB7zyMzw3PjWouWVxQfPe1pY
cBC/mDlM/+mi95UWnF/OPzG7EXts92GUCtHwnw5LEMi2CY+K2sLGTLNrLSPUSfZP7Obz5h/aF8cP
06tvlqRdW5a7mOn3uv1vvKtcQmCrGKloXeX4wJOxxRzRcVfAJvpw63JMBisxxO3Od4ciFinBnd4I
mG9c1T0I1USdNQ8FP7pxcErie3SNSTWOVxmq30mK5iZyLnjmixve8HFWv8SOMTjvlj4pRhZm7hVZ
WfpNOxMt1Pnh83ae6DwiXt7HTGjL/DglVFZzE8itaTYoX/3xcF2baqneP+E/d1GNAPEVBIbm2OrD
sSVRYtajB9z3PZFNMPQOb1brhjox6ZXyNWZDk8uDpyRLha3pE27Qh4tJiQ2cpCMQAUo9II9RcmMX
Z/+LqiG5WVD9d1/REehzosA7QdCUrQZeAO4SEEn7dVy3D5gVTWE3IDEmD5/pciZZ8zJcS9scrZTZ
lxlDfl6AoWlAIXRqMc7GY0jOTtuDbG/2GDh8YGqu97VSFo8WsKIGxxNggRMKMS4zrlR6FSWGkJ/d
iD+6CTX2wnPTQziAhEFFQ/B6vBHyep+S+3PcfZALFwlH4pq0R3b5KIlPE+0imVIwQ4GLYqOGLLnR
1QxdKoLRr0svCKkOWaQnF1hG2CMHzAFgQGTLG3h7gyDJo6aNUMO7hjOX4KH+EwiMFg7DqMvXo5vW
xM++hTfTfLXQ8zq24UhbPtx2VrP+oy8ON4HkPHiNv+p4zXOiE2Jl4Jy1kU3z3ptosGv0prGBoOqR
JTnJB1W+TM3ridlenuBvX5l8MZ56VBWD4OfPN+NfLAdFSHt9d1+detfvP263FNsv60+kQe197Exn
anNw1tg48UibV+URu8waB6lo8EvcsI6CPQPwpi8wqgspnAhoan5r4W9HWIuXavljvv1PVsbz8iH4
anr6/dlmLAKEy010WMGrFh6GvWjsCpdOaQQlmwBXa/rrYjvzBF6fk+IAeGXh9GCRw/hGeLMNWSI6
TRlE31b6uuWrKguB153JIJk7DVjmJlUf5GnJMRfiTRWfz0ErmlIFVmqdpyfEAxmu/RHIfhd4HOse
vvhfGGvl9nZe41/2kxxiRVB8toLIS+AFMYtzlBeWsr0LmjRelk3Ud/qE2dxRi4eFgN7wwlenlPAt
OTDagluM543NT5MEeNzFjDYyywTBwFfbFSIdd5Tf/mtmEwOYGCcuA0bSnA1Apeu9Iz0u8YA+Sag8
C7NIvv32Yvnzgy7X9jBebAnhIXYEMECMDx1Q0aKpC5lw96uP7YWDklraFAa3Ysy0S2fCUe2kWPDY
gnO4OzL5FvrzD/SxrBEEZwGbvxVYo2ab9DF+AfciWiWaDa9oVTLII50ifSyuApt0htcM5p0zmuKm
HtuzqLzt8yDIoaUAarFjrLRpyXr9iv+dXBUcT4jEOwjcuBUoAe8F3D8CIBIX5eBor1x+M5aF88gp
OOpJfG19qOnh5Vc6tNhZHQaU1dnVCd6WJzexI7Tl0zLOFTItdL68boX365qBmrNg95XqmjJzCbYx
agbPpCpHGDrH8Q/pXs8GP7GJfXm0ywqrll/eM+ldJk2xTyexGPh4FIilYufMGO1BiZF0ptBMlC0w
9k/RidwDJWvfgIAkUL0BtUNGRDhdQXV1hRKyqmlADxPkwM/Cpk/RyJUV5l687lWO7gDwaxj5YL+X
Ic+7k1JaNarg3Zi4QV2GYWHy/siyLRA3RIDk5yk7AGY8E0qwDbLZSf7/ENLvohxV/rQ4vADtKpfA
gq/3VGVQInBRX4pxCGCoqqVVkGCo9mJBtrfGb2OcVkAB4puw3RfRgLvgE587QEqBwoMEU++zWRmU
HmGFn6sbqw5ZG6g5X/ohvVC0lsLRJBwAqcZQgvmsIrBD3aUax0D35eJxKYer915F7LwPJx8KdhRP
t6mie9rd7iMysMrL2Z4Clxc6Qu4iEpdzxV+NaoSOl6DE1nJaMPLYj7Pok/oY8eT5d6MvW3G0Y/Yu
3980fwLUM9y1hX2zFxFpCWad3QawO2D85OnFy1NbcaWVYVzOTRlgx4P/+9Ty18SN68chzDj4t1d6
qOEVE9BKixZ3ufXQGA0BeOpFqSyT6Hti//FVDo/uCKgFuOcwa9407vNusWW3ToDpvC7Q/AJ87GZV
JCi+APHrJtIJ5XsiZzcOy11BwgqN53bKMBoYjwL/RKyDx+5WNxSg43DfRZUJByotSDMmP8wIl8OV
phSNYu3OayYTXhDWbBaMf/U5xUeB5ZzXk/InzY5GDq6YXQMAx+Ita7Es56t7akFMdDAyxf1MUEjf
5uwduNFNtW0hSaJ/rITRHkLHhpiYEvYeUkEc4i5I8+cXaumE12G8FE0ItukHAkEEJUwE9VLVOKoX
CgAvR6EhLVblnKu0U7yVhxjliG7Mms52ahenVlSvOvx9UNTdiHwCQj4CojzaZOFQgOaE1A18CV5Q
ncArhlyi7VaflQxMHUTYRNtrpgmcH5fe/XFGTCxvmltU5s+LqNjeWuz1ybYVxMasSlAmRqlEDTMx
nBIJkeS82gDxmPaoARCnd1C417GaLN1UcU5S3yUI3uIRKECkcLqGQh8uoFcAaPFxKBqy04tRdWqP
xihpcgA6YvBNf7uWvAywG7G8EA1DMjqO20tqOkEOf4kozU0/Q+hkNlc2GsOsCx1EmRTR1oiuP6Ao
UQpc+fMntm3wQGOatW13b0VnRx3oQIPgbXOiWoZtUSQNWK9YCUesVGeBlj50Fo6SYUz4jh0RuLfV
CLeGH2l/GGpz4kT82CtHJD9ntNAeKBI/EhUuTExVvGEPUAZcgiOk4HdQX7RvXsvQCSqDUF4dNEiU
Fe65gRbNzhTSsE1KrWW8doR/NuXCPFpnp6EsGnpsFdmKWn//XKOFASKEVhcyvXAe9oEEOoBgWva+
ib4bmZqH00qhOGYZKJNDLRsnAsYf1ETtfUFLLDAUEe+H4gc4OZoH8/akoMVsqC2FB/pwX9sh5rA5
0Zcb7KmBw+cn15vdpRfmlqn/8QJQC/CnDdFMokAwu+pawuhD4NdMfXi8jNaTgDMFfHUc6+glDfv/
wyKZJ7X93BL3GQCauFn9Pt7EiejpkPgHtZNBrm6n+beoMwcbP3QeUBYVboSRbjSr2XIJVheCgwaS
fCZ8aiVtmetbo1/4R1zah2Z+AjmW75zzZXN3JT7PrrfWcXGD5d99Fm6u4eQzQt6pKRQ+Lb2lRU11
1VKsfmQvNUGQzk9+/RTOnziLzGD8xWrypnf6s+d8R2dHaz8oM8hWhQlRz/ZLhQFxH4SVVHXCGu5W
A1ml0GJYSI0evXLEQo0snihJJ/S9zpjFlk0egZFJ6foFGIk1mEl5djfHUYJ7EhWzirGDuexFb9RW
sqwoyiJipIWcCQ5U/DO+R68T3sQvIt2yOqlGqFA2RGBdLGD0dJkJelwbUZgT8uZl8+MWTrVHlbPZ
Zu3ta52nRuegn+Gwi3RR/87a9+qgSkBwMdM/AoQPSw+BHGbqsd6qJT6K8bDUa6bI2Nupse3OFXsG
CuEl1/JUIlncziZegUjRGWnKlMNVa0AchpeCVi/IltFOaa5J25c5NJ/afnJAH3vXABqqpd/LlSLA
F4UPgpbAP/vYuzXBRpEqBD4a20JJL5Ngr2nedvRtwfL5z91oleQB/Mltqg5qpMV76IlpD5KVI1za
UGSm6y5//O9qRY9p1xOZQb+Z8NTPM6ECdpcUmI+Kq8In4wMRI7kaTckQJ1IYDOn76Q2jLOBTotOv
foUrugzSdfHn1FGHOV+UbEOsEkTp0aFl83XYuavauQFlUAlrDPILSorGA+T8smSz81rlJq1Gs4+V
OUGToUN+zTniDTTPjbEXR1a0VJQu7c2z7ID1RRUyd3wxbahN9vgRC+C/LIueKwtUV4lpXstRurU7
bhtmFcUCSGlpotAMhcEdQ4u/xa87HE1zkAbHtcMUvGoIwuLMjIUJDMb7wGpDADXssjViA9ojKFmK
UDbuzktTgqhnYKr/BArEsFbt534888QcI0LzbnHgru3Uxpd0qpRYQI3MAwItijEu0UKwH2REUtLf
+0u66s6KU72Vgbg9Q90HNQIX23QPdnD6tahyJ8LxZhVZO2A5NlC/bT/okImZDbv8AkA2ocNS+s+v
r1nyL768BXsbnh2EbK4GDS1maX+PpLmynIZXRWyU/y2r4RDsyAUg2sXV7Eo+He3+a79yHkZAdj6N
+05FrJ8gOLfKZNViZ175MHtHSlp7XnkQyoHZjoLB/QNofW+Pq5lpPX7AIdF7hW6JvdQANbt3581K
V1UnOg3a98JJ8C4IFoiqGW2hrpUupKuuYJ9xKAqbEPUh4kvDd89UijeVUCR2BYgVie/8bFt4ZWFU
Ak1UgGzFFbSi1jk2Kx864OblTEJUY8tNoVrRoZhKzUtOQywlSPI/CUzL/4FFWiw0+DCxDCrdWmMi
acTUYq7+qxGXbdR+xOGKMzYQPGJbMJqAMl0ttqsfItWmrXxYNXABS1cLdpIaAYcYpY0iBUO60F9n
1IDyQFPjekZXYb766Kqs1nb/WFrb65o1HxEAKkiVEK1VdGGfU5/vCnQMoFQv94CBkWB/qZGzxwM0
ZRwqb7hl6+xM0ksmGfT6S1rlzUPf4Wlp32N3XiU51X2DUefYSkeATvuPXkoojWhxV+eZnqsCobsB
I0oxKC4S1xarsiat6TaE3rj0KlTpbUegRWT6rpwT5KjPSsIWL1f4Nazqd88boRzvLDEY9kaqz1g6
7aP0Z3zWXjltpHq3+UHRdZVsdVMJor19Nf4dqk6nXLfsKtWQgrlIeKeSuP1oOPM9qqYk18ViZ4mf
kSgMAM2H9Xmzylk4y1ACNpdT3jcOCV7N2P7zInDzw9XK+OjWNXleqdPyDrdtCbWq6UyqFQfPkZvy
OAFzbF2fT1PSM4G+kxorR/4eoihys0Lmug4Uz8XaeT5/Gm4KC7TsOGH05g6J/J9PcGQmSiFiFt07
Vw2ih/mDzTJio7cidwo+LLUaEXDNilTstIoO3/7JDjBu5ceWg9mDSwPgX367FvkBRVIcOc5IlhHy
VxqM+yJ2k1JV7nsR0MinJNLPqMh75Fst5N+F/04Ablwi+xWRJSaIxBiLn0SiU1EUYy/tDD84/KXn
eW+4t3tPpXBXEluGXAJyPB0MyKJAf35zB432fLKSAie+imWGzm7BO4381Im1Bw/SV3a6B6ZWw8ra
R043FtxUK9/XBXocZ8f0p8Al0nNHQd0rAMfGjqQzlmHtEu9me1xcewfrD+NytWDUM2/hZd8ISc9e
INueZoyqU9Nh6mswjdN8KcIfI0qSzoWTRdvJ9bM2iM3y7e2eMZMcxXhfmBxV5P/uvOEmEYULY8j3
1KIqypYe915oEVdzepyU8CVauuHFnyodQGEwXfXdv3KqBOTTwvq+MpRxXSY0/+ZZJCk4w+tDDC+l
azcHwBrp3z+oXIMvqvHomMabR398IEFpTIGKQ45s1vt4U9kfbOicaA1b2FvsbSZeHlPXIB8xl3Is
Nu/mqKz5ndqA9D8hivdwA9h+hnbdZhkykPujpnrOIrooNIDXYUu99Jm0f7r30mXn4+T8RT38ZjjT
Uzqqm7Uo9XLLat0/PU8CEk1ocH+LjQOwXvLvgBFDCoEhugoW28DlyQE/r80t4Owje/hG5T3DouOG
7pCcaAeDqEX1Lgbcr2kMYDCf9JvgAROPJCNLSenQnyU43yXXaErGtb8T/5DR+KthQmDR2ygFrxQO
LpZOk7GOJAhtcRXYRCsJ2iF8bn5L4R7dkT5Wz692878K0d3DsiRUgYjwXShi+b3tVA4BBOstKEwA
QWVK/4c8GLIfpNXIf9XLQlxKdJotToLgBsc+0uauWEROpUZvvoJK1IsuaNm8FHgemF+KCWR+eQgR
G6LaJlwSwWUZQqowSum15dnTULlST2222qsDoQB9ijnyP2cuVYZWobGWz+y4JVYZXq2vdMoVpSW0
371suv6BkjiSIu8mCnyCNjZqVkitzRwL/+h3AgvJvZl8bjkqMviL8r9tplTH2J36bqr5uPUqhEWG
XqBNJ406xOP6wskvNbRkNOywHf2+BAQGn9144daUxncOvTyTTt6308+t0Cm0eeU1EU2GnAy7fMUP
NqxqaSxm5kHuyLG11hx1btzK5AYc50CBhJcR3JtIShKfPhLh5rl8PZW2uq01vinpUm7tyGzSo45M
lSLFs4ZtkxlF6YRIKzzevFWxLaqB7kcoM4r0k6T9juncN1DXhgvCuj7Hc/B8xPBd8a9lvWoLPd0X
IuWRdhSxapaI5Ne/5zemo3V6Nv4vosdnGNsEeOEnJACSxAgfnvThVnQ1dQItE4FrdyY9NNeDRhio
BSRLWonAYSpEFyMyx1Z0bNMXRmjdoAlZ3cFNKE/CviM7FG0o0DPHl4AOmZcIgkgSVwU4N2h9xUoG
9qJouVkKGft6t0yMomXOLLIR1j6P0zkLBSQLu7hYZkux//E16pTVDcNd5Xo/TH0wIO8/FT2V/R3F
qhQ8kdGwBU8a9QAT1RpmInK4hL4oMOKAstR1KQ6IqIzX7AkasOVLEsX7njGdgmCupStN+hh6Q64y
97j+VZ1SZZQwK6DWbVfLnAQsSkVHs58aET06xGI35qQBhvmCT42Bfg7vapIhvScmobhyNzhJi4/f
ONT08WTcPH+6lwSahteXTCVl0Q2+Qg9R0FrahwOV/h2zUtn3EDxR+qG39NnkMdfIKLiWVndoSXZk
4ZngXxgyAP43XMp1ZJvBpKqDdTBRseUfHGNOQjnPJf6OTTWkmvj7jD9lsTMMX6PJAdhnv4v0akI6
WfCKIppwq/K1tt1mXhH+v2lXBbWQD2l7Yhk7qD9ZoHvzk9CL9wXU6+1XSmu/Yl3NKn1WQ+G4pUbx
jzQRml2vPRcosSd8NoHQjNJHpMkw8aaFnGp2ZNWPpTxOOhCVbONb7QckK/nIQmPCbBCJyZRnGJi4
Ew8BjkeaTiHpJkVWyL9J+fQ/Zh+kQzan6BRa/+C2ZotS2L/Ym2ugfDtd/Y5BSPHijxryPcx2+wcr
j+hbgn+4emYr/K0v5XiiT6cqdN0d4yZaMNZsb90OpHQKKKPzoEkCQgf+1t44mnNKBeZhsmwTKDaa
Pqb+4HBkPoXeWUqQhOFHpha0hlArcVOAvWKYSHNctB0u93dvGjPKb1pelGBQAhEs7gIaeXwc44XN
UcknLNcrmX8GYFjrY03g3yI4zRoAEXIvbs6qsrlPpfQtQGqK7OBquJrIfV4Gyj3AvTSTMLhaJg/v
ZiML9uNQ7TvrdBIMMp1jZXjPMVZNvvAAc+0cZlLCqJ0YjnqvYhLnI8SpVa73+jYan0lz5E5eOT7E
mufb9+CTQFZVnmFa/Fm2qGarGAT4GrlQi+euhf5eoLGyp4gDWKCLSbXOwo6oYtkiIehz/99WtFXa
etb4TD+wXinw8M4+qVqcg56kZHq3a8mo3GZFt57lIx2LUYBvAZflvNu7RI0uyAR0d3LYKtA5EY3t
RnloRzc5vub4BfTCs94e4QSVxV/17bKJp97FOqRo/8QP2452gUcTJ1WJ5O31qePpCkZNQU4D+nzT
9nXlkxjkIYm+ebsYs+pm/twSAPIUIgcohYNdiBCVZURtHDaHzRF8N4Fq/8n9a7hdmd9hPYI6FdIi
LpJeh8HYHXj3behQSAXMPvC4hAPv5SvE8QHnxwKtD5bRFDJD0EMbbE1sh1MOZb/Bc0giEROHSQAI
bx0RbthI6Iq/zCmFclFNUa6B0yi1moRLmuv3QR9d8vP7wyTpl4DrAJmAkavXKa7IG9WCzTMAwo3Z
z3NJJH0NuGkGeQi/oR6BJkrA/wgz1Si9ZJFrdCrOVfI21mMEJlwvwvORGeZSIdObhXLcZ8+MOL3B
a9bkyGgPDlYkDyQhCcN3gS6hRFbbzMokC3+awyCydur8ly3F+YPmN8WiLdr0pcGgzFcOaIlrTrCc
J5lGEqHVsyP7zIu301rpXYlYfkWLuSA4Sz7kV14IWtIQHeYh8LbzuUJQjYQq/ERgTeM3zGcJy0SD
snQOWWZ0PizpFVm+HxSK6rI3MzfO811ki/q2PGw+8Edjj4hoVHT0rCWxlA+ZhTkulNeerYp2smkH
KXcnUyk5LF8J3yemlAkp7I7T+vLosuas1VqRYEj3DabKk6UoaC1lNkCl0BV3isfxqoiNTUZ9Phvv
GMpfI1HBDXrlMmK9lp1VrwtRSdbylRen9I4bKRar4VzlxiydNpz4x4Vt9Qb5okYzisZRB7HZaDnL
+TCHk8MDBhHo5IbnRv2EaSILAow2A57vDrLEexK5oAQGZCgHK67dvnmcURI0AfoA0wiSYpOZL251
DX9c2/mswDYcNti5mZzfQsPBP+EN0kJm8J7TSruPHle34b+o4Fcl6cvMCkwOzsnJmEbBCvVrWa49
hUtUmo0sU6X11frC/HZQ7LO3X2nDK6a4aXLbfy5QEb4PpLJ/WAIjkmNXniZuSE+muJseXANVTx+t
SyVOkMTP672AIO0lfczwdON8ntUn26eM6uDc1Sd2V9L6xdphmtIbzdIX+UXTy1GV+hi6twLd8ICt
vVbbbYLYUqG34AuPxAukz2GtqZPxd2Eb1k+FDAICOnzDMSefcEPUB1TLO/TkB8xPXdIdmUK3mEfB
lmrJrejL7k1eZwlD8XBNfigNZIHzVtxw20RmKnY1Eolwb9SpSqnjXodCWg3+yWTNuNexlrqRCnCM
eJpfj9Y886kftLMFXCtxdAv2zW1agr6Z6ENNGaHT1mYNC5q2/vc1X7HHrZdZ0rjcOAicetE98pmL
TxHFJdKrXngYkG8Jn8VhEUHjvv1JXivVFB3q5iJ+Oqhg6Ct5SEy4i8bza2E5bLyo7+Or4F3M7RG5
+UDtX+zquXSNK8LUquiDuI9Tj+mH5Sd4D5UMkOrtjSWe79JJIf2LyQczZIfQMdfe/OR9P0dhcTzY
qzpiywf+tSQvMjzrYYIfySDTsT6WNPX/1HCOK7GjgvlUZ6M5t8SsDSj+KKtEFF6clXW4cGlKFXGY
0Cl2G8tixjWyMNRFt3hwUWrpza58i4yS1gMtnPe4eKFr1vWaH+QIkkXxT6dBsqJ1zv2g0KuZLC1b
RmL3kHv0+cshPHCJ+u6zwGPSLrCSk4wRcgfj5+SM8ArfJfu/fc8GlgmuC/jt10ZHIW5JNS/cM48c
sxr395nblgm/tnAFlo8gJj2WA0PHodi91YMjpt3KwwkCmheA+YEjm2GJisaqEc1d0BWC+47nekZC
NGnIocGUGCLPwZH2XEsYqd995LY1cLs5QPFzHyZM2tBVUsTl4ZnD9H4gbRqBDqusfBsHmdJ37Pqu
m55wCdkHA1hq8ReqMk0ZApWUuGZjbMpO0Aj9+NRvt4F9ZQjG96ImjyFyw5zBXvY+rCAB1j79pB5K
Rf+pLcAiK/Ba13qDfEYZyFaN45DRuVx87aIvabfodTgzBtkhlFYTW3lZ0eQJaglcE+nRiymbYiqI
qOBpuUKAAGTtykc2mPQkYzyoubqMmquVrZxQOC3Npnd0yK5/Uqfw7W7loqpJXAevOkPvRKvyCWjO
XR3YsLYauvqBlfWzTL2bPgVfqPQvqpBgnGFjW+NMf4lN0kMzzzE5ter/AGHiDN8cvpwZNZ48cGSD
4qcEKkpZv/O7sKZpQgjDNshEnHkGxBUCbWKvA99N1z2XMJ43digFC/XPuNTtlwp3VdGPHDv0CuBn
bMZG1SNz6Hs2uoBtSXJ2R9IlHXLi/JdKWfuQEsirCSoteaBFkl15ec8toRBwOI9U6MBEVz5A0tqs
QY71cQ7JmMMna0BiJU0JWM8eubmnFpJTKjQc+WpbMtKr6pXGnYaBENtpVgbACAZnemXNAjqjqOLK
zuZFa5/9uawQIYSPXMbiFR+4mTo0QNj9OqDg7Q75M/GykgSUwlrn9V/TyBzGK1Ax2Z5XdrqOPna4
wr3CocKRGAPqSc3TzwO37K5irXzoo90iTYswQ9iO/6ylwCE8hWVGIp2DQk23/f0M46NCFNsdcbGG
QXKswzLiQ/FQJRq0eytkrudBpkIhfV0fpUynILt4Cvxnn5sUL0Bo2BaCJHaftZGghqbrGyE3ddld
o3bH0msijzkNTxMVbWH2G2ILnklWOPTSXXyQamt0ZSTYZn/RGPRYMSxOTL2H2n9x3YoDL2i7W5qS
4+han65oqcd3Yf/rWgf1zIb8mpgu+gOER0NeZTe+MhrS46A3V/8K8qh+Vq0S965ngrE4vXFO8lb8
cnw51XTSlX4jeikFAugBvR0q5g0+dA2zQhioM9wFzvIEZI/wzbQcol0DKzHPUP+oG22QlJENAJvy
qZ1j2v68ofkkivv+EfhtfY0Dlqj9CrrsMI1GJYyzq4RHL8vDGrf6ifFO5i4CK7T9gqOEvUTr9HWv
QgREiwX6Hd9IzKK5XvEWdDnDe/e1tCco+pmNhMQEichBtAX2A3+EJ/a5/dZlNdYtg4z9Pq6Mrz+f
sKO9fIHYyeLrjDyMli/8pfUaNaMNjSYb+SKuSkrs6LwreigVFMmOoZmfbkYe+4B9Jze+ZlIuBTNa
JnCF8zXnzX7vTwIvRM9k8jUZCT2xs5Tz/b31gTv+U4Y6Ib+M/OWFaFAv6wzWPSy8rm5D2BbHJ1GN
QYwOc5eotlBxNEPwGHhYzexEe1GO8VUev2aBS5+XHb9aZ6bzwvUNNNktJY7x26qmld8WEVCQKUy0
NUbQWzm82hXPL1AQncuELa57QjebsuzX3KwDdCXAH8H62SNtm4fcQvWtpQ1QQjXRFNcta9MVTXgs
Nwb7xFB3qlj3R1rqFzsNRhC1Yi5pQXtHcSBczEt7miceO4/G3Z2B9vjRSgQiaLiXRoXD/wu+EFJw
rleBM5Oul59sCS1cfLtCINSczG9RwIcHlvxAmMrpTAh4EywBGiQJ+sSyhxoQTUF70y1UrtQ7e1fL
PGrVxSrmozZfsZCJRZbnA53npFDk3XgmfXFw/d2nny/i8wBaDyTBSGeip3mfqQhCzAv0e5+5UfNA
NIJrh/OjwxSBRpQOIZhfhYVPi1Zody6JfLeaza7/o/JrC709f1ZglRqxvUdMWLJqcSkgoJAnC0mH
srdFX/nTGU5Q7vPSEyj/sWr2+iqyMUxt9p/zRIMEu5eo2f/3rmsNdPoKtGDuZegGm/kk1Kn0vxx1
sZSxFHe4TmMxTEOrSdkPdDpGrOXPF7leVz6aJsKOKRUqv4kXVuw3TkHNfAJQ3/jmOGZ2YD1g8q3i
GY4SpxepOTAGCa7FO7xI0ZYhdWKBOl+RpxMANZSvoGrTvCBFi6adIfqR9PpwVLxnOUp1IbEwi1YF
B/HDwCy5BWtOI+fmmQhY2A+RHEjocVM7kQ1tU2vKyU6YnGhGoYIjYbx2KEzlbQJNk6BhbgX9es75
dsiscFwUBBPfIWsxy1StBgoatEK1VoW9BOlPKgC+n+oep7Dau2T7vYobUMiuILqPHLu7XPvjhJtd
cUpI54ob5ab52tZNzbA6b6mvevPmnV2jPb75zJcXAhPzv/VZwqf5NGK56PmadmPO0A32c60nFUmh
LoHnG9UjGCQB/jDQttOBiFloG2K9gvr2Co8pVYNnxQegTfm1jYsZwTMV3gYmHfnk1sHmdcXbJ9re
E5ReHjWX+Lz7mJDTs2ToaMpcq6LHAmcEvTd2bZwqu5yP0M2dPazS+AhRp4LRbix5oVEovxAqP4Pv
s5/OChaC4vsIVZs9mKUGiBPAzxNNswAOurE2HTTZSVEjkyOX1fXbkjN3chghcu84YKqeo1fXP+C5
4J21cOr1usOB06LWTWvKQTnMlC4o8zjEm9TXZfH50IK3YH44BpLLQOLvURKG2fyVFIXW9Ch5BvHu
iCrn/wd6eFHtwU3NB+iUf102/KXqjGJpxKTRDvTClj4tboXOFt/WmGRh494uJQJwcXW91oOxAiqi
Sp1L9NJTyRzJbT4dhsxhwQ8d5jL1u4/ZhaFKJp8+w5vyOrspBE58PdLPCrpIu0JsYlUBKEkGEUlw
TOp/AsPdci05OgI3PMdPJV07tnzVzCBXlzIRCggH5EE8JunLJ7dgDPmXnJIqE35j+G2Llc4w6LXS
SruUvD8EVaMb4lTU6Q/85uRoCeUSh3dgEiopjjo3xJBKUq6V1GY9vo59PTPa8MhA/UzU6a9V9P1u
ObD0NK6I/uf/t0yXBOq5zkdpAHOasOp3QieMuvs5iGfoU04Fqf0upp9etSzQJBa58uYhsTdFA/eH
pbAl1P6EYTte7tTweRNuubU2N53Sv319GbrmFhbbtyfGhBToU7bQKIqqwMXJ1xSMJZWkvA0zGr0o
UA/Q/L95Wd9TrxJBI2yiR1k2E1LqRj04NrbvWJnlWiZMN2b2czBu6wk4XM+AMKhn8VTaoxCW4fTH
iYKO8wRE9c+Ek7XEbmZieedqYWgwpwz1QpbArZvRjdXQG3FKF7zXCX1o+sgmwW49Sv1CNo3fJFez
BcyTMW0V7vNFCxBfJH+33uzcsIIWa58Gu1sYbTTP29VvP2/7bU75aB6D55cVNbXrtRu6gM8bjNOD
xXUXMvy6ZFe6K9nwsn1Id/Esizy+CRuwfN2nTzB3Df9VJt5sOg/Vb5HeP28pb6FxiHrMiu0bB+c2
0whtWZhTaMj5hbB4zebUByTXrsYjum0bolk+CmmvFUpfjXgiv9VhSZkIcfCDom8zMHMhBvk9W20i
DfwvSTSPibDZIRTUrABQWuTy4TXNeZQb+nD/N9X62pjYwBVL/jm6NmTrzNFMdy+EoR79BCd/8YSe
ltspeseM7GHZDA5zdQKOljz7JSOuw4KnDW6qB2H79fJIbPUSqczjXuZLL/uzvKhP8y5VGcv3Y4ww
gd64Kts7YOdIF9uAJeGHueVQOrf//J0tyDvK1xXJAcx7r0psDGTathQIHjt+s9y0c8euGo6S7rwD
DQDk8+C84QkjIQKcteWIHCwTajFJfWpvr2uZEqHuxom1vuZ86ZR/I23D3TPnSUt849F3ILSwq6XT
nS/Il2ihIRJV2mtbM5sDnVWLVz3y2E9mJZAgpwIE8k5sV/85+sYS2xf5qcsPwCZK4dVJe4gOkkfb
JXFMyV2BbHfxUkVG7hbldGvcwWnEGdGXAn3N3KtozCtKwxTTzmzbOGia1Ks70n4U6lEGKqaNGtgj
V8SWZQ94B3eUmgrAfrwlTEBMD8P+Y7aG3T82bv84cvtz4TR0mq9daNctoiT4miQK5Y275WVFBfsN
0Bm8rcmdVewZDxn2p7L5bo0BByVeU+/TlRMCw44vh6FCi0Tt/EOLvKdOiL6vu1I6hXxX7JjzPzUR
aCKujHfJuMb8ztOj8H5cfjPS2rz4tZGzWVTmH2N7iEOhExy8/mvL9dK4dTT0iLra/ydUwYB5LuFp
H5WF+00w0sYtQmYulv1N65dLUG2fSKZxA6aO+IHmMukFgnZ8i+wsRzComuGzg0FakcMOHpZ8/w0B
Ho3n1VK87DDdAox32mRCJ92LQgW+txZLUAjzPEphT8dXKfMM0K4NGNUJn6MNz5OdW28Jsf4Ol/TA
b2matxMGRTVETWGtueG9cfylyl9SRNaMdA/ZZEEJfBB87BC/+Alk3YpDCj54YiEHUxb35Q0XfAse
eYFQvpnsUF0+EVQIEwx25vMzVscYDcQC2GrTo5yCCs2bwjhAAvzbEHwXxGqLeXH+cEXPPwdVm7ZD
iYnmm2p2iBlIyhbLKQ8IcLvtqxfw7li0056PVuzA9CaQQuV5l3DtO93DT38abPTZg2yErNjzFKXk
G6maR3MklreDfws0TZdKAR/mbCYzIu0j1QVHyuuk+u4Gqr7X1op+fQPQcFQfSlzR+NBXr4Vz6qDo
ND1yzxy3fqLkE6FobUgQ++RqURgMKY8UlM6oz32fvWWMGkhM0bRa1UXcXo3oZoo6wVvhn5EuuAJw
5iqth6lO+o1aX2iG0cW410Lz7b0ZFJrAw9ybJrVakLYIfMocKhfKb6OnCUsZSy0yExIZ+XbKiPBg
+Qip+B6K6ZhtoLTCv7jKDmgkmtSHBKpTQCugTw0cAZOyufo5QoN+wCx6Dt+dyEorYF2b6+GYNWpe
NvG3XBS8zXGw9CF6TPYxvAwB85I+XrNdzOowUpc4G1YLNNojYFOPxuJ7dFuRvjtpXTRf5XkE4DSD
ghxQJoLtUzEloymGZAZMQXFZEUvKoluh0HPeziuojdcuF77xE8VNIXXHC9QVGFJIAJ0O+15LZIvz
uW6PvsMTwrI6zFgUitJm5GzBJijL/aIwS9te7Au4YxOZsO4VauK3oZCfsiSjxiu65gu/IvGt7tMc
5qOtthC6KvpaxX9tj3wmiQRHMl8Zj6stvVE35qTZW60PA8HUnRyXHBdfNgFjIRohdUKkp66TSDL4
i2wC3zdOY72T+vGPdD7ALeNSl8BwNZsz4T0INF0RNKPtEmBGrlRrkOvaVt9vEOe6lFVltG+psKvJ
Yn1PLIRcD27WjITNuBH7oLZcyqEFhhO7H3b0HSA7BDC/Vz8DTGCODPp2wYkMYSrUHeHxHF3on2k5
jt71JZLKpCuN2rfsmkGmCDeJyWaP7xCw0BU2IQc6rKC+RQzcHapjg9gBC3g0Xf5t+WZsNG5HVfC3
8b8coPqRrwRkLFHEHOZLmzuD52ky6W7AXABfEKsA2UJlnsvtcooaeEjUzZrPXu93npNoBBJXScfe
RLnhIRDPIpFu92B5yHV5wLDQL6JMFtiOIWtN9dFLdZOviqdKd+sPsIN4dWE7+XVAvYVEBYT0bnfz
jwZYG6ZLUbCZ3naDW1guQnfuWS7pwdQSCUOOLs5OIMauiDDr43e5HEfqtijYXISsjaH+fkpgjI0+
hzAK536eG5p9HUZ0pGaEZbKwGfL3y6BOyhk5ZYovDsfNq1Z/Pk2Rl5x6SckOvh1F1Iw2gYX00BCS
5jgsS3hVad+GIPbdYPEtlAMdbmjzDdc2kQUSNBAUooM+VAU+HHRcD3DPyQ+OChDYn5/J15yOinxY
cpNEn1gHXHabelMHx3N342nH0oTK6ww6PPAHjP49G05owegMKjN8A7PBMYEJzk+hioWOsRqWKyMW
sTSg5Tw5HLxrKfPo/A5r2lQASPTjekj4I0gGuGxGiZhl7b6s6Uku7+Pb1Wq19udQhUgF4By/CX5d
wF5nrphogs24QBdYuoL7zOtwjfJ09SoWfxVS7EuvwhwzeALVQYZEwtPS3lbgyfLg7UlA7hBMrwZy
f2VYoWefKnY6ZBE/Yd6O6tAIA78wz7j2aiFX+SzFpt7HqIoWj/d8/bJAfPJAuCWlfsYdKEmu1ckG
Wdc9+fuaa2PRVfaElpSXqbbCcjFMSS7NUTQOP8xGRUddICalIhugR5xku910tkhZc5uniigCwTuc
IFNFgqGLn3yV2DfiTzTQd5aCtjoSNXF0mvFuualdva+D0mUQXRWA621REYxhkr9813UaC0K2YX+u
4o7WxhliNvuR2jPUwkfsV4RJXlc87MYenu1TpVafrbD4rV9GIuinbc1oLHNZHcVsY4d0Up7XaFJ3
e3qqskJ8vUy58wDwWCr6lb/imVsDVsAmVn2RyuE0EzUiQBqcmGRBCnNCLnkcuGtMCGCtn5OtrQ9a
piCZs38qINNDqyVq+ocDjqbZomCni8WIfs6tLYTRplwCxD/eKa9XU77pQKupaQqTqBDKgHHllYIz
N70J0A3pdxOfnszpccG8SA7NRxaxzzrES/YZAg+xDUk67Schqwn8M42hf9mji7hfaOqmjNe0kfUw
KuRf4aYlnfJwDW4tcwJJjZuANxjLhkkj48wfb5WL96F7xAb1NcjPJdHiio0YynPBFLDP4dD4mIHl
VYXz8teBdn5IXkMXthe98mLQ9u2yY55jJWyp2PvRS3ulq4egsGK2PH0FMi5bI749NXG/0OToHzp+
gfyegJGMW9JloiLGQoOicyvvW3jpFKUxHB2fXw9nIE0hdCfjrbFWLjeLW9wcVn32vRKU1aX7rLew
ANUxhy48u+fUEBTrvhYPxMWiyJm8j10RLjxZ/tUljFct/ecyMsEANDroPJ4pFiBGjgyPv1sHRB2U
pRvmJluGiv9vZm2L2EeSKZdaQzDLJbIDdY+x0scXSlEJRaCN3TSJ8EGMUPUqfPChrTt/V+om2NBC
RQFxJnRgNCmi3E4+69c8A5cRiIkU7vcN2NXk/0Crya3w7Pb3ztuiD0bOEDlpbVr47NEoGN9Sm+Kv
r1qRD5vou/C+YbKPN4dX3t9o3hJmSJYn3ij8SGrzIpnbAGjJb0vYzoCDa+BXedRH1UAydeOLd+6y
arFeU6znSkhFSGG5DyZgjnb7UiuX7NEJyjaUWaANEJDaZ3GjinxybVjSAU7afZVrLrVVspn4MxL2
6w+1Xp/MVIJ3WqNlmUvbMCaUFc/BqWsDBtqp73LnBP67atUbazq07NDyhAp8Z0UvS1V7NBKeYcbK
xyp8aeUlfKkWXEPazdVgn0oLwbUMTzyYxZc/ATnonrFdQERKfgj1hHqw76FJ4OyOzKlegCjRvK5d
GMDcjI/mfjUh99tHj3u6NGpYV3r7wZFxE6jOg9dsbtVGTxFgKzjkofkP9qhuX18DLyzjVJY20DsY
gaT0xIW5mg/v7OKiyBWk0t4svQP4IW5BJYgpXwhKarcK9ZBYpUTU/07+ewxksE3k9YRezn577Mba
6+6vWceBc9lx7eyMYE6CD8BHUaziCteJRHNTNR013M+xOZaage0eQk5CsIsgvmXUENEtugdPqtab
0kXLJMjlp5iH/oTKwagfyP/gbwrtgoOHh+rirPFNAOg/KT+4d7UoUb7y6O4gH42HaVEZgsiDF8hw
Jhx9SfCgv1Eos3MrTlkNAVhD1lVRBsmwih6ohgHSw4UKJzIMXjcKg95X1bHue0oRyhsAGdE4kv6Y
mLZ87OBiBuvnvcVjSH0RHM/nmVaTKcY0Bk7sfYuMd0jxhLQw/6sOVzyt86S63cG4ZekMZs+M6v1W
V4StJuduagerkQBFFmNrkRTIpGl+b+lezstSxaWi/rKMpjkwzivSagJiHNt74U0m0/k80WvS0IhP
YV2yUxCeYbIKeamiCeFfVm0JTqMNzIywwu0AzZ7M9RHBXi+PxyYtNKj5j71eMkHAHiir4oSSwTn+
ph7N37ekkASdk7KhyNLD+2tDYC607mcNlCBDmhefkgaIYYIpFniF38Y/xoRY0f+/l2KmiGajABqD
MJn4jPiMkr1cBZbXIMI5K0DEzf14qyypG/rdEBMa88OiLWUa+KhWP2Zeqpj3ICKqf65STsObBzwY
89i2JZV7bMgOBVfPJokWNT9O61RcWWWhBB8FmgfUdzWL0TB652CjRCokveTW5lCEI15jlRv12cr4
lUiINbKRxxXw32HnN1ibbwf+fNSyjCqMNXTpF7aSpvhBRcnMApmIqsSxs/7ITEMgZwIrcxsodAqp
Gls8DGtrJ3Sj6/8EPs6MFxWOX/P4zcGRCVosy8QvqJ8V6aKF1IbHv8JQVvc5k1UhFaJI+BNDmv0Z
0tjykl4tiy+tVxhDv7YtXoKravXtjo3QJytZcfoGk5n+Wx1rck/aB+40ibPGorDsNPb5XGx54g1n
CNAQ4EPc4P49n+7P4UgplNZD60w4qLX+F/JHwPWoFjxPdzPjsuE4asxzK82Jg7h5PDhvUJuELEew
Kn3josDrnYw4buBg6uPn0H46Uk/JwKxLJB1anbmoB6c8Xz/vKicjfmM30CTBFnFB9inT7UqYL2Lt
+4CvKzgJX2PuVGuMNLQyegBTQIpkSx3l09avgKcrEfsSGSb16Od66TKUb5J0lcdm7fkYnMBdjIIe
41YuAHiajAj6LgvnJwOPKnqUymcCnVmUHYtR4E2t6Tjhn/ymSqObX1V/jaQ9bbJ7YOzj8ISEIXtS
MQRT+PfHUmgh6mbsLqlFkQZpShF0JXyo9+viAGtYEKAUSKhLLlyohbqaI8LT4UYCFzxwn1fbSvnK
Q6EpzjKPDPCkSBqO3J2RdL4v2SiqGlswsSlk0HB3RxSERCLnykUrhjxZuaDM97hMhWxDSebYr+5Z
KrLIu2ZF4W9EG0mQaJH3tSwC5qdhJQ1L7otEEcwNyFyGUXQKG28+eoLkBj4It0trgw37llmKwAxu
0JbShDEylYap6QcsjQTLdPpPifCN6oM4mr8zFXUKX15v7xP+Xq/N98i3QWMwghDjJFY/IX8A3BKn
kQC1hWSQDy/4Ca/Qc6sa4gzDn/DhkJfp6fNrIwUaz5ALL7u3URmDPGpQ4nDW6ogPZLE6UctfbPaC
7wn6c6ghoBrsIS8fFY/eii0oGWwL8mtBaSXpASFl1YOY/UIkuTqC25LGJojQZ4rB3VlhRLrCy97N
+29+9PePw8K8u47ulRC8KMOI554RdiN/fg+ppWCo17DLewRNPuv5uNFgEJmNUDeh5oKqiwKdtJ5B
Lq0bospP3Lg6twkamF18uGSuimgBB4wKH6jWaVwHzGWFVQYwWbC7+EgX5FaYVa6iBlyOMzy6koMo
wAzvRo9RCDGTiQKoNjGUH53KIn/y0d4mjyOPtDELN3xG98sGI117+GNaXEa9V9KbKPS7D7+H2l5/
ECLjprOrps+BFiaIp+RlJBVvD85EmfcCx/1zKkNMu6FrQUtW5GrFg6r7d5O8zmj4D+Jl2NX4vxFg
tCvMGmsDxgOh2Wr3dFmvrZaC1QITFX2Xo5p+NOxzJ9B10cz/ckrIrvphKyh4i1ao+axVNY4hrqTx
ububj8CgSUXyh+8RUCt8kTXSUUKEu+1bODrVQHo565jY4RvTRBaDvfXvFjcGEgE2dsrTh3zSPjTy
Tfxs+05LySV+0jeuc53b7tPdQmHdQs8dUMQz0yVSt1NC2fUvTsn/+Fp6RJ4aIRsJ2mk5HYJTNKLZ
C4TSWINIm1qzq+i6vA/f1M+ZuZlwTIeGUHGmA+M4NxvSh+uXXK0IRHJ8ZGZNhhER1J3rHorVLzy6
sQinHXjmUguLG6Lqh6r6J4hbGGpr2zTmnSvdoWFY0fNL4agRYd2qNz8+WBGbLjl4u+/dbJeyTG84
fv3X90Y1w+YUAy+y44BTtzAzUI4VVv0BajeIdmvCXybI+658oGmQadXZSsZiJDGpZ62Xe+3l28IK
3CikPQ1DU9lMTxCs8RiNr/Xpuafwy3dgzH55Y+5JVqcsJ1H421HyMmNC0qavqZsH0KT0TlvcZrXH
fMY4ulJZTa4xT5HssjAhNmZaJkngnvtwKzHlzyckqnO3CwC8qtXdqX2QgprnhPtC7qOC6ftdeCWr
E+uOxSsgxD1eSYotnzezIOprbt5KQj03SD4KvuLmxp9y560C43u/YIwt0Ftazk3rzEMNHBOIVdZ+
DxqXbUbVGUKb5ifRn/X6d/lpQkyZjRNIRNYjMSPoWiUOmqQ1WnP4b7Yc5hyvPASWY+8oJ9MF3lFo
BHBXTuc7CtuVSHWpykfuztMU6ga0ftCfPLGYICTrGtAspKxIHp6nxkxsqNeGoXVXK5wmrj2HMsvz
bXvD0i2gG4zFm9LWgICByLml1E3wHbJP1yxEBzXyHuV69auAQ7XmkwAkbVkkLRFxSlI+2sCjcQR5
ze34NxNfzK9AxzGuIMMKA96gNCCEwYM3pRrlFmlXad09b00qzKz+HzqzY5RyXrmE8gu4xnkQWnBC
NMsD+9/TpZoYAJUDNMyF9EwDacta6SS+ICA+ZOrQ2zJhTSJsLT4HwxdjVy1zxi5ECKYLj931upGU
1mYpDlPWPnolDuB6VriRpKhaLsEDIe5U4kGNqjTEJcraIjj1jMJ7If2rjVS7j16I14Tv1ga/YAhj
TDYSMFY9+oGlDenFSddloiybxYYr2Kc4vvTJtfjtHiyzHTb6pkb25yGc1nxmIx2XUENTUspQb9Xp
rZNcLqIRNseBjZx+k6HQxId3w1YFgwabpmENzuQvkmXM5IzoRUsbaXOwncDtfWaKVf9EP4QN1T3i
RU1o0vCv0pYxmipZxyJjgSM1bI9HG0yboWmNJhcT8fsjJ2t6VW+Sq2vE48Y0IfSPFNKt4Zild+kr
cXrUHdEq8DNnXP5B8XbP/gVQrnpDvil3xvF2+I/+Ak23K00gEK7qhU2d0MRaU0oJICdt415GTDyM
kWWVn5OzYgRTLRKpQg4ReVzOq8LcLQB+ViOw9lxS3Xduoe2oQQk0JGQxtmaOftOsLjGiAOQS3FSu
6W/XWQ3bKWvD48c+EBqBgGUjmwtMaMv12FB081ogvPb6fYgaUGbrAPTxM+lSTR6didIY4U+mHVvp
6eUowoRcW/ec6CdjxuHC38HwjYqaM3CNpCgKmyZssMgyIL/gVKBigeXGdzAL/CTyPT0m1z0UGhuP
SqlCa4MyYNh+QY2XbMy5UU8futkuchGgfpTXKtrFz/vEHTLkV/R9L0f9DQdDgeKkOfhoacVfZKhe
ye6deVSWKVQkM+YGIG2m0edgxbmq6tFgIWyzWMmAm2efAob81GL9RcA3M60DhReE32zHKxYnXSdv
toMTnkJWs3lyziaMmFW2ptZHJ6UIz4tJZBpgidtQ6xSouu4VUZTZVZC19DpbNILMwGTfluwhHzvy
1Ma0EOOeFfXUtU9wqmdynzBuqEADaPSi0yMTfKd9AILmvvJT1k4U2B1ntxwzs+0dpXH1e2YfJtQK
kfyYNXppvwzGQofWa3vlJuF99Y11FGVK/aotZBVDtTxUha0aCSptCL+qoCIbQ1+FRR/wzkIPEo2n
uI8iYOed07A7vf4nVFfDA3UFogfAm7G+YwxQcjA0OnMBu/ZMDvqloHWYFAUE3V708qnt3nWqSIJ5
fpR4lGE97P2BUtOhCFedIvPtXH+M6No50Lb2MC4ifmzWOJ3G62b3EX1fOWBOYGoIkh8Vg/hBecD/
rjEMXEEl++dw9aQsGsWNkjII55R7sHuVqA4TqrNXSSt3fn5qcsCaspJeuewvpQ9EBasnBANXb4wa
dnLWwjj1W/mkscMbfh5Oo/uyvU4rE8mlMH63h8qUwaa3AfMP9FM0AXcAcnIlxUzCdt2cMucvX0Ti
wfCjAx0ciA0a2+CNIbxPlINt9NK0zjbWEmkAb52kGN1gco4l26J4n2y3fBrH838l+gMf2anUUVRi
Mq0lc50zw5umcwbmkzwAhpmHhs5nwkPKVhpM8eHQO/0MXbS1i4GsasWH1B6rXigoWmVWfV3uOylb
t5SsjGT64Uy/0KwOIJM37ikdsIxcjNgfYs7laxdvRTjirQ/vabbBY/rbNxydl91RiwAWo1x/vzRr
dtVByLUUdbftowepQq7cVEaI+VdK+6Qx0BgB55Gl2wqU5vhDsM+fUwgmwWF6c7b8ssUy6iULQgQ4
De+BmzUoZpEJzDF2C0w/EyH4S86CuQANbLxbdcW60+wHrfQOIOSd60LH1kK3ukBjFmO/MA7ixTRb
CYDlXPM62CsAse+ZCPzcQtXAPeOyekIbu2FfggosVMp5VS1zngCgtWx2IQg64R09wWGtCh0+xFC1
G73oiEkOC2qWRnGD5FliVyF8hXcSedposRQ8lIL4to9UenXfSF528DpSoJ3TLs8IpayStyojkBtt
YFXt5m+BmnolcuxckkisfNQz3b/PjbslCLjoDPwbb7AB79ioT97lhk+BuAyllZPLDaIRHMeIpNPu
gRI0gLatmVXN1R+2BF7mtAx8/d7wDzord7J0DvGcc1PeqUTlaDmFdTslKg0srPzAHZmaKozvi2ZN
X/6x9XI+jjXAGSnPeEgyy9wh/7LXKpx5vU/p2/MW+8o10ZUyirKMCv4Xs54Rg/J7HK+654Oa9Y34
Y5EfuqwEluTGk78lVTjUCcMEd8m8/OZztCSS3VrgwPlpH3bRhLgeTXolacA9xAzCUscY+MDP1sSf
1QWdMJ25OvVrmTUXLU8MZJsbdwliicJ9vsrJusQw20vrMn44sPFOIJoO5lj2OIVP6yNH4v1Se+FF
KqXNQz7iW1eKx+dQYDIIShCfR6h2BCYF5mFH1QuAnQrJ+K4nI9u8YjWnQeOiHVK6+KlwDjeTtxVs
TllDg7bJ+q9wpfNyVxxn+zELenXe+SsWnPKMBOjVzJj0Wt5QRzKAHTGWr72hwd/86xDsoc7plHmK
WdM3WgQ3ZKojQ8vDkUf2Hzi2WmVkUKLIaZ/kCIOdsAMqPFsUlQ1qrmUsj0rx0/d7Ju04CyoxXnvQ
By3tzDx8Ygdd7CvcjqqCjI4i64D8uvOJkpKi7lmjkUXukifEEHJRSTHT1Q3K46kThy5OFWq3VOg0
4epPMpj55Agu6dC6ukzFSfC5n0YVi6LttODWmE7LXsEpClJbLiKCuzwgV5Rsg3gdnfXLxXOGV6SI
vY1UPw20WBGFEGlVHu70HSmOyhYiPNL7LhykNbBJvt0q0D6ep12WixB7MvKuJlDFHc115krHl0YX
49lcMm7r+hxsmGtVXV371Jf/Dztwe2DncDVmewyldiXpgHCoNb61U69C4a4Tpq5fDZCuXw6SbNmY
1CA2eHx5UhPWhypCyqUd2zmlvYt6SLFeJ6RTLluMEnCwvIPyQP5pe9lSpiANPrumJkHqYJOknudJ
Hu/13zhggMN4W2eHbajtTxIL5OuLpfsjtgzY2uB48CF8xuUDJ86zui4MZJidyUD43vwkl4nbgHTX
bMdHjfW1yCE/nxEHOGgqrcaY5w4lYJhoi4oP6ABCyvtRs5dSPuym34sgeVgzpUlNz7J251UZdmsg
x0sSMxgWA3HxZaILwSyxdoZK7TEMCtLkBoJOojrJRZqXLSxaUSCoHmTv+B0Htl4VbkQMGPfbIi0v
dQb7XwfNl9w7WaAya7DYLz/nWpDxqUunreQ9Qr2njK1oPuoa2iA9uKk10HGoXdx67gLxVc7tglrW
7UjCPrkrH+OZZdmS27TOYzOcjVE1EHxnAFA7yP2B4h5TLxjwllt/2cSznfyf6kOLa5R9pGalfNSh
LHiOWYMcHsqjrzy4QAdUmn35OOkA7ISY24sDjAo0OEhrGIT1RSkzctKvLaKOSr8mVOgRJ7t5cUQQ
myUGXYEZPhCn9uukDZZNQaIIdhLk0bVb48qf9gjsc+dR67S4sA6l9jQ1ap0u0YX3Lzn8KOf1pLdB
zHC7oo0O+o3fh4M4Kifv8hnLmpFDSPRDxkAB8DcPEV9EI/ZxOW1iRlV1P17BSyHPVAiIEPkgoAFz
l1qsDf/7Pz/8ejffyDcCuXnLEpZWXUIvxE94Rjbhxr+jBF4LDWSM82/NBChjX3tWQuXY2OxzRdOs
ziino4O0nqWzStOta4CXK46Fzi9tOZa2EenA1dEnxYqlNNgsqxzYA5gtbZ5mskKUmwzdEdzKOm5x
LQDGoWMdKTuMT8SqH55Ngz5DW5qf1sf7vyJ6t6V8z6RQZGRWiiTWgSjTWR9cyjhqWfNK6A9dOa5J
t9HhTR6QSiH7ibsoh9Gsp8yVUwBoyTqF728gd319Fmw9N0ZXrUbN5BMouQxRYb58B98Le65Lwpaz
NX8dK1+32tReoM/Lf/7zed5PIMqpZKYtMuWStU4SpVxYnUH1F0euztPEKohFu4pm1z+E86V7V8Hd
q1tPVfK20NvH6UwkWgZNOOsBahTaUPn0lXr94l/9ZvtlzuDIDY5eGLNPL35lCRlUy8GCXgCA4eu/
UV9fEihoeeb4R/rKrnbc9AE1OcVEtx9UpVotO+96ixK6VDQYcTJBtPgJuuomL8xuQLoSkRRWvY0c
Xon3TLIZfppr1zWlizy4YqU+SBNp6/L0j7dv5Q5IqFRKEqv/2lNDth83cbN+LPTTlyaZZQFYjmpH
McI9u50KpQSzbSdEnZOWWW+9biHpRPBu1n9/vSvMCptmAo9flERB4W1yYCR5I0MhNW8pyRrzj0YE
lqeSH6u4yeFI4VbAcT1/z/uCcFjQzcLN1nbErKxmCpbrJ9JXakzN/UfR1APmfn2r/L7fcR3XtG4Z
Glj94H7tGb6HnLDLRPS2Il0tlHidq9eZ6wm0jA4koxXjKlk5E9K6Qyfd9G3yXnOSociQduTcS4f1
iMG+HCq3Lt7YERgDasvPnXp7MdFgqzlIRyIm/0C4fLHtO4bKWI2UeBZXPtE0rrsbf33EZY/7NQda
sX5aUXa3GcjdyVAYQY9p/SfCWuJE5rIcdcALp6WEFvBXmkCsQfl3uVcnveKdVvBFBjA2HBh5pzxs
StXyVK1wptOfBddFNctGlDmtYUnmxvOAHsBmjys9SVrfeZT+xcnI959lnDELjNfvmxArTdTlhCaF
6mtPhBGZpzE+uwkJcp7OQDq7sJRJ15RsXHj+gV+K/4J3bZT0hxHajZNe0gtyC0Bmh32SX7SflXBS
WUFih/PzHWxK5CpFrRACfNhJVHnbFG/rjSWZEzU4nhlI5ZSgc4D9t5eRpQ7rDEVmN1be2fHGWEOi
5mK71H1uJ6KM+ea4vCxjedH1MNJvVuJY8OEnXmwjUDpEEWkxNRFPXDBHRzM3m8MS2Xda8G39y9De
3o6YT9L18WD5NKV7KJ6C9Dq9I3FOUWkY68z1AoTueJ6aBjWvbLmfMODy3/RDK/aDiTbIGU26xxcn
7vqyJlo4bJEMomP/oEEBNkpgTMsw7fhcZCxaT1MbJODNdoj7tVyOQ70oVJHtusYD1HmKceCfwt/6
Sgsr7iUOcBwa2faFCMoG10wlgFqnUc6wYP+1gjKz53v6s6XZyq8fqO8knlbIBk0yuLXhIW/VIRrY
ZRzHRfbvkXm4oWHRcty1AdEDLcPjCYId7vICYONUbgNULXX0I/K5OnmuSlpkE+Zi+7g8M+y3gBF+
VhEGZPcetOTZXFpq1k4FchZ9+kBFzau/Xg0t47IRv9NCgMQ226rEI0kfbjLdq50aPVpkf2QQKw7B
XgWiVQZjBc/M92+cViCxYIWRUvym3iBGfCFQZWRl+1hPB/jeLnnTyHeQ43kz8QrwaJYFsV96Bg53
T5EPAit1Mv81QksZ6MRUuER31AU5U6WI0wVu/QcIYR3eCU9mjlWuJeE7YG/NajgZS8+7qhuT1iT4
iP0Q6UBYSTsCJNvFYyLL8/ofVpSldOBhBvQe7Bgk18sw39IRFE4U67iGCLKYvqjArqmmpW902VBQ
1NR+GvOKiJtDXwUdPJ1zBqrKyqAMwBmOA+ZIleouL9HjcY2IFC29OuGi7+QGh4vmOsFLxbhA2QfJ
7RUqGdLDq129ANfiK82a1ViPJldSnnjqyULPG2ukGmx2uhcCsHcaoinVMl+N5KUbLJq09W+9kz0W
Gh3+xXpDgf7ufW36/j1+I2fc1KLELOwGTMMfWmWm6fVHgrM6pitzF+C0sgFOrAJV/GUNBuM2Fa1P
y/20QIjydCyUI3L8TzTyWiGXN0nbB+TBj8v1yadoWJSQkCuPIXvelfuxerWHDsGskmsnsHGQakmI
ngzpgI+WCzO2ugheQh2PlhR0Jz5X+QzQjHmIaDMB/Tpk+E+bemPnLo8p4MA6mkfyTqyWaGaOsnDF
ZN+lZUPW04dPUcSEcbZutPq7FlGTDbsgZg421jXREd1WnChlr4Yp+GCRerm7TxfhjXV/1AXWPgBu
ewfAX5Ftz5fyQhCeViMWdgIWuyUB5lnYwY9A/h1I6a0YrqnsLaRtBb/molfu3AGD1/fDy8NpK2RQ
Hl/mY29N4wTGZwKjfEwLSoZGl9PyWn7qjYbr0nTDuDEuL+brDGHCawHRb8m+obW2u3vBHpm2VD9I
k1nr1RZu5NSPmxJ+u0mFFKFXoTa9Nl9HDvTxf7BqmtiFiXlZVfQgAWXzpts36avYDXql1pkGijP+
j1MPBC/D7O2SZTpE1DcDQydnnc1KFF01ZY0w4cFG44lEjTEI/WJ0Cy4iR0PtM/PRk9slxjcAMvXG
XliRZoELETHGGRlBebPv96HZx1Wjw925G3HHwrPm0r7coJ/filybEfa9jgZEYn5oxvbKxvY5FHOv
KQBfQcIEN/hu63aR2IamjOJRckkbeHBeJigd3jxYgstvZnaT7Ogq9dj+AWj2+OI3fCKZOBJCr93T
P3AFVHNbk7ysOfKYkCRwdcyTyulBYE0DZnu6TioGZO3IH9x6RMhJAAHX3b64L4FziTNPqT3WGc3Z
4EALVPOGIKAhOg7/cFiq/3ZA/E9woccDr6ad7dXjqezltwB+O5/osJlImdxY8S7ECZf/OawKpE0r
C6/zeWFRYASehBDvUzC98IU2Y4/OyVPWPWyeZ7X2LVakXq1Z1l0QNxYeDWY2giMiontYsFIZw3Z9
6GjsqbeP0S9p3oyViafdzA45LN6fbY4LJvdrwcK85w/PvgKAUOLsGA+masHhwjD8KOtojnkMXkMt
EB9ROzUM1N6KKBTtC6WfCIxR4jANMD5358i98XIwniqfhXrsKOa0EWfgJfgooTOm4IjaqXPxRifZ
i26G1tEeKnyT8hdMQKuru58Bx97SYDtrSzRjiyXTreXJIYQ+yp4BJ9wnv1CAP4FrXsN2CxUbqpku
goQwh4U/FeIcQ3g5AkrM9hCoaOUxVinVTWOI43rUsWLUuzHlvjfkqyS9ndLPCYbdfUDufjudpjlN
TOIxpRm6QX5B0WX0U4htr6hRBOtISYUkVEEB/T+Vstxr5gvB4jnH0dcVXzzYVVJsVmWfhcUtRsPl
eKqUYofdukDr4LJJmThuulUgUCCzyUzco4OL7nZhmV5AG+rjis4Ru4G1AjjY/lZSTw8UnSpHIk9j
fC/6GCfyl0LLaFJ3B9c4vjvcp8pDvxZBrB7L0QV32C8PCE0gVC9/6R7U9q9a2OP+TgfTX+gsfqW6
Z3oZv6NBi7ud00wvnQfsYJTmNuCTFKkyRErA2+Q4NLemHTeFOy8SrSoibskuXPb6pDqLTZU8Qmi0
A4yNDNdfCuJJ48OP78VpqsHZud+UADKdtKx1JIvfHXXuDr8rv1kIXJURlTyolaUF79FSCkvFf3Cb
uKvR2UMFrTZZuqAO3y+XVuC5+O9mAWJNgk/1xfKxl7MYKDWjJeFI5Dee6bDo3GetUtjwnM2Y8UBF
xOiJ7a6OSFz/nz/dFbwyFMtq1Ml4ZYMsVv7gY+iaei4J+NslPzEAV7QD0KErUB5LtZ4uMkXwJkXU
EDlRUd5uN1+o1mWxA6Vjggmi+CLYnyjsfrDnRLXW6LqE4rUHGUlqdbAvbCj7PnLOov4B7kMm+aTI
XiwNEuZocSGkPifgOx9a9iq8wFGRacPZi7zAgaDVCrBUYL6qpw7hF5wexPMvd0WxEIT8fv+VYDC1
bR1TbnpRTyPomEfSBQd8VAyqr1Z/oWTNKwNJhMmTY17nOmDGld3ecVP3cdgTcu4kp9SZ2PnxuIXV
StDupc32VrYOlnEBnt2WV4S+oDBYBScwzZloxZskts9vDK88FM3UyyosRP1ccd0LIU4cz5cfMw3S
x1b+18vmp1WvV7LFPRZhRTci87PUfKPMAca+UqvatKLblEPp8hVB3Yh3jxy6pKNlhi59wmv7G6rO
7Iu0vaTWKUpVCCIrDLtMbPBPl3Ah8ad9Kf7PkWouV9rTA9geZZXffWFJ+2FrSVOuF463VJ0Aatur
1VSPBFrDFqtXMkp3wq2BlAIjt6W2q9vg23fy+96x2XlBaIhTABH4hnHZ67xkfg3vo5lP0Bq1wu2o
9U20sX1hole67FI0AaX2GomV5MHbde2A1u30WN0oZ5Kn+7hqbRRVIjNZIOy0Rt0YBVxqrKMfrjOB
JT8iQgVMvUYxV9/zVqwPjRqRUkwEtJWg2nw/Yl5EVWy0hk/HW7gG5EdJ87vLS3E0pGPAyUEs6OF/
LV/B6YJwTZWDu2igBcIPokG5xMpSPVow76Bfo7+igkNRSOAKDMNftUhpWV1hPJ9Dz2IAEUI2Sg7w
dztp7OH6YMjGeKKxkCIV9HtPUE9GQUsLOpYibPBSYcCfeZxMVctpBzH6QsVaNa+S7olru5TQ38EO
uCJWl2jcLN+D0ieIkn30PG0wmn7Qw93BnuNmr5zhcM/GFVpxbPM9MFvZ3OCJFr9J0xgNyxEiiZqr
4NSOHL+uqy+e6zdfib/aQve88A3yNJotm09Ozaj4X6Zl3JvBlEKb6YsdqPEzRMc4aE0IeZ1sV+QW
+xiRbZ8oVzUfoofBVvh3pndu7DQULnTcY3vBOuCjjnh1M2zBnnLZ2d0JGYdv4MOoLoMtOQQD103u
UkYYNyqkyAKWx5nLwmhDwETmN6mgynZg4BVb+uqlntw+rlUctGCktNpjW2Vgsm5z9LfSSeQ+MsXT
zLf1n9s2xHRRsztX1JkFxMEMXdGZ5lSVWY4mb97Km+fRN1nDGv+stW2jiJOTnuJvzeNAcC3Z5dwl
iSqdKghBcYu4s39IZNxUkDZhz+pV3fHwCRCE+wjMfw9gtvjwM3zYg7as6kgQhsvoTpM6ekZs5yPM
UI4VSSjHjaZzA8gjCg4pWrLqleXYc4/GphKBECNNuBTAuMMGY3X8AAFZI8PXkMKlWwCsshLURjQv
gZR5hKzbHh03S1USF0g1kbEWrJ/rNZaX+zZ4aYb3KybEhVKT+VJl6+sjwXrSfy9jsmPQRzOzQaLi
7BroxqEOs6Bjocano9DlNKb7vdghN0rGf3TXqWKUJs31rlWuHk5ZTYKipHB6a2qeoIXyxZ/Bnmpo
ajaHhwTqTOzkHk2r3CfNthvfMv+mOpH/LRe/FH04lcRStDb5S7pwZzvLiOR5vlTP6bgJmpgoE1IK
nqXRsZJIGTNPOVqsWZwSg3G4DtN5P56XXAYiA4YV+t72UUMLLfEifrzl/sr+76YIbGrfDuX5eRRz
TSuVHZJR2LEl0xT3+KUik/v3G/vi5IJpj62O8JDft5K68gJsZQw4yTSwES9cu+6kisyNCQTkcj6e
WVE7nGI9FngA6i1PmRXI7EOER/y4+k1btG27Rjfg/D0uwoHJ6KHpOj/df1KNBCAPrtDNOHadjLAT
AbYhCkAzoxhm8JfskugAJnTSEVlpbx6pO68MnxK6mTIoc4REV4RE1RBzk/TLEw+uGnH1K4eZwFuX
V2GwCV8oEFUENhtp9DonU6LgSDgdtqSPNVbzsy8LZV6sztfdm1AUAkapADEa5iMtzBPq8UP2koKF
cS9UgJ3YvZa6yyMk43SSrdtQUHscnHqdsfMtsJOuQrpEwXTtzVm3K6KcnqvXbDZSdLai1yBAQThe
IIePbjf6YwFyPnsLtk6uQ3ogIJqWVlRhyZG0KEHXGQktFVz8CzNLgfCetxB9URXg3nlXoIzvigzX
TpFpVHBgtg2HZsqY9pviN/+sYozH3qJj1ISCttSjdLpgollAmQGf0Wd+tG/jRrg17yEPfJaYbpIU
c6348DrHw90COFvUlmc4IxjYHZ2KXsLmMcJmai5e5RCUrmhiLaDer79xkYWg/126+jhYpjVdpGDd
V5xSBEA0YnAqzsdtSWInoYRDFI/Q3n+ynFiv8wtbaKAPr3U7HqoI+vmYQSfhvaBQpHPESkXK9IW5
HTeFA14AxbwU97wWdUlbZ9UDZye3xe5Z2NW/7L/jYdF745AGHOKmC6tnTv8wtg8X9nCIYpzEWQ2o
VmOwEa+36QrS8PyPmccEPJW1ru4k8DfGl64hDEBmCgwI2XHipfKhNKYAKKbmsuYAxYSJ3k/Vb4Ax
Nx+uVp0RmKrHvXRSThgt9V0jLSh8qRZvARHE7sPWF9EtgcGzZ9JyOml5Jm44REfMmsW8cA8KTsmF
nVIcDZCZFuWWaRSn1B++TShSazUzXJwcbgLq/WPX2ePhpvrrKYx1GdgBXv76ZP7VM5VbyVF7Utj7
p6dZjWo1Yz+egIiaY8iYA6BFgMCWM1H4uR9ncJKA8RbO6eh44pV8Rg4UjQvzG/HG7ZR5BKfdErnN
d23Ifmqy8ZGBR+OS7KTlDcZZOKn88bwFCFqE/z50yjsuQwQck6y5avkctLJfx3JNI0v2NFzmZQpi
SkeuJ5F7GL8nR5HLBPn/8MwvM1pjR/mgzA2bg03G8ul2yCRwcIMQaZFtN/k/OMtX+JlRbPgtB9DC
h2sx02DiwgHMcXJ7GoETr65sp8xjpbAAcF3lKFHNC++QOnO4IejI+02dfOa9rDVUXLbS69E+weyq
NUT5+Sf4gkjEfyesGZwhszjY8WhPLcJe1WQPHI5BQ1sxlKymqrxOmQLtu9TGCVIEZCC9jxWOWcpy
+c4kmgCwvI29vuv6nfdappxjQ/D1ayGzY06ad6JWtMshz3iQJTBB1/2hnbdPy4/kQ0MGmr0n9Ih/
BpA8jShDda7G2oZKsxPn+4EKnKhKaBl7DZkrvhk1CJH5oifRfh5YFhnoW4CrOj6HNUD1yVEHP1to
B5SKCUPIJU7YFiP8g7kAZ3JdXR9aVp79o9GgsEuS5ttvvH//4X5SqpTvYrt5Q31DO0OGtl7nfXVE
5p0u30EAe6Ol0vYJ3fLIjLeHDIrPV0gdDG3LXmgMkkUAMFa9fmHcMppG2rLSvYuRAmyiqj15De9L
/iashJZvbPp+jmHdVpc3D+gSymAA8G/HNCz7loIfB2Ibu9wpmcKjt/fC9fQONF+mE1US49ooYj6c
mStkxGGWqNRY8fBflPSrNyPdJsFX4aXrTjBrk75MZm4nubtPSEVombrhz+Qn9uxJyGLWGP/PzdMG
lZHneR+o1HqybwM8lSqcm1DgkWyjj+bxKI/NwojZrazYl2fuJsz5ZKNpP8KTS1njK0sfpSLl9yQV
2Hgvi+g8VLWkw+i7qf3uHbtYP9Pv/3VHFTuNE/5RPhddhxAUJ8lkOt8/VhA5Lnxh8XWI8YbIeAmS
z1fSMx3nyKD4DanZjKjFtAWpigR3li+LEwPqvi04wlRxwVUc2KjVVdqelYOIGgjbSwYAAcJSoRy+
d100mRRMKJ2UFLGE5XysorqGSOS+mjScRqpH0Dx1BUznXcIw5AQxjzvwN81GcB6ejV9duqgXpxh8
bS536XNM01TPtQCx1dOtULSE5ZwP5FIGl3lPbq1SP6ZaICOm8vs+3iNhPm2zCMW9WcswSj4qEqPA
gTTSoulA1JNJdQLdtHzU9K0jIqW+ZH0CcZ6T+wSwJGl4E6qMsMIcvhqnISJ3r2seiuXHyKEv4aWW
fxQcKxTaOpDqJtFt/A6GflktWWDjNkfXNucUFWdCzNJUPWZaJ5IlkbXbLHhALZWLfpoq0vWRlOeR
oMJIpYWWazADPv2O0gfKsV0K7HkrY1bSZKoLtoemEo7GHrbM52srK30W35lstOYR+n5YB5U9l9JI
TlvTP1CpN4HGz3VGb1/KPt/AnXw0EUmRLu9xjg7W/30s0rHM4IPrSv9Wdgw+2+Imoty6Sv1avTfC
uIKjOUUVmgkEu8Ic4Nezwy3Y0tN25tvhKtM7XqHkQwr12X/x5thDOTwVINp8TwHt7voTQn9unrJd
7FqmdJPVKn1cahCBu5qwrnGkhhCNq72rmN7IE4UMGh5qv2/NoolK/NnrfTYIkgyLm/7Io+RkQltl
qqroYYABcbLWdNTPXeWonsK2TTApYz6Cg53DQYpRYkqAW2/K3As3q2PLaMviJtgbi61F5BQcHzef
AZse8dnMnNTeycbPJKq3mzoikxvkCMjWuIDtMYX8cJL+Edmhhn0EXCfxRq2DN68pllWZE7wv1BFw
5G7GZTvii6sE2qkt78wkxXlxJbDYUiGOGzFZryhHNdblEg/51KCCg1NK5iOJW7LCDXWSe6H/2ubp
eGzpoh3LaggsIGR6r7Zc5zTI+5gYs9LUS3vfOtmWiRso55Id9bRGAjPNTDQWtqxi9iobBRRJdYi2
638SMiqL40ueaDWqHSsrseCcU53ub1emRdJ/1Av0GHrco40vkTaRtVTAOpisqwqBEj9r/HKTwYxf
o1CroFGs9a4N5UtJn0UQvLrcUuIRtGeVcZO0HkQWiT166+QqAvPdbeCpi3XlIXBZ2eJUONg0l96/
0KqwEOxYzekUPk/V/DmOHX3b3LLDB8KyA5wuTYEG+8EcrAzGtcLYulMUVsOKRQ/MTHAlZVoIQzOZ
X78Qw8HyGXJFAJz3tU8TNOvKOIwCnSvjTUd2uUGw5uZ8gGLTK+L/W0C5HXF84JjlyIs1UW10XP/u
SlxdqbCwVdhi675q6zM+JHJsGSK0xzya8y+Lgk3GCOFtJCRldunlKyVBrV+NeDLK4Tm4DKM1RDpP
3KArz6Um/nm/eGAm8LXQccZDEHeCMOKA233v6PQNcC4pl7Arhb18IgDKKOx3hgtainvbbK4U1q3I
D7Y5yle/CWjjO+yH9QvvyUHZhkJVYVQ1E93OfEkTUJfjVE0jOdiaCaYEO6X46wkqE28ruQAw4XZp
BiBFCCniLI4jN88w7CyUGjaZG/N1UMES1+HsBnVAU8oHs6aA/m1ZoBRqBXVSTp/C2A8J6DguUQyS
gdAm5YO7SV0cuN8ZJXXMYIzCXRwrm/m+pPnIUpWYLLTLHSvzgjXiwDBoEp5E/79+QbjfgObnRcUr
wnOljMx95YC/lZn63VwUPM9nSAB/3Gxq+6K+eFXInTHrBVLWfi+Ir0PVvIL9fqvK2PciU6EPs9Zi
EfdR3UHQHYMBbJxqD2GbF0+dkuIJ0IFnnlDKZX75uZCp2C65JKDmQEYztSNMOUH+P2VD/DBJi6Kf
ONLTmfoCRJQoJGuSNIu/X9QJKhdWcZbU57FGAgAyXq+KdXu3TefPTTvCbn3ibEYzTiVVUGUuJwO4
8q4DD5N8CAs8OgexdJObj++emQXcGXfIcud57lMJmPb7mwsJjH0x8LqrQnMaYKTejNANhbBeder4
HgKRznS1m+zC02yOqyIgBG2B1y1qkrI/4F2BWT9gXKAbx5cwYyA5E4LH/yghGj/ezip3IaSR8srd
+TyMCA8aqOwIL/9goNMq5gYIn3bC6+eX8M+Iq7WDlIJ2rPhnaQ3Alm98bMOxwwe+xWANj8K9U0YH
DQEnHxMRBig0cRuD/zF7BM1QKLenB+VCsB0BsDIRPU5spohHogUAN4F262VZZU5lqkZHvGXB/qE1
Qyk/o7jrYchtARklP160y/o+essVxbZxtKf+SwJnYXoO9CqqZD2xmoxKkK4p8fdVFV3FCZnGv54D
PUNU/ycyJ9iUpgJdJVXNbg0uxKQbf4CQ6ONeRdqf77oHpQ3LOp8MVEKJTj4yhlGIqJY/QGGXtcZh
rwz95nyXuHxYAYJ5bMRDzRmOqydBJN59fniSWKA76X3+gpLVGqmaUqw4R+IYddsTogVaPXA/xlxl
hMlL4hZh4o7XgXXWYrUBf8PBKQElJSsZqlbinPesL01JSxZ1Qs0o9XdpL4jikWVpiaTJGmdOTmLK
E8N4Xhk9L/WO/UtK8HIGIVODs+imH219qrxzJCdu5Ck+R0JxB9/Z8N1vxckji75len8HVUBmAN7n
7lU5zTQc0rGXLUd32uRuNYNj9hi/q9zNybjJcZXyu0sL8MVBTiO1tnU+6EBydBbUeX/MWgynOsVg
z9WLWCAfj6dN7TxHlaHXWYqkiq+ULo2Y0Rl+CtDwfKsVfJbOn2/tCoX12HtCmpP8J+xHJZlzWAK1
GMrVJRXwTTDzkKoI1NnXh4+0Qz9Iwq4zLR2JOV2xZv5NLH1fjNcBllNgAlEY1cEZtDVEf+Y12kRB
omlC0wghpOghDSF7WAR/OrD5ZKVf1opJyP6EnvJ55H9UNATafbsesrCRgcNkGl0WTO2SkluruTqv
ZN7rsI9CHcU//y/akQh65/QfJtU1G3Q4R+NNYJMh7BX8cN6dCP23MRyG5tSNb+O1BK8f/Z+uG70u
U0ZHcrOa+8RQN+sMY7WAgDYU4+sIpMa4FFFwETPF6PKDct1RgyD4LHRK4B1J/KvNk35RAzH3NPui
fL/X2UQlg7/nHMJeR75Rya9nI5K+Pp2y+Q9n9umfhIDAxd3mthxfvcp/E4rS6T8xCu01G1gdZHa0
A7jweL2HGMdLLIigxNKQ5etstIPCRfurYKEUEBJNdjpS0k+Tq8PA9MMoNPguhWNLoZRpQ1MzQSlF
/WX8iGuoLAYjgkOxc1JMyduFpK/v+WRnZsYHKDwwEWVayL280qrgFodPTQKBptiAZ4RNdRe0jAbF
1En+ooegH0rbq+sdtRmjPbh+W1AJgowFX7bD9abuxwq6anONzsAXDHRYdlUkKNwM+2nYizQrE10O
ROcNPM5PPXCPdU7LvQke+wWbSYcsxz1eEk8+9PxrwKIqZ2IWKhdFwvhUK6tMO2Togq4pA2FdcS3P
HgZobHHuSev3Bs5kbmyZN37C06HecK6li2YlMvTq1+14RikhHx27IsU8Xz+9+ktnjKzyhLZfGD+r
0rw6znDa2hlYZEVBk+M4Hg5MrKYXithpnLqWwyS2AUspM78SKgce4BAMfXx3nghdGI3dIFPEMAcA
XAcvG3gd5rdUrxuhzpEpZsAUrkLG54a/4VmAxXGzmAiEpTH3a0rjuaUhtcVFyDnBud0FQfkm4noV
u7ffmYlx/IO0qIY0vzFj0sGd3fra03d/IBlfk0M7BmmrTuYs9BCkR1esVOEkvGrUHQgJtmzGtVCw
Xs0Qj/SPvflNfvhzVf2406MpGqMnl0rhc3I+XcBclIOQKogM53B7ShtVS8lPwYKquEoS0/yt0KTB
264GlQT5fpxixuR8QZIyn8pPIcCM+Sf5GTJuS4Lc1D+q+wsmAko0PO7MuO6ChkP7K/MP7HFo40kq
VqpK5wkx1IdDOZiyqTp4Sf09y93BVazqM4svLEPglzVw4Fei384UkkqVsDrnjD3M4hRatOlKuIeD
1106mpcOyJ69egshXhhIcWzy/3YQAxiM+5N7pxGWBcqwbq0yJppNg5Kk+o3mYFSA0x0nM5GuU6Fc
68E3wGVLLLz+H+n68Eurv4FJ2Rc/B4I1cMWYyes9+9SMhshEC7z29r+mlICPF7kTpYCTOL31LNUN
efeThhr4Bh2huZv1cMS3dQLjR7lZj0xId4dwukZ6ki6YI2Y9e7fFzMt0A16OnAjQBvCYykMs8oGt
g+QWh4EWN932ls64gJqNTM2xgvvzJGUSuVX6LElBgnymD/NGhMUSDqEYlV8bKuZIaJxEuzrLhXPI
E2g/EaJZFbgWEqnVrDpfmKCXD/vtz1M9pHpj0yoW9Xav+WMV8BB7NuodBsGMxuc1Ymbhr6Rr2tfW
EvtJkBFxOw3rJHB/1NNrqFzCfUPcum6NiyZEi5oe1B82kNyZ0ngqwbZhp0HQ3KwtYAHrqjaLv+Fc
1rvW4I1JmAEgW2p4NwIpJh7EDptvpJ3UKaUIfd7PxSt2XBfwpoPhT/Rjv0r70CfrZpGeAfVBVN3c
3+8iJcAVvriLSYm2zglYh1JPomKmHOxRJ0365tfFX0mUUXerdmn48gBrpp5cjoIISg0kfPZmsTLW
7UjPdzc7ApKnzh3hQaNik5qozm5rRxc/h2unbI/88dLp/DDq10LtgzqttZGAIgooN8LJJFroVdRu
Fhpd+G3bI5UM8dwwMDsMrk0sjH2sG3tIHNifDWFP4A+epRJzPKVa8Me6LJ8nxyAgVbURr0VK8dIx
4H8e3LNkXc2y6scqpeS1E7njk9jqzsXu3oWfthrBqVLN2KiZqEGMsMedEeWJEM98SdFLf5w69Vnt
I7BnYA0Mko3uQYvRqp7dkYI3RlL1BTazteWPZpQIhAs1JYbFHH1fyb6domR/XUvauB2w9MUUvNea
1xqCZbgRQLbqgPoZBmZxyJhoj/smoGqm//eE6eUyjFXpMDb8SXtJB8ZsPyuDMxz/oOsQZsUu7XR8
3C2s5GWiJ0RVGhyBiCdBdPoJ1+BT/IF5nmZp0CijO7AgF6JrQtLl1/mto8qkBs1S6ya1lFDT0oeo
3kEfmYLhUfv85x3DCIb1n6TiNGBUdv3V51aVH/gaGBHYjKUJU0Q6fyrlwS2D9neQQ1zj0XgkIAtx
n6jExn3sDbpbAKGBbmX1K2ZLxiKIF3kPk5yDDFQO/+MRxQ8iUsLCaP7hQvdoYkmU0qqL04VBbV9r
9/Z4GJKITABOBw/oj6AkSkmwPbQKKWmZouwNh1jdHewA9/z+MsoP8EtG41e8mDHzP171Cy2uTSCe
sikLxQfCw2aB8mFoDxKaqoatrdpNOSBLQK2teYgR33Qmcr3tliKqfP/FqoLDVF3+EqcK2d+N+1RZ
+0jQwTtP5VB6E+2RAPiZbJ1dEcDrBdoVYzLqouXwiD2PK4SXLHSBnX8VoLJYoMvSGzrHZbcKlbsc
/+yNxBDODRRlqRGhJzret5P7Rcn8a0ysur1DSUp7f61Eg8WEdiM+hDCGFT+3ss6mVUf6GoJde/9+
3UN3KEWNEewArPJI5FFagJ6mc7Y+qO9+bQyVYERufvH+5K29dnLm5BYCYlBYWQLyc0lL/mlcn9+K
zwRUIgSh/TuYVwmtu/Jh17hno8eo8neGeLy49lubHG9BYWtHdYmOuQSDvqrDUpAY0055ncZ2vxdI
DEim0Koa+0MOhqbf2QtMIRDDRbFFk4ghxIhRQ1XYPeBC2woBeImZsMBiabVtL9Jazej/UTyPzVEL
N+sgYluBlTtL/dqesLuIrjcsNuHSV45YlpqPsj3CozGKuCYKMwFaU9pWCN4t7LYxuUVhKrneoXlX
lASd6L0vrd1uB8HIxDhCpGRENpGBkztEtvu0eUb6phZ4z+ujJgfKYLGKwtFX9dsYwmOEgTa5zvp5
AWIT973ykQ5C6E57vpsPt+rFhiR3okJ6YBruenjcqGpT7/gmLLuGNV3cKv5viK8BahyGC9CRhGAG
k2zGriFFcxLNFT+QI5ga2Jxppw074h318mdtBuqS1LYU5gbJ+KYbS2Ea967O1fyl2Z+7BIpBmAF6
7n/bClDTbMRAykgQWscu/44aAcar9W1LWK6NIx+8d0Axa+HqWnTdCdgSzuU3Fr8pRXlGM7SzwEBG
T3zh6azLBjxXHVaNbhsfjgKx1iGxrTX13AqPw4S2EJJytyQJyBYXGJ4cuOkVdW0G23I3I38H3Szq
tV8VilKgrP1U1r+iiWAFgpfqpKMQG3sAYr3S+y5yD1sdG3qKEwE+u6u1gah7b0vVoCjgPCmYoP3B
tEllO6LfGMQNd47/UqnK/M2B/wZDfPOxmZgbYnEnvYkLTrVbvfuEe5iJZD0nFJsa/dm5k21zYu2z
thInKbwTsoLfC9gxdfeTsG7eRjXJui7gfJibC3edTYub9lv9xswh6vqN0DisnkuZVw87MaI/N3SH
CyAAuSDuPdqPDF0aEaohkXmLTq3sMkkrrn8wo4HlYxVbbuuWhuNXQR0GPNoK0gx8P7b+7aswVgIy
3YCB4zShQv0wKFadMeg6BVuNsnuocsLZ4fPguL/Yzc7he3lrMwsLKO2Z8O8yqEwbmAqSgmzT8U3D
tYkOvvzMy0PxE/hTm5VFRHHsTlfUMqSPeXD2Zi35mj7KHgHz2oSVbNfudM/ob6hJWQFOHk0jbqMY
MaYWZgP/1k5EGFTs/TrGx1Iuxx0ZNPP/lZ7X/2MPFTIUMotPfhiXw3/1xe8PLmo6E+LKYxJc3aty
DqrastsEQ4TMxeFtbNViYWjc2hHT2tE0fABL/Y4uV187e5ymipRAzrbT/VHJbgT9qqg6ORNf9Ex8
hZMQ84y5p9aaueJq4XqUYddjqlKqlSogWaZa0azkMUuXxmfCLlVWOMlbXcNhl8ka6x85Flcmh6IF
u7QKmBjyaI93ofgezNV47BKc915YSHogEsK0nGcGGkvwNN1tI9kXZYE0REAJ179KrRMJRcGnFhO8
wkvNK7kA5wefEKLcWC1bGRwB3TmC5zA/s8zVeT0jJQT9gFg6HrcNs5hwF6/ZSODSOUVBybOpBjy7
K7SfiQ6jVrUdRIlA5XiPXthXpLcG2afNoND3KJH4bvy9sCrYjNvfVafbm7atPeLe9NhFheRbDMVn
G/hD4xhi/VZVi2xBr8N3m//3bxpPfXTi2dyRpXri4wzLcaS6blNT4G97ME970MxhHRYq+Ach2fOo
tzmi8jAWn4pUcNAB/CXHwGqRUIJthv6xvNQsCCWbJBJrAwFnIX4GZx3szOeT7GjTJ4mqKBNlf5rA
GUlC5ch/eehP4AkwFfXTtAz7y8pdALcsFbQKfnI/vAcMbcnEFbt2iewv9u11yaNv0HxfFy37veiL
VEKCDweO4m/nP0/QRibqD98nOIz3BPWwAwFgIHosnZ9FJp3WauYyR4WfHJFociH6pQn+N0fpsAeP
eh18p+WLvNxsSO9dJLL8kWyD1PfJu4thISe1Jaz+G3TQQGRBcouYPdlFhdEUHwSQ3cBxnXuYbTIO
lzmOuDDB+MZdRY1dz3/qYi6TCcFXag/bLhytvvV/OITfZnvaURMG7apVY2Wo0gsECN51LKpeaQYD
2QaLsiRcgXZhhBuVDkOTDnXmbPGFPEAcNSertmRANDdnWMZXzuBIPLCVpe4irfUjIM/Zw3osLSCj
kulp+RdZcYlciibnaBrD7gA2pkEzICEMxDYhMELQrb+l+4MmYOJcvgYHCgb0uVJu4VjK50RfNOML
b2rCCSCNxVxkX6pZChKRyOpydPBVZiufzmjiJK/sI7Y3F+6Z7yPwS7BBCHyQev+czRen450iqZEw
Bg5bLHbhRino4SfWPL2wZ9nNJ5XkLaSBg5rpI6Ond7Uah2sqw24ZQdJYZVzvGJpyL4nnTjgPGkuE
j7MAqg1EMPqXj8L6WNxoV2QsAcym6skVRXoAhm7XKGMrkZkhkE0/DW8oGLkkrVqVuPUa9zqcqEIv
MMNYcUhcmW2qSkRnGXn3c+ojR994y33YOHpQq1PAsP6zNgbl/zlHb6fSCzL096MDYg7sO4gwG1kT
FL7eAnuBEM01DYJtV89bJLyBeACt+Ow0Q/t9Ciadu4hEdiXFc34nzwhoUWeFkaUprrG9ssqKOwn3
zZCnfMSyop6UDbGrj7teTjOwE1nMBCjWmWjUD4RDDixUv5BPKrzraznDJcSfs6eLvEpLL0RcVTCA
5l5Ehf4H+s8tUZtxNbT0TYIcS05h53BlQ49v4P9yXyvRynnMmuOv4qWniviqPxn7YUliF9cVddy/
GYwV+U67M22OYfFNt+iRvJa9KZay1RYh0cg75nfAVNIyP4XB5ZdZPvclXfbnDiXDF76iHbHTjN9l
SxzJoTuzHVZlnJIb8NJN3mmG6Y3VEp4xMYLZvkdz4qiQZHsMsryFs/BaIU3Il5JOHgPTXYglgRcF
X/dY5kp7fSlG4eYZydjrd+gfaQwinGrKzEerhCHH0IyDyxK4R3Yk7WOCzhTNlgW+8EDZONFueBs6
KzyNenZckjuWECGDedJimOjVg6hBPbTI+TWF0i2rvW7cBuckUnIhGvagZ1sEfB5SJowangl1gByl
xy+xxlbZQnuokOSRSBYphjjheQjVyZvVleChzeRzjPE722uBQHvXV0MAUhmlxA5Kcpk10sTyfDDk
Z99DhSmT3SdrRWw0l98enhQV2bCN1P1su7UZRmewjoiIJANoDMlA1hmEtjIzK3QHGzOwxt6qYI4W
RpEU7JT4uAAv92fjlKZ8GGZkYItCIFe3B3nB28zgAUozJpQiKh/taxnFe09aXaCUJqttg2C3VEvp
fQOqeXMYE5r9osne4sJ4Hs4/xpOpmvX5Bop57qp9UJkX+GKsJb7Nq1acXViUSASvHpKjHVNF15Dc
qwxCW5buKNNGfH9mFxSgPrrqQ8OUgTCeQp0Arl0kfc0a+PITxFJXpN82akXU3zYuNfEUDR6zLOPw
VuShCiL5N4pGo6WzZzEOuk+viZ1oaspcgwXYdN7gYrVIMCxVapLBbnW8POWp17E7vUroN3xdq7h+
9+ScqunuzvzI5rs+mLibOj0gHu2knj0TKR2L0ut+NFe+RfmJ+2DbCWihFPhQwYAbp8+ePH+3GFAg
wGIljXBJ6DU2uD9qn0Wf7PKkjDPS8oFbt/U1oG4jdhsQIb9uo+9Mw8PxF+Ai1o5Of0PaL9XWlaai
tlGnn5NBEC5ICBjNlxKqoXws0m60jgesVQ8j9wbqal5Ls0L4l2GFs38cG8lvevK2gteQVQUEZZlC
t0QdcwNNbADWqI9Ul3HdRNeD3jR3pMUE9zor3LuAnWQl19t8cZcNYuANYEUasJsslPqkLpug03Y7
O987XG2JNL8zzhHQRN07IwsiOtCcWrkeNRoT+o1BMoV15v+VvUuZjw2cRnnCs6ZXNkTEyYlnB/zi
Ub5zYSaHgQTAuA/N7nA3AVnrnL3yM8HGEj9t8yQPktr8x4pZCcXtyLT1baDpe74Xr4ESQW+u6N+z
80CEQ89h5MDnCSyivN7geQK976FRelPPWy5adLIcsPtL7wzt6a6jiRCH+FvNVw2DASvmoHwOT4fO
ZPBYl9zAtlKnPUoWntxRVC76Gi9TQv0uFI69QlLPG1tlg0yfpKF31AcujloYCSvThODh/J5xJA9W
uDxwb1MHHjZciSTKTmLnWB9BouWz62J9EuGz07mU7/VamZZxx3qaAA/VQZJxw5lNNAUKrwx8LWYW
qI/NAIf9w+I97niRTjithh6kYBDzJY4j03GYomXQxiJEEprROv3ZVl6zr2G2L7oCnSMkrtWFcMsB
O0ir/OiOFCs9wRXqGpmUT4UPML5sdgomNylxs+fxsRlcFr20kB41i4koeGXkH0VS5Rlwv3ytAZ2e
jYvAD87H7HRIEy0fJAwKGidE25H1IUSlC/JT9Zolv1mOPjiQI216ig6txP+D6J6vNa67prdi+TNb
ZyYrdFVdfmsc8Yr8fseSI9B52SzxU6oavO5pK0G3kd5wI16112+qty4MdiZq/lieG4g5BCErSgPY
Yh0pWRDc41JOvwVzCXRoUdsvUXNDqeAl6Iv1uWlVi5GZ+Er2EHo7ku1KXheOmiwfZyrsOxhtjez5
4TE/6As77V0R7htTdb5A+e7PplwgCTNy7syokECwjNeGHCVfsQXWqYNCo7qHZiIeXlHE03YqUf6z
8UzRUzJHqFjukxuHp0xtp/xuKA5w6n60JcMDtnBWLDraBNOr+snezSG4IKpetW3q4i6j5kAoZk1T
HRJKbFTkIPP+/TNR/L37tgtWESwVUZ364nmEqOndr1erQk7LgzBnPdXX8QdCXDKSYyz9m54sCI2G
VeycEH9WxRCDxJi5bs08OqDwonJ+fD9bwVfgTsGJs+DfmXlkUPaI+CfG8wxYugILV2JjRo5hY6YO
bssgx87OOlWXLdj/ml1h/htIv0xa6DGOquiiyJ3WsNZ9oEJcy2RYb1RfZtUnysn3Wa8wIC4ShfAP
ip82Io6QSP3kaSxYpgEFP0m43S/6bDzwe12dowXZcbb7RrLXgYh0NX4z6UC0YTB0AaAcvhIlkSmn
wkwpU88KSOxkqL+MTXoWHzxFIPp3wgmnTpyJzU2alVFqljsDXIiUjV/TMUhEF0MfCD4K4WGhbwg6
zvJc31nhFBynNJrP5AFhgEUtIsH0velz6mqm9lYMomGit2psLJo2KHj2rNoKzriLow2LadgJUWYC
BB232MRXAvgFMzgImBNQ0PJmmbMn5Qs/hDpgVH0fYGNHACgWRUoUWVNe8W76i8F2fvn9CzsWs2hH
Ufq3JZucnXHKnow9zXelcf8aYmi15ibUlvyTT2YM8e/f9JtTx0hg1zU8ocI8j8d9rTF3orohaiMT
82Dis7DdXImSTRum43lvQsfsN8+eEZ3Y3aUCUDPO8qzoXNlxJg2Q8Lv76Oz87GIt8Z7jkYIpBhVj
Mz3uTaoXt68oWk518/Z+8L831VdWuXnNOYHoZx4T7Sn/ZrBwFNWXF2lwvGSNpyXLXuA00qR/zWBE
OBlLbXSmIFxAmAiUz4m3wnBLPdqNcVNtXMRu4ETJZJFhi6wtKoi14yTWMFzHV2IJAGHS7r4yCzIT
tzrsBSKafBYby7KeDX4Wx4ePBCLwXqin+jrMTTsnqczMcN33aZQ1fLIH48yY7Dyr+OMM2h8uNZLU
ZD4fra62T45Hg5/zJrHn1TJ6XGoNPmNuDLObtrChZVxtv294YZOp9VojYXzODNxAxdP8cOvJI0Su
e4yqI1iKoTiwD9qPYvkjCxWe92bC0GTybIiKySQi7ncV6ZUtaqROsXVi+Z1QCkwsLWtAJ45RIKJ0
LqIclYcKZyPcennJ1EzR0TwC+bvOfoWYHq95z36FdpCdv0EJqXsXLy8PtJoq/rTSLUq9qkZo5UmR
w30tN3fqUpeDT1LQvds1i+iZvdf1hf2FLYc+LlbXI7GaYDEzQCThobQYe69U3De6kLNbNKjjwhZ2
Usy0/oOJW2kY57VJWu0VRj8NlVJAK6eslZPXNbZ9gUYKPMdMmZo89x2OvFuAZKewzX+mAdESGo0v
/oGvG8M9eT6gILr/NC29AxiXkdk6E7i9gDEnlSAj+bwDvsehtYyW93jhfwxLTScwYW3lmpJSUruJ
7Q0Uu4hmuCTV7s1rh1pASO3CL+bDg8wKDQ4/uvwCs3WSizIsXOfW4KYKic/rkYVubOo6vOkjH+GJ
Tgid7jv8xsO+rLy7f9GhDxjN/PVgP7A9kuKpq4VV4p5DfOwO/keunvZwasxKWSCzMIJT/YcNm855
9KEvMca2vGLXbTwsLKFYWyXutveyRypyy4TRb2gPbmf7zMLdZtrFPPukSbvzNadBVm6eCBqE0dzW
uzyXlbnBHrLvPukbNeGTYtA2dkg0aUSFHex6uDOftXNR4aAA7rCjEEsmw9qzEnMQWIqeUgKKpsH5
GZ6WFxAuJIcs2ooU/TaBvHU+O8ppYgste0jdjOREjlSUkgVpF3PZm28d50rOtbMh+MwIJcj9Hapq
wKl40gIf1pbZZPyQr81K4AlYkUU5KRE4N87uMUv+9oCj3xqXg06CAflAnOUmB1NXWTOHXg12tVp4
htyS2xTLILILe18/OERPMcEEbjiriN/nlW82ALjjC3vy10KtOF2IcVOLIkmUNDUS4zUAlsiB9Ls+
oQZHdt9EvNC1rjXZ/ecyW9sUWlVacA4y8OUyDl5rvVmETwYcg09AwRYfIqZW0jVp8c3wkuyfwG+u
YNDQYejOUc6kh0AdEDEqcFlxtj080MwFHvjmdhkHbaaOMfpH/Cthv0CRteqV51jPZrYcvEsX8v89
FH2qt32WRppe41mgEnz6RTvE+XFGoWJGcsYKJl+i9qpunL1PNZJl+hQeH5MCjG8wtPVkskopFrM+
KVxu6kUOgT21jG1xmV2YTE0q3a/u1Uod/UBOLK+67oPBgy8SsJjgQ4l2EcrFSiHigh6mUAgnbmJV
fX9juIs+Bk3dtz4xQZqzqLRxbbavUtiycGzY0neDwAZLyQQhEz9cmPPp/rnQ2rG9zFjPKLVTCu8Q
GzXIPL+KMS4Z+99EdikESaQAoR69UohrJoF3GHBUC1WT/0L8E5yZAE/KTafFJ8Qu5xLQGWaSrsWZ
0ljMYoc2a/g95TYib3IVhQZIPZ1zEW1PZnIKTrMvQcMKXXRTRaykVuJgjQkPagt+T/18NPs7iz7s
X81jekTfyGFvQ/KbOPyrYKrQMtL3b3BD2SEUAfbpjQYFWb/61t7x8j6I0olFh07mZEQsPkfG/DSq
auLsFaLqOcLarPIKaU/WmH71pu+8Rmrrnij8cEFCNkRWcS6sTxVnaDwXJ6hZIhq1ohX8V2fdspEN
pOvJusVph7qOpj+z7ppb3Df67sg62ufP3apyjVgb8+6B88efQmjXROOWvatUiQqiPZXg1QjOAy79
+my/j53MGd0EU/sZXLZ3kIWKFnZF+W//lXUWECibmu40Qb4juW/U71VHsnGdjp13Pd+hTX9WSXfv
O8sIFrbvqoGeXZ3HxSoyEfWQFDQn2A9YUpGGL/z9b+e6+m2FP2barCFNeeF4eRoM6GwCpBDicCim
WCMTdkDWIdESh4wcF6kVoKfG7nLTDViK3uLjBuODnQd3OTUYB3PgY4k1vHY/dgiHUNErobIOZW03
b4pC8c5ct/U6PLup0vqiDSTu83Hmw4fODw0+q+t//4lGjiUQ+yxgrzOqDEGH+iVWYaieH0hSWebw
MGzvO/7s+3pNub7i7pbBud0IWUsaPOMkP70mFYUkYfkvrtn/k/Q3NqjxZGcJ3gBngBdjkW8Mrh/H
zcNCeLulteJ25yPFyyvecPk6ZaVanUAzugm3Cxp2z9fR/sfbm/ZCoxv+RMVm8CNzMAhuj2jKZNj0
jl9wBwFNHyhed5wx/AQGmmdNpyJHE7f1Jnu2Dc6uRfVoxLxCp2TVYRxF0RCoKQEYVhchH1HDOBrL
lwsDKRRJev8Y1pkUwO+VhrDBCcfC6F9atzR1pVpAYRNzDcg16VnJ1yEhOeN7pA+1ScWUkgSS0BdE
/pEG+u3uBbOKRh99+xci4cuTNnp1NM+0OlM34CvpA5KVFlEXse7L+kC6kYcQbSu3YA3KK7JqeKRg
nTRw8CRiyt5CIk+TuyC+HnmTqGLOqLC2rwkx3Aun+2oc9/+6B4OAcB7tWmIUj1/VkF7WH6VXNJub
bFuSlATHd4GythewLU3542j5CELYJECHkXPTjnKO6397eZd/+ZKQI/OzHpRw9/HeFlmooPrbOUDL
1XuGStrLFy+M5WSR2Em9mar86sqy3qc3fsjvGm43AO7Q/hTqThnTMjwnkjXTFVatXBrcj1vdgBYz
+iLusdbPE5ggGpAYfh/2F63BBu5awfq1NAzjygGa4J5Ard0splQZN1P0zFlCUB4nbDsXatfYlS1O
icmfsrGPNmiyx6wQI7Nj/vyhf1N3sshLvW5mPEwzGc7W5sJPGKGXYiSQFUrCVqx0pXW5m6xOq1DE
3jec9lJF5JGCP9h0zM5xgZ6VzS5tlbCyTeIg9dFPY6wsgFez017QbvR+r6gYn0RGBLe24PrAHPUp
xKJsqqwne2O9ssMedUZrjeygg1Q8bQLuY2y/qrL+V5T+mDOX/KTfcol7FBGGiTko6a32aivcUoFz
q2wA1z9WjZTwe5D6jHgLAGcyeVGA8s5lBkYF/dDrcWJb5dA7p4A7bbx1e2J38g5Ic2g2wEo7zMIz
6bgYlgy0WUoo8nqClgpk5bwPecqXCx4+tlgvVhvQTtZ+8B6yd743OtEwXBGynbwENf8aIkj4Zm40
X5X4hKqIZ4O+nDO7yJ8BNVx3+g/5ukI4behDP1coxlVYQoz3VjjL0vv2DcsfIGVl9MfgoSz1399x
lsPNFKFA/Jh1JgiqdMqTBQq9waXUTt/U0tuzx7UpFx568ODcnuU1nQD+jJBRQchGPapLGmjmPH7p
c2IXAhfC/6bCAsFilvK2VfK/ZqWHrQmqV1YKQMxXkiWeeVTm9WaK2TEMKlarMOShC1zfLkMMTPPf
FALZogJ208Juup+sFl3uNJ6Amc9Fg2dm/dNUdPt0YowHQn0EveTsIWBKHkU6mcaVaEGXoI++05LN
eJcRSQIyIR79dh/TYVQoo4zj/ooWKlyRorm1JbkFFiHRgIrrXSNNbVUEdDn3mW/9zI9wIXoFfVt4
UCnXxzVYaPqxo0dKVKu9mNh+gs3SrZtzfmdo1fBuTwDNGi7iZ3RuCWWRZz8xopI9G3Ax181W2MuJ
v1BlW/HyAszmFSDweiEF1HERYhd30Le4QxlR6kg8niLipCTUiftNdugZz9BvjBm0PM8vVS/2wFM6
uSQZ9uY6hQ7qUJ2jcpz+NpLrTHCQ9IBrcTyDiDQNadZyEOGBYI4E/ojLRF0chmIMuO4bvmUVOFAq
Dk9/3wghbJehhXQGBoFVJ8tOfRdMJq+rx3T9saoAZ5uI6mw5NWPiqTf/9FV5ZZL69SCB0FTRWxHR
sBK6IqRqUcpv0B6liAtkj5nNPMHvIdyEy69mQOyFCSrO4MUGfnLYTZlJZUHoggaViNuE4voe+YEV
/EWOhqAEAsjlzHNRgT0CyRy7+4gM3k9AwD1gPindY+Oej5UhrhMucoRllfuTBmmoEpC6uB4dI7gD
WfDrYORlryLW2FnSzD6dIQOvqTcEb3WDD2kEc4zHBG76W91jQW6mQUr2MCJWKckKvu+xKEi3a5nP
3H9SNEhkModm/ocyC9SPBOpRlVjqxCDW2TVtWbdRnqLJL284dD/6ev15X92xxKH0tYshENZGJQGF
QrOvQXQP8k+PdOv8+KErn9xU4/ArtrbA+1DKC3F2GA+vh7SBxnfaXpGfmcsf/C+2J/XfU7OG2Onj
GF1D3sPc92dumxL1T50piTk5128U31RnMhwHi1OH6+1uVrRvMBafVlQ+2CfnHI+kD2yEqheEjYhq
GrTjUFm+ehVVdvxqbVMJUw9AE8hzzOVQ10zja8OMpwmYhTb3jZCBAGrPOJQZ+402EnWyFdYMKvZT
nZYJ5lJyuOmu/5iPhGvq7Nyxm6SACkIbbrEmSNQCxmwbYPd84WhY9YyehkcCFiAyxGRgVmRTRdSr
eQO0v6pw7t3B8k0W9DZOoPay2gpvN6H93U++yAWN07nhPaISCvzycK6GGk+1lODmbSdPJu/Vx2Oh
IAoyenjuImEMUF/NhziJp09rtTBeR/fG7loEPj6NYr/KabECRbdT8r7B1AmjOJFKpisPLNXH8eA8
XSYQiy1OQipNIlPLyasf1zEIlw5bCxXSOBKBQaWuXcIrz4b43yNMX+CtM8UZqmiXAGDJRWLKNqWH
Ki6pOR9v0ouyr6T6lLnzizFJgNYkW1UH/j5l0Rko+U63zHzO4+kwbyi9e8qZZmAqMYR8k+XvSQsh
u767pgKnMYPozzWMQCXSO8z6UlvbuP2Yz2x2vJmC0wnpGdFQ6jh5oUuLFMN/z2KDdvHrWRfeDWKE
OBNK07izDZDnMoEOOQQdB5O0yNus+2/g14n0o/L+86C4NMG5Gzw7+ka9oEQ28qF5AhOyBfRbbsoO
FtyVDSjfnyZERNZRARCLbf/78aLoopqgRgeePNOC5EMlQ2yGI+EWqvksSxp3vnhpHEFigLZuMMkF
kQ3L0VsPoDTbukA9EHskk8BaPA6fHWUPzOCT0y//nSMC12lfRK6PpIbWzO6PF8TivUOUnu3rGQ2q
Lh2CNSGfBtQMuQBISY52vVJs0GlSR+FvgmOpgckFVmwtc07ySo5Orga+m0zZXMrF/0E9POplgM3z
3eKsBtPczTXn3GA/0fPXEo1E/mZnGFJZb8hSpkHNeIo71WEZidoh/mFXoDETGEEbEvfTcpRhRj4k
r7f+pGvOauK5us5iEJagbn6CgtnaslYzX4bo0AWo7kEUqBVBRkjDJxmnO57PLdPEVYelLEVFE9w0
SiQsebrbMlFEJSJBWAgsFPaMlbIVIIvTPZYNepTEs7+WYgQXqPXO7KkdfT9uALbEU3P+ivkKN2gN
FxphHsa7MkuluBeckY6qUJXgCF7KSaB0w5AyZuaxQljQd/4Cir1xYefex5yeCeOrRBXxBfhZ0C9e
LKw/9abcEa+QXrfdoPVoKSWv15JbuIvQGX0I8jSH6OFa5ogoGWaenakB9n+YKaTBotjVf967al9z
/SfdZLWAh+N+POJK+zsYyyHm2gqVf+GJ5+ljDpJabNvPp8lNMlc9MeKlik4wPefSU2lsJZ8/ZO44
fj1jBg2gwxTjm7I+5eePbJ1ejIfOulKMXJ3D1EPD4NwH7xGh+XqTsazMO0V7eSKRCafZQq7YjS1r
6YF2bpaUMiZptAQIwdO0tiOxxAvG3hOjWQcZncaRRwZjYVRilUaYpeudqaec+xlMEfXfOHDIH1bQ
lUWradWP69j7d/EpeNUXaRnDj8SRmQj410taxzwjG1Z99WyL4BaEJqEnx0AZL2jlYxVsVzaDBt27
kub4F12PUUKWOFYE8vFtaOOf77LZmf5kuOQWa4YJBUunutUoK6qs24/yVbv9Sa7HCkvUQ97toaiP
DUGJnZt9jSXCjcSmYTgxJR+E3JWbGpqvvldOy3e3SvwRqa7LZHjbJXDWUbvQIsi391Rlg59j3fOj
VReCDUz1NDMAyvj7AEQ8irO/h8RcryWtlfkO0a3WV0WD7sj6Ctwf9ApoJ0ttGjR3gj7S19lMOa1u
n4Sz4jgDj+z4rSfotHP7nk6Jxt+7Dx2Las5VGSU5v4ynuVMJYgLAYz26vbzt6G52P2U8ZfEVLwco
AhnubjcCWCBI7lcH1iHYzcJe4ohWaooBJog2wehzYhKHm9jhxGUjxlLFb+OinjCiIvaMTthpTKzD
StYLMZSwSctwZfp1+09AGXSaEYyp3PAQvAtglZCTkyMm2xAf5RJ9MJDmwbrJJsJ+CqhRnZg8PfeS
hVEEviVxuVqcf/DdB+8mZsTx16KXootoa1fRa2OYrlvRjA/PmzNoJI5VNKLBomyG0RZ539Zxwqsf
JNZoeIvdTC2Yp6D9GCP+yLshl4s4p1sPpU1JAlUuFiAczY/+ezSlj21MuDdURlm66sIw8de/z8P4
N9sdsNf0Ka7Vx1PYIUj7l3j8dROYUsvrEww5azpzjFuAH8a37tlQIb1w1qeEDZHymN97COeSYdB9
atf28tBLD1kpOj3vwsVrDJ9mWWnosUYBLqjcMFj7JxgskD496cRLuKtAN/HdmVvZK5qieq4WbeAv
tLBylwdHUlzLj0znu+1Emed3MyDUpBuDcV0W+KJClOPHtdEQ9NiKCKBOJF6OJg3B2x6VKzpeQ9DC
9xkkerRYbYv+PwjFv9YIXY6Qhk8dbcEGJhJpsMiOpKERWdcS7LWOy5JyiNUdf4Aj4+oOHCu4t2YF
kAkYq4bvWJ8KIlpYUcM9773+3a3Fpw8mqaO8E3n9/YXkmDoSmyAmauXsb6BCce2a9q4j4Yc5nno6
IZt4LxFuY7EFV0XATYXyhz0OW7h2AABqU31oN7TZIS3+dcC0Ohols747H/CRvF+G9TzZ5M2lGImC
a5OfFq+BTwbekxsGZNhaDRQMucDKYARjuVl+rRiH+gqDE8yPerpWZfOIkzW63wVBNq9e/NiTQKPm
Yv127oMe7l9hujyI08Vf77Qltlo1B2g+xkJa5ABlS0qqALfLP5iIBrdW99Fzm8miFliD9VgbHDRs
9wMyCetMKOWLM+BT0SYIvfyeJXN04zM5a9BYwGB+7OFx+d3t7MlrzvyMdDP3MAbzrq0tkl9GUpeo
MduYKh5mizQfXPMrdGCcuUUmi6XCK/+ia4DH61qk/K4HQ9gaDNM4HUkXjqAcXQdbWkGmjh4NdQeS
+wmAPO7u/b4dL6xEPgumjrC93hiEBiVyha2USo4Q+hzVl8ni/WURryj2Go1bMMjWovJ/tbCZJAJp
t811OIeyG7awe40IyrT8WooRkOodhQPtU4TKhQUTh5hlyqeA3EwxCCTmuLo6wJJhIMYV6jD4B8fe
ll8uOxo3KLFjL+/6R9n/D5VCX4K+ntlHdJYVYKIENHAnDH4mwy9Isosro/vMJq9zOpvBGX1NFxer
6YMjvDkc7QBHAWZ8u1BJVRz/mYi+gdO/+LMNKL60MO7JBeucROQ01/wYVYAgtcz+m4rHFHeHJ/xm
iFxFIVXf7wUaWNZbJMf/iqrHxCiVkS1TC5jq0c7O/UQZWa0xXHUsULVenGYRgFqrcoO+FxsJkoAc
G5ex/kqdDstg6UKSEaNHhLQU9MvHPcpYBxzA1UPfpRVlWwUWfCYKCGtVA8JV2/OEfPuTBvpDuuah
vgaI/wcHVT88A9PGSwdhVyg6bLROjGc9Va6Drz0/0YPPDTMXBj+z3/D8pzCvuekFXBHXDjkvEzeM
jZhlQizd1rVS1pWd8AQi/VyIe3aDbPpdzWw0w9c/K480r0TbUXNvfChxQ3QzUyDvU1dT3Zh1a25L
70SNssZNJY9HrB00KibSrnCpPJG4EhGGYFh4WKT5MQd7Xf2DqZm8wGfEQ/5o98zba1PNfx/w4Efr
VUsghKl40keacRW2qfBHkBKAScHdQ//xz2yeFMoX3ZkBEhZ8fcSiQqBHmzbT6yfKhzJtv5YSUcFj
IEGCglRc+eO7MB1XFQeridD5BnRhPfwbjXdnbseynGOI34ZC45N/3sijjZUvf3OEwO2z4/uFeGUK
jC9Kk5Xf/D4dkr2IiFWRMnmg+TGfySOs9eQJEMJrXTPybnHBSOfy6HrOpkyWu1xLD+IrBsTzC6x0
V5T6io20aDYpmfhMYm0pzOKJbCOvM3omnJpX0SvoDIZ+VFyv2k0wFYVxBtIGl3IUFxT2bnpTFy3v
ZRDOsiV9JySo+qWeanvomL3xqlVjn3UlzKlMGTuP6VR3+3HG0j5XVx8yGdhTbbotNkVmULH2dPxR
0VOylOU4Wu++JFtQhmrQkL38KS0kI9XxmJhXZGV1yqWFdnY4SrUWNwZY1tkL6Z5XPZIV74P5GmCZ
VCEj7qDMycJ4I474iJnb3m5QToOvZYzV24D+k/+VmD/oi0Kdn1e6dbooIhLC7TAXPHiQj+jK9JFk
aMpFZ2kznVdiQ25lmTuV66UGOROPVoZGgVvEUl6X0YKpeXkb/I4lED0wLsNmiEKz89wmM1wXzY1/
5WepjlYWcAQsSGpK/UgqHMfBJps8UAIuNJDEFMxntUuBHr+DeEXMALbiOIhn4n9myeia/AwmMyWb
t3/WkbQNNIsmv2Cawz+6Tdklv+OrAC0B2eUNLP9yMMxyILoyJEnqFVKPnvKbN+tSBwGRjmtbXeTt
tEjb2GS+gHuqgdNS9W2MbPhOIVT/Q4OmWWRe/tfadMhc2ySY/TgqEiCkeLZ2WsdrZS1Z8kTUAq8E
4tPxXRdSEEgSmpTW4zeAa2r7ftOUTVs2NGDHjwzinZrJqT5lEKO3pzjyEerxRp0ZAbcMD6xpND60
85OtgposrkXCl6MGRnQPyjUigg+a76AsXxe4anowFuALUcK1Xxj60WrthsTTpdjrdchVHIvJiZRD
rjdoTADStU79sHV6H9X15cG7NB4/wj32plVYvndLCB8cfbCxBONIGpPTQgWXU0aeD3Vo1b6KfIMk
wnGSeTqORlkok8cspxyBZCdp9rnowvU7YVfaHbWTHCdvyKCehzEAGbJKuBC6xI0CiddhOQBLAjxR
wuQEo9katfHwJqEm8Na6DGiEnZUUEp2Ul8OW+cruRY+iT8YVnjiu8x8Q4vZlOYH3xMXSdhyRk9WP
mTv5+xxQd6aax31tatARVOWHfjuG2J/dUzcjt1UQgHYkTp3gHkRAsZj2x0FZaEEUKmgYx56wSrGM
JE/53r3O/3AQMb1+6ZwmY6MqlaEGZ6vzpWTrdvvEAILKsJlJNoosxpV3yZkukSXTwdSZFOsJKMOz
hsQ1vJcWEEysQFUrN9F6AKwPqH/Tf1hMt4lI/48+h9iNmmMAuZMwi4zqbX5tYAFAkyhXbEKMxvoK
Ty9hlKiKTYERpxenqXsKt3QklARtODCHESih4txSh5mGfe2sltMUjZQlBI9qU2dZTt8x0YB/QUnT
uPcOchBuWW7kQX0kpJPnu2b3cedG3Hd2bPOIHD5XRlI7jHwGihiPVTvPVvS2QYaFkZb9ti8/qP6a
q+NcWrI7qQbnAOQ7MjvrGy7KDATgJQ4BuxX/d+RV+3bfbCmrHC91vnJBqzm4KECrucuCRO2oxysC
gLeHS3HVf0Rh+RmHBN5iG+fZ9JLf7LIHVXoqUMDO3yF+J8M0Q34lk1bhxgXW8CSd0U//15SmSH5/
onwWZBxp5SMWh6IwnfRxouTS+IFgLKz+XxhL7T9DHWTebLjHtm3LsDVY6QUFmMspEsLovMWWcWjp
G9oHpOISR/0iHYh5EDq3IzB1yMp/VPKMa7m2b/cgwVpzP7z9hGRqD17p/zOjxw9vIyn07vxv3xc1
ZFyxFUXZ1IGrmH7OxMooutC39LjqbGlutBj4G2YPq20LTuzCmncxTS0Mt5nH9ohAGOzt07MeHpqA
sM8zRHNDKyjXvygVemIYIGZRqfkM377vGXo2XLHY2WhJhz3eTygZR2JBH4pTnhjMbDwBTUCqesKB
/k+ruliLRNPK5QsxH0BC2U57kQu0cgoFsBKXo7dV3h/TUSklh3RsZ3HSZL71IaNs41ZpwpWdgNV6
gctyO+cLW02LXwHHukwB+iHw79AtCnZ115fPCZqIl1eLWQbvyIkfJOw1wlROS4YZHf2uRM4NViy5
2sMQWaINlLgbxn3s0GRUE1im3+FDuXQNbE8SN8A68s2CY8bUTBcLJolrz8BGdC4x2nUYU1qylv9H
HQks83TmVFRBmJeYGtoVrd1MbyukJ8GOka+0rW1FyJJPUVBdUK+51qhQAigBQv21BMqFAfm140gs
3oyCUEm1xTpImzbkAJ1uth2BR/fDMrS5mNYC8CgQQrvfM67kyh8DWpFUlR6LBdhTzIrxdg3H4ziq
fufwxDgszcU0xwnXx6On7xkSC+Mz84vXnwgmnG1MLJMF1Ic3SirRPBhE/9nB2mZHCrpe3cO8E+az
zEsjXK1ehy7baQC/sevGn9l+UYxZ0F1j1/tpOIPXdr2RhMbycvQ6iXiPRjMPX7cHxWe9oEebw3dU
bltAOoZQf5RPcqv3tDgN5o8kKjuiCPtL/nZxZ3XlWkVTkkXqvoC592om3ROVakRc4u1dkUyD12HU
yAwKJegCc68jU4fuAeu7cb68f1VrFJc0bQpP1vWfJm1Gz9b3IoqC1Ai0LZLr4x+wBGCCsg+J05gB
n7ny91mUkE8YAU2cpaeq3Kqwr1wTVizd9KdNZKspON6Te5Tg9F6beUffkLNueFL8Iwdz0l2NJzev
Q+UccI0R7VFOvonrgr3w0+Mq4ZvYZgAX08LNwisTuFVdWv2KIBYdD22ey2ER6bocX8MthXwyriyW
kOkBdGeUWtD04uuiKBlexdfRWNQx6HgYWSwoHxSA2/UQZS8SLwLhKd8a7a+nRyEYyAbKMBGoRVTb
7hYnm8p6oyBOgVUzIty9m/kn9IXZXBFhE137ykmgzulOrhzhNHBbnsbKwq0Y/PDp2fnqZmOiFXGY
3RuBvR00SbarDgs/4PalGYESyKH9jUcO2D3rQ3vPdP0TYTnQAQrU7xrw+tLjw2e7uik3INedJsbJ
XZH4dWf5P99yP62TT1ljkDAygGLLaNJ8QzSsUgkOo7YLFt5gdxmYmejd1IJpvGK94QmKP8kN4sKE
DxaV2QWbYNVgx5p/xa4mpdc5M8d6nGKe1pBR9VlmTEyxmXfrj9DCaGUL4DthQp+C8uz03qPvtFsB
+MdiBLyzWVNtguh1JGjgbdNWfKG8+oaEqFxQ5h5UuuddC2XJt4TOqHx6dHwkDpoRr849pmBdFyTe
x7jtoqCktiS8uwBB57wL6jycULjXWyf/aTSc3e12wAMznwg87Th5fOATpMo1E5gQNmw1X7zk9ykt
+jjyga5fBmnRvxLRNYzBBwfyhCMnoRCNRH5YLx/Hq6F3uZm/z701f6vxLcO4qr1IvnYpZ6ecN2K3
oh174RIBh7GL9bQCsKVvWlTNr8oB1cItfTd4K6JVQf3YY3kal528rOws2J1o3jBNlH2RTs5JFdNE
vkIrkarEG7+VUjR98CVVNDGpnI7gKatH0kOpM90ZdQL/bab0Zh/b7zp5TNQWBn4HOT7s3V/atl1V
PXANaHA30l7IIH5WKetCX8mASfS8OuHb3RjFFaPhJSJ4hh9w8cBcKyNNjIFOYg2+kI0Buwzj3W3l
I6kCwNzZi2g7+lH2tr5T1gBHnrtrN1on7yvvP6pTUqKhnmxm04g8vF/OYlGva3lC97VXDpYx95lX
frAdT1EEshF2hg0JPdX+RQ6XWJpCKGR4FA6AK30Zecf37h1/TG0Eb7fNI7INWBRl/bKFaDR3FHfH
TqCSodNK0Kmmbna3QR9aor5U4ws8yr7yIbjbm589tRNpUsW1GG40kqKmwiCoMLciQ0NTU5fm8sx8
+xDvq0DsSmMkaWUVqek/8YMn2HJQJFuK7yEmLfR1CpEW7M+IMb3tNqxC5/tXJi0L6on+GBmQe2yy
AET2tx3Zv5+isY4X3Jd+2Fky1IRV5RHLhhqjMg8hGE8gz94ZnJ4vF5zGl8XPtySibW/7e87jhAEn
BfT/WmmZfMAPVrJwOKfRFmjK3zpJDfu+Q+b9bGBLLE5McirSZmp7qGlR0j9ODRdDzmuvsFJ2y1/U
DbVniaTuYt3Gxs/xy6q8fHT2+QbqwlxfVyFilpjxrSPjZwQcSU8b1IDtes+e3id3DvI4Ij2IdPqd
vYPng/QAkcJ5oPAODZ0wTas29dAvfw6E4EAyGdvjmlDf22LbHSMee3OR92c5g5oipRkyDKDyIOBH
39K59o2BYGVmXozMp69Vf5Xe7AfUHvrsLePh1hwVpPcm19YVOoUYRBJ4w/6wTdyu7/SvELcEwUwT
cN79Hmr+EifBPK50z9cMJxYyCObUN6DXEmCpanIfHux5XdQxVOPUH5dP5Wxsc+Z8thdqsGPcttHF
OsQkQSdVw48HpwmgTzzXwAGYlYNXT5/Dsav7cC/o2NzGejPslREmGb8LfEsWZPB0n8FOkVhlzsx/
KVa0S1uTVCIA70XkCj5mE+MJNLjdlEFQ/Y5WEDTr8syfkXHCyBfI/aE7lwC6ZziZF/dHuvpJnhzK
856vGnXLqAYbtRNnjlxRSTfRIeWoIN7yk6SXpNSifaXS/Os/pPRnT3f2t3SLwQTS/d4+jY0Vf2PI
S4/JvRFR99AUWq7KdwE+AtLaF7lRTEuA3428VQTHbDyWLHi4tdZZndInxUQUulOi8axG7UsSAVBm
kA2wJ6rv1Y9ym3Kxo+bXhq4NOG5F0I74jbexBZeUlO1YCUe6azMc9dHuALt/bJhNcvEmyW5mCcCr
OIKFoQ059vMnhY06Rwcr3ezRKXgfjGToLdAW0+9qg3Sl/FJqbs4L4nBltWEK8b2GcuFuHsbAgsJI
hxKMFp9zuwFyyvsyp1WTz2eqXWk19F/2VV1TmAKrLzjwkHSpAjwkSrUbnyp/IdyFsWg2iYYaZ2HR
Sg6uRgja0cZDgsk0Krko26dUOKUc/eV47ryVJx7QSGM5QmUq1uF2cimojlDiWiFLfI4q/MnMc32N
grHfJxm6DGHKVeFfDYP909pfcFvczfkxJ2DEKnX94zkkXEaQK06rjObu34lw/c6JQ5Z4t+58r1qg
FKt2m8kedlHoNRdLb+uDAttm0xlQA+0ESR6VOVZqS06TP9rZmvNuZAN/1mGpFAP7tEvxmVE7S09u
mURFrKLIvEGjZx4N1X/PSrL/wlgJkds41AM1v0mY+IkTrBPyit+iJOeE7PERoPcfKSFK7go9Yop0
m4kOx/J0pfwoK48witEXeKOb/AIDfNHL5iifF7Ec4z8OlTb5VdWqmUfT/ZYnprj8F4VtliNfT5oz
wM3OZ8lvrAFRNeeTNyIVF/NllqhUuYKHiIprFFzSSsHPMSeZbpaDCe99TCRzgoEAbqlj16xYhCsY
iFuI8zjHvgL8n9rZ8bevj/f97DE9tv9SV2OsW7prQlSPajhaiKbB84Us4ldZiR8+fi2n5c0g8zBS
CFqWkZhg9W78WhunDbwytc5Vhxrp+ivvmisInia9Bq/02/w9Tm8APc0vtPNTdf7b/rQ43Jj/vMWj
dJm4IiRchPWWAszDtCajS8jyw8sPu5s2vxgeRLBUm51QnAc8zrT+94rB0u4GCdyJNQjdfqS5gyEw
/sp4M97Mr2LbxEgWyD5W0y5U8KMDQ7BH21JaW3iLmyk1rnHf+zc1JIG1iBuSgbffNfbwKWEyKP9s
zlAmZ4YuBjMqr/rG/OAiDDv9jmPpt1Et3KIAGXWkLFutxw2J8imCYfbmtWrX+8sY6wTUbFXfBQbT
cMqo7LljTjckyTCFRuZvWFU/YSKcmx5NrqlNLxhDIQ86m9/7zQz2bXOwkk43zWSJ13+u5w2u1V1H
pkzNnyTP5LEDg1nxo7NzIb70CPA8sRglywjEkl093BWW3SS7wAiGWbQ16iJrKtI6HZTG1QcSTh5R
yQO/xi9V7ODVwQEp8xAOPpcXHsAOTPIk+xe90vN5ReMX+3npqjxhOoGkdvkbDfPCyLXQzCCF8Awe
VFBrUw8YmcP0G1NJlr9QTkqFNIWYUZkV0f/8gNvaGS057KniO8DsuzrBt3sCyU0p9JyCmcQF1Igh
GjwWxXWcRUsXRIDicCapLufMATmd09/jskwlhM9L8w5CSPcDXL0ph6qGSvU+oKKIVIAD7a7SmhxN
B7VnI249lnOCtRjyGxzyN+0OG6d+rgLps2cfcZFWx6bWztDd8fMNxrnQiaND7Zr76El43r6hw1Pr
fMkTOpo+r4SWoAVRR7T7Unq5nAi1ocuSeeADelGdQ/bSuX71yNRzn4uOU6s/fc9cL/0p0ZBHvxGx
7TTQux+bhf6YujBApcVJdN2s0jVK4GE0qKtmRYLNeV7nBmXMiSfqjDCB19FFtQZIkW0ge8WRdCqQ
IduqtAa6q+vTKZGkNheuVmkk6ytGpb142Oz6aLzDRddzqS/3+LG3ogXyesMH8UvzHB5d8Zj/3yRI
IE24eMaHFo2FfIr7MojGojnQs1ImWv418XoXc/vTztLz6I4qlMqjuzfI+gsWh9SMpZMn7LcsdLDx
jX/fuRrs5zyepWZd92JJnKwn4Yrk1u/bDnlPLHD296b0I8BA3e2xG6hHgjThfiWLdm3LGCThijRm
sAIU4sVEkCIQmUkw2dwNJkPGlO3Vzc8KYMhCSyQ8Z/LPRATuCog7dIotDyV4+/jOtGxT8vxNCthm
Yzmsnpd/i1kONB3E7dXnaY88lm2Yf2kj/AJefBkN8I9kGVZC2SP5pkHMtmp2VjhvO0hzT2fsAZYC
tPjkpQPmJYgAOU/tafo6EkQ5QdYhAzITjSS6vvvAnIj6RSOHvlgxJspO84ogE7mOrnnquS/peBvq
IblCk2mVVAg9QO0mJwn9nNSBKcZqPxK/twp34WhtvXvYcwqItnU+Tvb9DUHMKZA4F9F9dpagUhdk
0j2PxJX2iQsjYlY+wrdbODxBxCVsOd6x0gldO5P93bFQ5Aoh3wjH2cLWScCl/mKWg5LLRrtff32l
VFM3EoqD7P4waw9WXiS6EFpJmz0o0iZFhbq9u2EllmPbfLefcD6DATO/Yw7A/aH0qRU6bG3MLy4b
GlZjwsb+lomXKibmUIBYPYF8mRcJFO8iWQ01nC0HMZgPrnPjjiPamzuSbqdk/5cANCmgOURO8qZN
SjSjW11x6XDYuRD5/AIdnY5uPXwls1ydMoaC1QMAqDOaCqCxQPjtrjUCeEhdww89C4D473HIz3kc
+Yr0vW6+Y646AptVrCNApaYCIQSmIssh0nJaH3Q9OP5e3+aXsWF1ADeVUA+Fum4XZx/VDyMN/Sh8
0yadlQBtnkW9og/RYZLzT6pSMqgdHFfbrLTyuGzJdKTvKftkPipuxNzUPwgLVJ/8rFClBCsyqmZM
pz36y+oM2FmpLM+NVal1EvbULFs7wFJ2yfROWnDtCwz//yKnDWQ3AiuJVeu4x6COEqkGGawxvu+0
kiGuuYq5peORSSJnEliGz03inP0Ifu/YtTs7B5fn3RpucLLU4gdgARvghiQk54fQ/Vv5Kjt6vO7q
cJiOCT1+DA20KUiWDxhEooGMF1g5bmi7Gq/pLc/YXFyY68MtrMmDbp/92Fiw3aTrMLLhjmZaX4Xu
3/xnwmNIgcG6DPTMQCe6Mhyl+IrLUh9cXU2aHzjUaVVtF10plF1NPIgRy3YUt5yhu5K1pr1HXVSk
TLSImtXfnIdwpZUxouKR9r6BdPfswGlFbX9mDS3W+gEQ6pF2S/UmbyOsPkZC5EoZZBZZ0+LWs2xA
KFLxDB7NU5wR58Pu1nPTYUL9kdN4sqn8/daDNpqAP201JjWeJ/jgE5YlyL8occON1QdlgjlY+Uy1
RkWZLJ3QIcU3N20ii6lTrLY4lHRnH2FQTd9VzNXZIgxv9cM8lfrQ3bxy9U0sqLoEJPozHbyZR+d3
zv3JlQlddgv3UyavSqfr6CSRQtScuGI0KiOmgIdvnfMv4H0KC3wBIkkyxCYef2nUegXakY/OdtEj
fOUSOhNifTs6QunZnB+EI734TWKwzPOPm2Y2D90ysGQkwHVISTr25xoajc0DJQr+JySIoPGH8EMb
FtXl1fGgivepuiCeKvlY1PQR/h0d5ZicCZgebXuQmi6wogb5LbeYPgjJCOCDsnSxU2xXVCthiAaP
sTM7iyUvkprp3KFyCCbU+T0Yf5OjOJMkl3LXIPJCxpEVu8se1gjWRu16bOqWac82Thq5zj2MMXrg
pJfjC16S/oku0cZJgxgd5I+H20UTvBf+demS5qtvSSy+tR9QBQlt7FrFZl9W4MOtxSvE5AhK7c6u
cZ6QS6zYrvzyWK9XVhOoZpfLUkaEyI1rUE8mGEwuE820wV/ipNHRX5ym+QYt+eFMoRESMdt1TFlQ
lLB0Dcpe/Wip8jSK6rKjdLTE4A5AhJbZUbolHhvJsw0jlZJOenpUGaDsHzBS5+x3myRspbtsuO/A
yDwnZWXYMAuMe4ViqMu9GgZoWUATho1/0hXwCfZ+jVk6hQH29WXYkPfQaAjJ9gQ6v91mtWNr3FFV
8ukL1g3UcMeV0KVUhkYc5X6STA81N3xTQ28mMe7EBLC26rGNvR+Ai3l9Y09bpKtmVZTDJ5blEE75
N6+tWUNyQDQd5yW9OEugo5e5FrpKlj5WrNJqYjMUt2nAKEMaD6xT/tTYFdhPS01YVZ4luAzDb4HA
vDC2FvwE5tLWcYmCKDsIZlwzTZohvds5pkfSaZ+HJsJLo74JDs81U05G4SMlQ22q2rpN+i6vqR0Q
6FkkSBHwNmk0mwaq+rPRSGHcsGuW+274pZxHDVCSkGQRINCP9nffvXIwJyuIJ0vGP6UQ674PXNOB
yrL21Rn6fcyBziH8FtgLLj7OF6D/9WUNIz6nAJlzrsy+78KHiTgczZRhh5n43XDHwGMErVh1t2l3
cz93hD2rXvqe5cZiteb1lik3PSCjhn0hsHj3dAz7b4nV4Z3oRxuJ9m12tmAt1v5/Iz4kS63zhftP
TOo9NGFcXBHj+kERgtyAQWmny0okeMmNUJ5Er71M5BO++KiBZO+aS7TeZju2uz8di38GXyTxZU0n
ayb0eN64rqQdi/454xdZihIbT2qT48uIr279uGf5WG0yEqi7Nj+U9Mzt4f1qCEbNme+EiAzHYeDR
XpOy2/xzNPekl+DF5EODKZ9TXsjehIsR15Q5TzwdDJLDUxseA5aCcFm/O3qFwk/ICdnlJBOR82lm
Dlcm1dj4g9tF3fw+z+657RMpalVLuZFpZ9+n45quFoMD/4JhNUoAY97k8vgmYJ+6LZ7YtHxrkSNH
OVNmjq7BTvzynKLhFTKK6SfZ18HZN+aiFxAwnaIacHpJcFjrxHfBogHqjh18IvlcnE+0FV20uSQc
qQLpcwuTSgQDRSXP9ZpzVujm6ANi4SH1P9jUfOY7H4qunAtU32voYllXKPpVuvXIXDk3+O0r0Mc7
ct0tIiqjS93YN0C3vhfYwxF2fHO7TnWv6npZmAx4a0/xLK2SBmVkK7l7Fg2sVCDwZaTuBGHvv5IW
q2N8dN5jGh9fMwLX4/7djjyUrF50JI6/4eNZ4u3AMSUv3RdRdETnbH+VKMkP+1muy/g8ikP27jeM
+NIlc+VLSGIRCNpihHvNLlWreu23QmEBii9XGIexd5agqkLvzKkTqX63WZzbEUDjApj1yMpIJ4eZ
SGM6h4LjUWKR0b16xYmJr+adntwTKwHEkusLULuQAYhWlDN9C/AcYzMhWJi25BbXsS+Y7ZpM25rZ
DfbSIdWu08dWciQ/N16d630NFoBK54SHO9eNSK4DkAXf+/ZjaOmVap8kgVvWfJWf2O1DU7H9vXUt
5ELSpR3d3r23CKKvkwD6b5ZdLJXUmArzFg5AATqmjHDs1QGI5htbNESJs15QUxaYEJ429z9S3s1c
HXK0hz8OFk2LG915x98JJ8cfgSQ9lvJdeayj4FkMkmko3r8lHJU8UZ/Gysrfn1a63AxUW/8lVUB4
ao3cea/+fl0qp27fWDNnAUizqP7uatnqnG+YN1agBYPr9YF/K1eBAgMR8MTLW6br7XGEfPNIbw6U
yIVoeGPsNqNrjUYb2d1TfpmS5mmGtnv8dUnGF5t9EW4bNEAncS27e97BLAwjuiUdyh+6V2866MMc
5i3eFDC51GekCtgkr3ArigMNP3K396M0a/QjXP6dJL483cSyezxsD+rX2uecXcvoRmo0D5mJFKl2
FQcD0Pdl6HqzHO2REbsg7ji2cT+QXiDfao6Zw8S6B50Ca4JULb9JUgZvG3UoHkZ3qXRjBWwuGMii
boA7UqUPxJZDmVp7V0TfF/8LK+ORA6Y220r9owlCZvUNLQbfLMbRyts5BS6y6rmntXQS2EfgL0JT
V+XWobr2qKzhogAYyG3fOj/5iqKOE+mfY5xQnxOPY9Sqmzk81LIeEwKCLsV5vAGGT8ilJRTQoYNb
ycVYWp1KdeWOE/jWitbKlRsCNrcWOQoFgrrfM28SAmPbNCb6rF1GhbwLhk5J4O3a0Xwlh29kmsS0
bSyxv76JBTbssG51CyP2kRSFqwxwPaFBbS/eBs4Ex0QdPcRl0/G35zmBpv9ns0Kcf/7qtRvoYhWd
AT/gB0y7wToOoVH9+OAytc4GuVEbzXdQfbYVB958/fGXBM5jmYQRDbMa9g+c7mkS0acTDNL/vXBy
XU6IJyHEVuTlJEDc5MZCOhT4qCfRuK2/aG7BotzxP09swbvHNOgXfgMvpIOSo4AYoRr9sBu4RoOv
whFJUeam7LyQyAmeXml7zgdFEitGtC1Gje4Wl+DeeSnQq3Cv8HgoUsaZbLjhV92rP60ejQK6ZECz
SR6rnlcl2o7RyvGbhLXkPjKq8nb8Bl3lbM27vgmnKV/NqSHf1PlooHqZn+CIuI6ZiZEsgQ6qucG2
Yfw53emPC/Wh8l1Z8FagDadNDgWaMYngRacps+fCtGIpP7v8faejaY4ZyFlgS//dn9wGNq4m1Zza
Vg5ZdOnxSJ1zfGRvpMqmP5d2CHvsgwr0pCXiZ2AO1v90n7kN9KMb+juCX8nSvwg5/DY82eHkID/q
elad5thvelHtG8NpyjaC0FU/QFxpOpu3AqXQAqfMvph8nRxzhAhWqYOqnCv9znchhIBUUwwfXBEE
jXhbSus0NeM/OETVu0/aK9vBjG/JDC7jGPYOvAHkb6A/Z9Hubill+cSGwVh8P0TsBYxd+VETa8UW
eYOjYNMzx0tpKIZgwqSMaFWFR5dcYhyCYEAywH4gkNSlzv9IrLtRLFY+IYInYt1vlUAGFYyd+MMn
rMwp2xsy184NfxL2MGUiU+PYb4kOm8fBWz+i92PKlWsrQ7xuMTHV5XwZNgHyskhPLBHlnsuKuug4
ZUhKj/wqPYXw9MErck5EaxRQxXVqCdeaFSCjEftRjyvjNOFeKqLl317JaO93S/B84L/uLanajwkR
KriShxx5F/Q4j2MAC3Xi9EH/+//JnCq8HpHr8kHXfMHruqAitHdxvyjO2rRAEozWdB+qx+HyPj2s
GlidJnfCIR5tMR9JmaEIGDqVUowje0zZ5SOc2sD49AwCDBEOAYYV5NMR5RAAKHefUOSlNzJLlK3i
xg9rCVSmUXzjsWiD8TweAt620HpzZYffseoEuhTSKWJHJYHf5Dm0F8mEF+D+3TxNujS6P4H5txQr
OD9zig/MW0OjvSElzzMM05qkrZBB48j2+xRURqA/XXuW3rOuFBi99afNso/aS5zQK5tQj2PQD5kE
/tkFSjWJX4sbVdm4KekBVWdGxNGuPXF9M+algtuXTbyOBVFpkNJ3o/HJD3s1HsTlXVR1jMOQiwfU
/ZjsX5OXdsGpG2DtOH+al0xl+X5CetkKsxpd2S6ad171chAPyqTBMrb4FgHY6LUCvzwX9Jmr/cMB
WtJXL65Bp57XdWaaRf/VelMMg06SZ+tw56hSD+SYtFvWT4RANp/ufexzJxD+HKCvSHaiyRy9MZuH
4zpibJkKgKhoOdH5Ucau0QRszzSt2/VsqCWpVGGCBK3V0bN84Zb98FOWog2BC8PUYlbqoruFC/fz
AhNWqxwe/yEQKLfOzufEDdMvqdsEiYuPGzDXAB9Ggz4siJhpH1lxIVqNIRR7TwSCI76roMiLZrTg
uzXQYPA1ZRgvw0oudoydkTCagcUzns+rOAlfWqmFAgbgVXmwKs6Dbb3TvyUhGDr+nivL9zpDWMrT
yrHmhn1kDKrBiq/M2XjRZHGUytk/H/KW8SjO7gzp5/39gT3I/JebweuX+AFXsVOu2XuGY2S7mw1N
N4ha1sTKis7bEjeGgJ64R8/chy8ZDaYx/W9ZlGZSBRA0EmwhR+LKyf0ylUcmh9WSceIU04DBeD/D
AQNXA2nOqDI2uZqJlUDrRho4ylUCCS+8sGqSKIWYJJSiy8Ut6KrBJblVuBog/0GzX/nv60zSuwwo
/Z2uiFVjl/LWTfpICR03Jgzj3CNWZd4TP5h3a/MXfFwiZcTHv3owv2tJ1POgq0FeOlT8xDqUTXc0
6e5pwdcOsN9GlOedJiSvka7uBT8lUJ0JuwfPSF61JNSYm5PXsSrBA3mhWzAMMefWZPNlGW9ogHeP
kqr5cNI4WIV9J0mPnD34z70NGcWZbqNOUjzICXjuLcEiGYr4r8gyd9MI799cGQqcOrtkfH2gjjhx
Vhi7ELsuJ/bQ2gESITXNojTl/iNU7/W6oXv8wM+2/Uy6SIBU307Vmbl9Z149Z4Plmq+00+tj10aj
giyy895+JR0u+5W/FN9Bn5xzqczgUUIOo3sngB24nIVPR8ZiAZHKdLb8wRHytE1MnmFGMNDl5P+C
ADyyRbHWgVeCKwc/fyYgoyDU5k7cVi22qAHn0tBT/XlNxdeLyI2nsy5LyZNMUjZM5KNy6ks+G52O
ESmZDpZ8MJ5F9y3Ptr6ufydna3SGeUJjIeyvOicJB2rYykU6xtfX2hE9GNYNj2dlHA+sVZl3Bx+H
K+1AS+jgxPxb89d63RRiZOo+8it90mS6fdtTxxZhedf8xdAjvI0W36g3fwI272OKSwUd/Qd62ev0
zRZfCxlXwtmsVz9UIiiKiYw6G0n1vSkqPu4QmwUPoAvYhT1my1Iqf9PHWY5vxIRNZRL79c1WMjgl
5GdZoQE0R+XllV4LCMe6UVdylv8JDk0mswiEkU31WmV1HO2L5GZj90nqa5AV+mJCceV8tWRe3iKA
mTbXIaCEh/XxjCPG66IQM+cl/SWnoNAXHtChXPQmsVYK14HiHJ+0ebDDEAEgwmKv7czfUQpC5ZGe
9phG2LIc3h06WRcEQW5w7yAYBH95rTmH6haossrHIAlnx2EVJHCS6edPBmiX970j/MTa2ZJdV3jy
r4U1Rw1q9Z4nSpAIol0x5Je5D75I/rPBqcKLlmX1bQsM79ue+q3LC9L/Z7+1StcR0q8VENWOCN7j
W9s0ovjsu5SWELmBQ/f5RH+HmofA3cY/MUyGdHqNCOvFtaDKRNp9jmzIpmmGxHzHd4vPo85OtYUt
qMWTLrcL7ulIPfD7V0uxlzbWTgmLsKSMXTk0VeOdMh5+mhPzRXvNt2gtL7xSRuZQM4V/HwKjQmLc
snu/Xc/sJ6nR12TsXlK1GfJ6zGkVYFwbKjdUptomwlHM1KA8VPX9A20xK7LiA5L6E+vr4dFH0pwj
m4BO+jWoV0yQC14ZfgIjmY5JDuYGeJAu4gjOVVRK1PJiZyoErax9otLa/f+hEJrgxQ7wKdqqxMlC
uxnK2hxc9fm0DosZrhUQsT9J76bLwDNapecyOtTQQockWWPo+WW1Azrb1nRI2CpH//KqZcxa80U9
xBpfDloNuPRO3n3W+vgNLYa+0OzIFJS99gMXf6vII/pE3e6uqEwVMNths0Fx5RZnhhP79atKrlfP
DXvXtv6mp6lWu8Nk8IJM/odJKCBMDpYGN6xLTa7don1OZKsP+nNxljPzWehHDwYikaOIvKRT1CZT
SZe/7kfl+OBX4EQuPcQxp3k4FgnI8yRmgXuS4bND47MQ1+FlBnUNPHt6+ImCjsIyBoXyR5TFkxSx
Dg1WcwCSf1zjGLQXXqtxi8QdHXcGX0N4LZmrW+wcSdZXDBL8kg1W+rs6WmmFWZR+XgCfxRqeqAwq
4HCjuMH5HOgcctu9M31kG/9Benum1DSriNapWKxnu9TD7+pyLNqgpn2tQPGpWy12GFQfKtLW6hPQ
LMUsy6PnrKJle+t9I38R0uPXVyxXwxOI/RIKS78sPByPVBFqmYoMXRyAgO/Ufiy68Tv7fENSYA08
roRpX2uR8KOj/hiWt5d9iErsxzYuJxJii1zFfTiRZQxKxGqfGfwfTXiepHp4Ke6qxMVpb4N9W5l5
vUNQMrNxXllus4hF33iqGHpzcsHEFGsnNwMxf3XtQT55il1tojcgKrOgU+0mLyJIJUSAoAMOOi54
0Tpspea5grKSy+sZ7a8Ni9Nx+E8927AEz9qarzTw5BeoxmUw7xE2fiNY90e33wjvz/idg0P4ZoUj
s40DZN3kq9BSS46TCeDfAutjY01LKy1pttEJhSR5uLRRs2mgnolNI6Vw4P7KiaA0SkUKTE4iQlG2
JabNXqUF5GweRq0N2R/mXjp3G6crc3vOJek2P/+sFr+0dE7zAxat6BIBipMTlYgyODux2oYtt/wm
VoCgiNOquLu+8Vx2WFC/1eTsRaHEHSkTQLY2VUCEImDst2ql5kfxNVS7XJ2PtR+t/H0Pkpjz/q0i
LDIZy0UL9UR0kNnkNmO/XQqZtzK9nmU57qEssQvou+kGMlWtKLjv1hTTimSlz+gDVgwN63hHtLLE
O5KyQFC5m9rdT/16K+rac4wsUCv2oRnXZo1wa9uJBeLe516XckELUh4Iy8Bvlj3Gr4YZDznqJ/au
jdVDlpJGq0YQs//dLN/1fZuROF5mhYqXwRTbf8Yd2cdBpFETpo5dNEGFVtQwbWCLnZ3kb4hRWeAO
hQ/Smp/3sTfb8+KWWNyyTw0u2gdCpsxcNNFOp4JPmkxypXYLc+kDrxtLJ0wnfLfIYtFuswp7jR4c
1yratKasOYflRLS/QY4J1bh9JYnArSxXL5/xE0mTByZFqg/wZMhntM4flC2EM6W2OoMNisIg772h
0zFvg0t93b+v39Gyefc9iId5JOFZzenYKrDWZTuwqqWYRlQABj8awbH9Ro9A+zxQIoCeJO1Fx/xA
8DTXG+whcqxeAjUVkG2Va5Vh0JXyNlzz5djo0MYrBDz5CaiSFGRFcfEttLS+AYX3+F9uhpDpzCdV
/kHDmDYAD71Gg9quBlxyTZ4exalHnPC5cl+WmYRVBTcYgmlLItvaIaZVf+3Hq3fnxVh/s3fgC1mC
i3Is9LPkvyeV0+SLTTe/gnSQqm/ZScLsva5JLEW3cpCM8+yMRZnHzkSyWUzsh84C3BzKgNC5nX1i
jmJX9+/oPcNiua9t/ufxJYBSiZ/LtXRa3pI6e0y5AkwOav81Ie/JHOQz3ST/xRCXfoWPdc+5G/9i
EvNDSVLMPRXytHEaOTRcAbNfFnmOPSAHAk4vZ2R/hqB/jJn2/qu216XK8GAXF85TQT8oUwT1a8k+
CruHFtc08tyvvAubR7ptN77+3dBDdz2gplScOKOl9tcwK/00K79cvFPv3ptObsZ07fTAWOrvTCA5
tp0Yyqj4HP+rG0SNgsK6SMwS6POz0XPCafVPBc9OUwycNuPHeY60GUrnYKFh7kGEvD6AMJxwKKOB
iSHw2kaUssE9l9u1m9lgKzYlhNtUsMwQ6zN0XfugXjHFMyK62R7JuhsaRKOJ5am+Y5PTI3DwvOQV
d9/O1+XEVNNruV8oo5NzCXOiekTH7QN1aJrcg4vIakYWtbhJK3eS7enLTQm3Y43ogP2kGnFgRCa+
eJfT/u/cD6uCN0mjwrl7VJbd3zrY3DUNAqTRUghkCu3uielBqqA5I883I0TJC3XY37rvMcfTGQ6J
1PFiCNuJElQXELTm2xongD+JUYbaoBoxHOM9/0W/bB/mfzOHzd3eZk/vCxy3Gzxndh4tQOR/1Bsa
1gB/YgaJNeVtU3cq2L9fKeRnnYtHZrJFGcGDMOKD7KXebfTmb6lv3Ri7yrJh/mUxGpKWXZdM78Lb
jj3dxsafTWXxWGiDMZGnokyns1Ukv1oV800YN0DIfWPSwxNcmnNytxjZqfxQz4iAFg3SpaS/cTuj
te4mvPsfNV4dgZ/GjlCim4tcYpfNBaN3LoB+Ue3VExaZeI4AxDkKnlyk3YWxPJQlWQJX5oBmjVzH
zKqj/SIVRKgAfxaJbwTVGsMoM62aRqzEpGt1RoyxSE7KsB/5fP8gaxvCJXZsLxFGUAxz1O5+lmm1
I7VunQc17UUJC7at1ZBcCJsNoMmbbP7bxgauKJNg8OTYbwOY6QFiBQYCPSNVpYRMkSMP+r4R8gIU
/HA/wTbu1Z5zW2yomEsqCBSFuENZu5Q8A1R2KW1MTV4v/jtKmfKurU2g8V8kiO79dIWGFpa56Rpp
7XeIgZnS/kLzMN9gQPIR7lfuh9f+irTIywJE5/iMMFWuOkF7ShmLqH69HwdKcRU9N1sROjKnbzRo
lDBkhYUtZ5ywhnbGmFWR6KLwh+RWUjWZX2Pjev6AsKJ+ydVWEz0WM57GET2S9Jv2xR5ohW+zkxFn
wH0Cj/GfgXQyyjfIkoo2tp0+Nah0+heB/4tW4N4T7fjf3cM4Z4ACChKTagnAIsZs4wC0lR9lS15w
XJHNttGvtQBLYRkLBcpGVKKYrgt8o2fMDWVl7L/9ekcs06bPDHfPenTVDovYEyPwS1WdRt6fTMuL
LEzyMdXHi27SnZ2QA2iAg2bN2X3loggFCZIJnM+zK5xJDyiFrWhVFuJxzM1bcy6maUNkdvkdomSo
WogKQkk8SZpiA1eXeCIAvUHlMGrCfILmoDT4ULvagAFD9M3xUnws//1gNoBmT9rVj2yQF3VNk1Nc
0x7d0ifo6NZPVFDI+vJttYWbkvR5wkupL5dKthHJnhK/sQ4LkyI9P0aNL3/j16SJvOyioK6caAPr
rj8WF4TquXiEaBnQTjAodTzQ6rx1JXmQjFB85FdLgrJDZI9eVUzgZXnFeavsOIvpz21dRvHhQCaI
mJ2zITNYRYcHiC0B451pDQic2kMJgPuJsfKNUc0w1jXs9bgQRjNIRAdokr5cfejthlb4YhhY2kdS
9ilUAXWDzSJapd3E6XF55/gEbxQCYfBapbSVWB6+7ZRC2BFnV8wlk7QGmNKLYIb43+tVMmZCWcN0
rd34SQUurv2oVJltw75tbusxhLLF+hoF+Pa0yjWyo13JDy1UkYd5QFm/Hl7pcsjdsgatc6PiBJZh
PgJyhaI5LuRmbz4DZUtW1nj8cbGem9vPyXgN1qlX4vCuwOL9QydYPb8zSPgrt3NRreL7q4h/RAcd
icdaX8uZMpI+vV51hpAdTScqI58B0OZ/YhsYKOKXZ6jKSV80ctyZUbjGC5SE7j6U2UPOnRo41K7+
tn5SvzLYTTY/dgXPgmmQ+Emc2DJIV33oo4VfC4wDWgOYRFOwpHaToiehw7G6i5mTO0awD8mYZhsS
NJGSrlLHOxfkCAva2hGuciqBzE3/GzFmZV9ollxHFTM0doHnx5dHt0Eedac4Ccb5IcAe9diqgiEz
rUJLsQaae24Wu3a2Oj4p3DfpKIpTqzk96wTD4J/spQ4tuMfnmb/2DdETb0adpK8UsozZv3zRNG9s
qPYGL/+blP+B7xY0VWTODgoB7ceJZ9+pj82neOiarn4YQOMXydWeaIWd9nWz+Tyt5JLXV1ErrenV
J+wJzpfRZ1ZvVgceSoxttwhY4cUH+exgDNqDdfQFqjnNSJ7BjXHqH8lVO/patdzclVhZuSB8Ukra
/RW0FxF2zak5Lm/oMNTrab0QaQN9IMreDiV7ngS7QhtzufcLpfKrvfswYfyclhGRuIdqdqf6wTsa
pUThnulFwqBwdHbZ7GXs8HhPYznmdBNxkUXXiLkC+w2Cf+K6Vb1nCcXKPtlLvC5buBReawOpN7C3
BsOadaAmJPkw6jzHThYnvdY66/mAHamZhdkx8RBGbdIwGdUsEoXPzKdfV4VSGKSEdnc1Sa0F1DfO
991cvpM6bpoKnaPwu9HB+8g9tGMkCNzeVoxIUdjP0SPWdAxn/Zc+h29nG2QUp14EOXXbPlVOp3J7
I0fslpZoh21nWuIdJcX+jnU4L4pnWj2JRLJVN5+xTMPGEIPS+K76cUnmfaLt2YwNu7Ys26JRdd14
TOv0Mqm47Co80pBjX1qglroVzOf41Gs1aEHQ+fNPvjYnSFpAL9HerEAqr8rFLk3PiE47NYi18ZDS
YgB5EX7g+FrvVPODfBHIQZmrtNec4Jt0AwQBo38nWI1M/iVNfl3onrueTyaasN/1BTcvpknqsuyV
t0C+vxI6MfBh6BA44kqBK/1h1RiiQOtmA9VNgboCJ5wxPDrrIzt3rWhbqAaFWXwfvr1H9cGea3eh
3+hc1kJKTaVOkX8MILH4uNSEy0ACOBC0H/DtL8NwbmacxWV4zc1T6YU8g9FfExD+CKB3lAdB/Ese
SVrAp/79qLqG2EAc+N5I19vyryRkxkVPhZCmpB1vylB79G6h3ZBRkkE8ly+65zBfFYK5mhJrCf/I
atVYQNd9rBbTCKTrBUdCsejwF6zJuZ9fopEId6bC3Y3xhovO5cJIrE62N3viBg3fDYuIWRSNj389
0mp0KiY0W8tvyL1+Zf8Q9aFQIIgwpsLw4gVBMoAmSY+Q60MZvY9r+SqQ0ew/sGQYKrCLrJLved3V
M+j1hqo7vYvg4bRXnmQbyXB2+qHY/PdibtFFkrEJLUYP9BF4lQ6aXfoFX3eznquPBTC5exHYHAIo
5HY8H7TQ0xF+anLLuow+9bjK42XFsXjJMiMJYAXpwEaN4jsaqp11ipyHsSy3ZR6NXX2cMaaLX1Mt
tgZGMu2qn0GkF5MNwHZpZ84FZhm9kKkiFMyjfmeLsj6EvvjaIcVP8ObFy1pl9rVd+Xq8FOvavlNZ
e4zM1hFpg7PhSCKF2FP9rTf/3rbtDAyiQri4N9GLtkDWEGlxG8D1YI3b0hLtmHKMDX1KbI250RZB
lLQjVNBNyzkEA5XklGClflfosMifNnuM/6J34U5WPKsuUa2lr3rQti+blDVKGQHTmk0vRt3gXWRX
hcS920CvLO2BXMz9quR2yS1CvunZZRIYd5NwX0pwIsAOKNd5O1rBB5UwTjAtxcPb8OGTDFYk65wo
NZyY8gXtv2jWn7hrAicyjAU9ACGswX1Odx868Ru+rgXS2mZifxMswtFX9zmXOl91UTbK9mPmjTnV
3mtkh+w4oLcw8JwIEchPJR0kG584MlaSOwz/SpB1azhF/hsXG1+i6pXeX0Q9x3inDz/kPeQ+s64R
+pWMfFHu8Oeow4vx9BXS6U/ysteNbpfJBC8oTnYCIWkHGLEPH33I95OUzCfAC9BImokCMEVUV6CE
79lTTvFO+90hSLBqYA7lY5hpE2o0ZZ/e+rkWq+sYY9Z+VRwYUsqSyd5F2fxkiX2PjUKOMYs2nN2L
9wws8y53BSNS2KB+FE5XgxxB8wUQkdozmLsgNuXiGJSyxCmuAaIu9OhfWCLRTQoSGiBIkU/QTjjP
afi1CCCUpypTsCjfXz2iycRpSnpFnUsrQCdi4rztaPszYOVEWoneupUOX6K35Zjva2e8AmoIimij
wyLvdk07QPIc2hsNcLBLOVdw+rTTYnUzvsKpml/KgEfSy7dABTHnVDXqE22BDhpScsmGIPTsl0DK
h4a/3NTm6GcdrOoDAIvnEscfhRZOotnpYWGzRkKs5Ge+qLxPBnZ/mBKfi+upx/JrkR8QCIdNA93M
K37z5Xsm7n5NyQQNQq0diaZrUZH2sAMnMW8SLs8O246ingmtAgUFBpVH0aNm5FoKOLmBvGKAZBGT
hsyobv550bFkPPgKPRduK5irxGCsG3P+iClabALAawYL4/jEVau6XVMpjgka5fcPaHViD0gOa6S/
YANcPtpslj55fPbI6tzPuYq3IP5ViL6sopoTzb60PMCSAOcP/lFvuqc+2dqQCfdWBLQrb4TjXIgf
ENPZwnETbpqAog2tiHxImgBHHCZDLobvWf6HmNgSz+f9RE1gn9Q9lCEPnqQG1Wadrd00RYzZUwA9
1AQGWE4CcMgHTLM71WfUaZsibExZ6swe79/Htf7F+5+0XhR3FOdKMKuoSEIXbPfbpggBZKMF4SRF
RaPDgsgzSiUGNLpmj4fx9qLanVMT9pOrE7ZdXGgA1tbBQWNrMrgZZflpO8orzdinLGJ47NuB6cIi
PrC3pXfuN7myBoaZXDZPPJLGGTM2ZWu7zG205JdlRn2l2b2jNUwuOxLPFbHOmdhMfhs57w1fCrZ7
pfIqzkw8+OrjSqkHGkYI4211t66e3vcRkBrPxEdy9cXyIWEJnRjyRifbLpBY83LxCuKTsJxPeO9J
+I4Tsgjb1vl3BzKLCUPU4snRKr9pt2083aCddcowvz4v+jcRwIa7PMUfZb9htiqWN2KFs+NVYeGS
XYEzm0NYsIg/IrdnKTdu99bO48zfSQb71sWRZ4rROwD4fzJx82MuMWRE5g8aW8V9a0nty4KcXNp0
7rntKbeO3l9z4TYzxJJpHLDCA9TGBThkCQp537LTmj/QQkyTWn4P4ctP62+yGH+ggCr2Cf2NAgiB
v8fO5ALwj46rCKDjMpGs5+kK/WVAY5ZZdHDrJd5fNOJLMeLERiD8SN+eh3BqZgPo/ogd+csyT4XD
Je7N9+fwfAckUllrQWwxcmf75V5rZVGvA7rLbh4nutigLJAC0v+VJDye5q+nXQ98Nct37JyffntB
Ik2rv911+sp/47aB5+AU5+4D7Rvw9zdjWOd7DVdrvQ36iqxfSJshruCxzo43spNwZ0Bgbu1VWk4C
PRQVI1szfAm9xOWeLeKb34tDAZSbuzri5PB5I9awH36EjaYPXgt9xYtzDg/fFL6usbx3+EsYaUjA
qOFwsBzVDvpYzNXBK6heRGxmBSO5n8w9zrBiSWzU3ttKtNnpI0Ho0+nUkYEmzoD+6rs33IQj9htI
+jzirB7FIBWs+dQTPjq59gpUxhVvTBpHMjqfYEeRPVNcLQ2BQWkwwvA9w4vWZvI1FJnp3jX3NEmG
5KlInD54yUq1ufLMl0Z8otf/AXaqBy6LWXIDjeyA0Kaz4F8m/qv+6RqnB0IT+vLK92sv5TBQjp0+
/hAh/eID1BYLgxCNPkMoipVXqDIWVu/XHKe+RKi4gkjMEacCWa3eRgOirNdiwNxGTLlSDCICU6cg
aaadVIG6xCdmT4nHD7UIgz8lfkKV/LbVRkwpj9sn3xWY2bE3UYUFoG0ZroGte+q59bDCv6wn6zOu
kBfA0ygvv2n9FUr3T0/Fz+SXO5JEsFvq2KsZ5j/WWnithoe30wlfoQ7wnrRIiPfAJgNEXviC00kI
bzh3h7n0vdCfyMQ1baXL+upk0ZVlv4GBy3zEmCkps79rLtu8k7Je/hMagnjvHLHWgf9uNocb+TQ8
m1ozgZSAqYqWF4VrztT+p6BKXUbIJJMQcPfumaRQFDNPQd5+ycxfiyKQ9DZe998WHqyOvtf/mWsa
qI6KBz7OjIXKrsQFPPUXBTXfcrOSXuUoLF5UUT3alVCPy7OLK7nFVHPWO5XImIIWWJQcKyy2/kHs
2KOQo2zhcSxNSDaU4+m6J9OiYb5IWAdJ5iHsQCOCwv0/YGRf0ZHt78w0jVC/bqg2gDv6LkpASeo9
7kfdaGsZAZ9GjsFCMspoF3prpV7mMe3+MavJ9Rphgll4YelcuWwcPNQzyjQsVXugsIw7nhR1Dtk9
B+NFfrPCAbPCH1SQc/HV0cuTlNQgiFc1G+DK3ANIKlWZTqg4Zjh7hKtQqEeROMtnEJu1y2KinNOJ
gm2rm9j5LHMUChldC+csF7ZpHKbQfK1dCkNTjDSdWrdZ4/1duyk8CUuQwBZ5SHF8+Y46jZvk7dDJ
kf5UroTEXfY+cST5QMJ0m+9u2qk1J57JVGuJUo3Fd4cOVjdESB70TX+c/Qcdzr83W3xRmFELQTbq
rfW5rU9bjoY9AZIQyva90bPzBXMkODdhpYcWiNahla5wBn5LPGGlBHk8ahR47TLCK/U7jdQ7qnde
RYdBDrHe0+FL8cNs6B2JiJRyqLhrUTrUIY2sYJlW++e91qA888T2ZUOGTUh6kf9gYG/TpAG/JUPk
WRogjqBDdzA4C/nC2jiqNrZ/wf9SlLOKKHZH7Eg+l8XyPC1eRMEwxkT9StbZkH4uGJI5mYFux2/I
xZrYDR7bqvt231/gT+ZL1+KifMUbROC55sIh9oBhv07Cz2wWCuPmp/fxuVvmvz3Dy6xOVvffOeF6
ItRdI3GPa887cuyYqM0MeiVJB6TcElYiwCuErGYzI7vjgLycfqXpn+gQhOU9+6zSszIYD7Lc65qh
+y0JEY7p359yipzSCghra0mm93bVqNcR+eH65p8FdHEX1aX5F5H08D/W1yor47x0baTbLwox94Dn
MR3HQnpL/PRREgdS6rbOiG3xro0LDRLkekKXowgA7k7Rt4XzIBwz0F7pi/vQiViBWMPsrsBkBFG2
EDvnetSMUCIJIeht7772V//btw1AgFDkyt1sy4CqvAF5gGhOYpLcrGY2mBoP5njo46QEZxsAYwBt
ry8lfCWFTtQKnhQMIoC2gnrI00XZXSVsjAsH9/DU/SOcTtcu/gD/KCBqd+TGnVzo4TFNtDYH9uRq
PK21Ad6ygF2WFSxWW8ukb8kvKrDkt2F1g13FSmfk3mKm80A45ajvEoNEVPIWSgwwip54qWXmNlRC
fns+mpCaGFs39pvI453JK/cU7ebBJgfg4ycGKR1xCharKsF9cZFGArCoK+FgKrdE7ZlfH8AoqnWx
y3P8uK1k1+EMha2mBxAlQj2kv2PF2NE0oFTAmdRntirtOtt+O/P0XIyySpKMR8BSLBN6pIi7Gcdf
WPmgzuQiyp0/IR/0P09lSBZHV10AUJ5vcmJfqyV/5y/mpeAD420wmMhNJ+8adgnGXcLV5k8XZEhy
hJOFaaAGzrVaN+jfvCNyNS4AL7RTnGb0cadbTz0J/3Fr4FM1k6qHP42A5lEKOr7ehObvck+LWNu9
77qBBA96B1GaUY/H3rWFFD07A1iHD9WtdvdvaIe8jRDzm92euu0si7Czp7wo3+07+HT4aRzBV/bn
zs6Oq1T7HvR3cPA0wccTJaQQJpbFytgWva53TCmSUh5uSEeWi7Nto62pKGx0XOXLEluMMIK30s0U
2joK1Y+8j5zo2Cwqme0hZT3VzT9IxARhBFdiTR05S4IfliFnN6kyay4g7+xSDzCXqLYR1ULv/mRO
06M4uXLijSbFwwGFNhQkDlm7Gs6Q86MuYGD2v2ECbZxaaq++JIxqTdh3HIzVhqQNkiTahHppfwzG
dMU/0AAfC3OJiA5DRsarLs9O+/7gHQ2Jp5Fes4bxfIqUu1r9+2Cj+4G0eaewPBQkn6XVhTS6DaXE
BUY4w9QyGxD88XclqFUqbvyT8EwaxPFhQ1jy1aALghGeHcjd3xPRleMjDQoVhW1T0nvwqA+E2m2I
EC1f7hmpK29YgWN3YE1rdAI+svZ+b+6y0JmU2tyVpwhHMF9dpNn/HLn7vZ+Tefl9C2n5MpiAMFET
gxj49arZOB/3VmFFyFYs0G+D+UOK1k9V5qGLA51hZ7Pr7YqJfIDfjIkI+JF0xrwWRBhiF61H/KKo
NJ77LPR8pedsiyQsNuGpeTI7loLMPutPiWyrCFJ2Q0Tg6AoFx+kmrbN+jUaqOgS+S4HFcDGgV+uD
sI7fvaM6tTeQZFPdlyLX8V1/sy5V3FutWnFGjDL6ISB9s1woXZ8ofB4SHzPhQz1xosGJg2oNxwQa
F2hAvIQakzD9bXOvbmiXV5Ab5rzUviiui5PYo5SrjATInBBVh/J/z0CR8DU3RnnVv/XUceX8739S
IPsnHDVHi5VXE8zmxhGoYZwi3vM0VOx+aceCTrSmJ12gbKyxg6z08GMAIEnwhWCQhrT5XW4Gcrq0
hyRPDjgpa+NCbpbv05j5Itt2erx7ZKwRRa3lRZs8IeoxoaSIaVWCrOzE1CWuXWTezW8D+J5Y4W/a
2ITHl6/0nA7og5FZsoD6gmspZOhiY/B4mVvdCpq1ww7WKHmRNwDEYO6qKmocMhBjAmDdK6CaOM+p
dWJJuwDJaQL0mYI1pwgKXaJTU+BJptaHETrjQHwVr17oiue01iC1ubIWedtzyNlNddI+R+h1Z9oA
6NhiIyHPtLaCwKtOzFKofG/GK6gLIctprlpl+/ZXgq7EGeVL4ABvZ0EFgzNINivDMmV2iYdid4jt
5+fvHDQTiGlfGsG9R2R9YL/kZEykUKY4gJhD2ilTGRts5rhOICD+sJS1cG5zG47/fxdbrQSw2XOP
Oj7vVoPdztDZROCk98a7Wc2I79Hq1GFPf3A/q1jtZ1hqzxkIMKY4x2E4CcXQ1D4u/I+CuHB0W0EN
zLBXG43HqwirRmE7Oer/UvZc0A/4+3to52i6DIb0Z9zcsqsN2O6hV1FlNwUj9wKLpnWSi1hriPEs
bPHISvDbDBfeSpsaSvor17d3J6oK8GM2lsG1p0iFv4oIUkzFRGAtnNZNX8kX44s8tgpuvZ6M916u
RKIih37VrJrjsdA8cFYGX+iYzf4cjcXJ9yfWwxs+pE1FzoghHR8k8i7l2vSvoyCpWknRPqvjK+kM
E0pS2zCHY6EbIL+gd9Yi+xuzxXMUyzColcSlDJj3CfrmSiKqsAxcmJiTO/SEbI+EyIfaTlh116gx
R5z4bBSOz/cpPfGsnaf6lrm8gqq62Gdvs9OPtwSUAIR2F0Pmq5xt9Nceo03bNOHjiG6I10XCyS2z
MBZbR22SzCHR6owqKzdRxVHQcG4ghvMoCUIV1hXyBahyAE9gZb1uq5JlnojnatV03xonSIMl8EW+
GEYQUGCV4Mwy0Jxmd3evIQlBXcUXVwybbixh+T5dM7QXMeGQe9ynb2b+DK4oiiqwS4EQUsULMFp5
sWpMppYLmcDYpEHK0AzUwQPZA0jhFZla+1AiiKcHPQv1uNWS4/zB5HqFIkzGpUdo9wgmP32PTCdl
R38YEbkOmEbAeEtjQ8k2M0rX9ZonrtLpa9rU4xfAExRkQGMDzbc2XxaxE6upqM6LeHgN1azw2fIm
wiqc52Nb+SfDq0xGK0H+BwD2KN7wr4N74VCqBjk1UkX+GHqFT3pXo/C5UFOp8zcVCRINgXhIqMav
38+2CiFqb1DjRbnmAgsT82y22lh5mZ6QwsVUWzV6nCkkYC81V31ROpCVs0tR5teyUSM04jTzrZWX
L2LQM64Q/rE/6o2Cd9afYUUItZlF1Gg36mPkA79sMS4tz91ttNfHxyOIhyuIzFKZ3Z9yHMXk9HN7
uJCWe99oVUGT6Sp0Car/Ac62mG4ifLDubBcf+tK/PhJ9DcJeBkoXZZLvf8HtTTT1gcOmhqOdJW+8
nYBHAdAAjgTrH7Ocp2Ln5IWoZx3M0TzBrUyMw5g3+DT9HH1CxlMO7Bu/+9jIJxb3Dq/LwOXvvpEd
RZbx6qw0EcmFul36EkM3yY/WYnBa8/sy3e75tFlcptErYf20/VZMSMFmhFEehX4tT+I+wkCdpo6T
xp1U2gNaJHqrCQfAx7R0F6oP6xJMVZfnSnWjkc+ed39312FZiYsYQtW62JU9d77xc51FTlsW3+cB
Z/qoKPy+zQ+cpfSR1SOEZmMD61Agb0ZC3RwLbVZlIcMPjFalqC6Om2lNZN9P6/ufvipSRG7KstRf
pJjZs+xfyU4QQ7EkhuPqP1rwfG/9M/q6kqNBqAOURyZ5cQpzpGbf7EcipFEMx7wnIgQLmPuRHcif
Hd3zXIB0K+W+moxlsG6iBVkuxVhKpSm1VfdDA/k6ue4D1dtsag9VP13jiXG7t477PmjD+GS6Zs/D
ly9MBnukrjuzP99DpiicIYj9dw3B/VJAdX55qqtEzY5opMfR35+YVmzJfYhtGGFVCTDMKxEpqtuE
nYznB1gxmxryLHcbq9MWpe65VGdSNV0hVznJuV4Za4uM4ScoGJz+ZKCR00qF+8wv5Pw38RCjX14m
zRBusY+90FKaip05F9qun2dsDvGl2e68w6c3fgIzLAY4DuN07Yj6I/tRD8cEhBDzDNF5yFq7Txc6
rzM7WbOqspXcteI73qVgx/E0+SEwq04lJEv9LuSJ/et7SRBwpMW70XSfS2hkhClF5+Izd6PCPKeA
XGy4cfOZlIPV/rm3rIhH3yHSm2RwL4DSZTBNIlWOm1Svo4vqtxxUJg0KEewNWLwUPEekMKCgFxEE
utC81QdYRD+82vp0ZN8kaynkdverGyoXfRLqqCCsrwAkFiZLagVd4XJp6PiMkwmGm0wlzfxu5/V/
raRiHuM5PNnLZXRBwRdVg4Kc7T3ccS218vsiuMyep9JfUFNmTrG8cEDj4uhGSNme9gXnz/qXqiHM
bSTdm0Z1cITIVQgTga+M4n65rPqJaffZGhPHJk3/oKY69I5trPJMsR/3CwjL3DYQyyknUsEVIr8t
875FCojIPdxg+TzWyrX7sgwYekl6jput7AkcybgySA/+rUtyVp31F4mUw443WiNfltfO3fpueBIr
knEtMqvOEG8/OCT8lcKbIyBXiYSCDx8e3shQ1AK8KQ2DdDRH23ro8KmIqyIye5NiCJXf8meMjjB/
h3jeTQ1u2svMG277HuwvA/AdlizE0nmPBkNezi3T8zB+BVXGvH8tljJdE2x4IO2CV00xkkQgwakc
FuksTpCXFwuDKMI+VvPjKN7IG9EJSzrwGl2S8d1UvT+Hrk+A//DkTLmxvMeYwpWIWdVF4149BGnF
8yTcV8m686XFs/HI8BZqqKDzMns3BzyN2q29E6CoV50lbRWpCZUiVA2mOqCRvhsNJ98sqM0ucxY+
81rUynax/LHXm5VLJTVXXIDA9qnZp3UDUVGkUtgLfQ6m1m8RwWWyPRkasaix4h5esa8Bu3lxJotv
8kdNY5VFAdrI22CvroZZ4XinNaZQK/gi0Jjud7sQltJzaucIv2jWt0Ef8PXhHGcODSsduTwP8xX+
ZnOT3qr210B6MwjSaJv62ECWRNRy4ePYnX1Ya7ceCXeMnwtf5C/UgHAwnZ/fCaHS1/Y5Jblb0d6f
CaTQudBqgjLP/nPlmLY+XLcqCbG3YzabGhzLLMd9eEAzizuCOqfttun/2xWRkQXck40CE5AT6ODW
SEiKmbmvl6wx7fzf/1QD4oISJXkl/IzGVRtT9aPX/c0bLH/iYzdm6I1c36VfippK3LcJUfAEMqZF
kNjxQJoMIK3OhwAVkoKO0oEq9I5B9hwuA/Cd/+BMcI8f2J/3PJSDp3YO0iIs646vkk93n3DyE5EZ
MVc0FZZxXvRjfmFwR8r5eKEHS5HXjuxJAVfhp390DlauP5EGbYPsK4D1M4/RMCAzeLGBtQll4xg5
jFbuJ3uIq3yeLKnrPO4r0jwC3ELxL7SxjNYFkbwBgUDtCtVwxHvx1Vjwc9b8iqwSBPuo9nVX2JF8
nVhbMtndqzUIRqqsVJLddt/gxEk8n81M5mdA6KL+0rqVSOkeqX8dpakU9McN7lGwNSMwnrSL+qD6
AemB8a6wr/dnBaK/eMJTrjC58YsKDA5WVIDttS3YLRUe1Q+0IQJyw8q1Bzcoxf2vEDyIbm17rBYT
k2aZ8t5uMoVUKbheHWqLSRbTYoZkdlD1wsFtmlLROK7ebmlk9/S4QW5HNDETMYRMAASKCK3DUUmj
8jcGOpVWU03NGAkfqChfTCWjDEbl+N63cHsofLcDRVOFmlsaVblXed8Fa599jdtYq4GQZV/mv0aL
bhkQtF4Oo5MVjtJ78VXNqtx1m3BT+WNfAvN9OfYCBIKKhqq9N1Q8nsfpQpqpHUlhJDM2g/cX753q
S5L8uWIUgevWPMRuoGUnVMYf1FS6mzHV7VgF6Okjf27/7xRFFS8E/6HRGpXo5WmAumDG9622ZRsM
hskbOLjsIzRk94igTSS+ABKolkghVFagHl2wh4AYgUzsSgxNMajydA48+ONXmH4SJIqHchZda0Ho
qNQlNKBXUFgQL/ju7Ita9R+MSH4nE4eX4dAHWCqV/Qhgb6JzlFhMtu5YFiIymhrVS9ngxow1PEvW
Bs73ExDGmSVtf5bH6JrcEfDBYBowF6G4c+mChvvf9So20nRU9dpeFJbA5AGbndxAVFasjZIqzldh
fFsQKdLcm8jk8dqwp9kZ2JFj8CV2glv74UXkWd2OvLAZX3oD8EF7cPTA0Jl9fVWMfTk9NHvbix23
/bZktsaRZU8IJnUSV62koOd+zXuCaR/p6sYGMKQJw0zoQhIpMY+eKMX9B8FeIxAS3K3KXBJ8HGMm
s40+7NylpX9gCrDqUyx+p9xLLHwkjXE7nY8NAWqW/0lsc/Pli4zF/i3cUzRnnizTm/uwOs7zyGG9
j7ZIEoOQBHl2ekmwOJ2FdlDeytda7wk40sFNc5hql64hDQfNfqD8npD0HasIEMFUax+pEkI/Es0U
711m0v+QQDiU7+0TfZsjgtzsrUGkyDeh40VM4GHOXmHhs6Egk6H6/kD6lhjTd611vZCkkTRTUmSq
AfrFenlEJZcx+Sm1mBAOLJWBIfOixCtoqn+Bzdu80aKP8tAgs9y3qltza58Q7LObRhEvkgbOvn/G
65IXEedet4e01Pv5k54t2yQiltu4s0IWOFpr4NR3qi7NvAwOj81cP3cNJKW4do/xGtE4/qdmUUpf
Ljyv/mAZRB9+JLYTkAoH8sZEgfsBv1F9XUOdJONT5b0wGqDFiwV6ESyG2vTrY3z6YLrm+nEL9a5v
WT3bhCWSsuNUTj1/EJLZGzQqAXgYHtBuI74J4PvibjIArpsxdSIN1cboLus8dLjEiRk0eVMCkWZQ
TolxUx9v37Y1nXfyj/JVI4dwAUiQeUrTT5eXWTOuJb9xU/DY0b2tHr7bwMs6bOzOmAj7SXK7lzJM
HxTKCrIiu5jPEYOhxHR/x98ab720gJ9wQz2v/nV9qOvt7FGBb0vR7RTi4uYG/YO/dM2jEz0xYMzS
N6fRT27sGRR8kDsFJz4IlssckElk+8aCbNBChgSzZM6bzz8JNby1uDM7EFSF8YU1W13q+H+OROqg
IT7YKxU6gb5ogr8xELri38VINbAW+OO0px7+SRIMY2cIjNtEam6hmFSEQl/4nYRu2vcEBoPls/Tl
NYUnezN7PIwWd98O5BOJ8zu3PmxzKs7jExq+EGvXbxMnWaf0BSnu1YTRAvb0iLEUjfOFSnfW4rYG
Z55yEHQXFEk4PJOzh43bJn5MFbKY6KTbwnNTHVQ3je2Z99ZuPeEf0MCatoJSOumiPf9ehEWVai1v
XC5A1foeQgJ4sRTMQslHsyKSL7K+lP9CPAZlYCQD2bVE8rrhnOotj9GxjY8fVewsFccZGFfuiNAO
an53eePNw09uJyI04KUCHqL2X457VSudU0g8IAiXk205jeALOrxeSAPAGoxCRgpnuRhHhMrGJpFm
gFbv1krt+6u0z5FWi2Coa4ruYtxvYOXA8DocI5KEH/nb3mvxywlEacWVEPBa1/x2YE98M94EgrlN
LFNscWDExMbTu7bsnf/A0xQEiy12IFH77wVG2wFE7NPlauQZYVs+MomTGARO2aSZ7WIENsDfrVuf
gjbfPYMz+kxe14SVol4GdwNtNoT6NYs0tFaw9MGJvOmL7ebMDyCkNC6VMmg7bc5RtpUNKrBP+0Wx
FAZqrdmHu8oyNzkf7t3pYUOnmqJK+VdwwCHzUsgsAvKkPWwAG15NG0b+45rmnboOUcfSPxt4YF+A
IESlqocOaHkZxeKkxWGQKFTCMLGhaTXpJcxIVTHQLRafyESh6serrhoqaO1dLi8tK0NvyojtIvno
7C7GZO5mBuV6tiGuC6iLk8La3NPGgvIKKPiWzHMrlfSqIBk9dQiveOvMIY3996GPADTHNe2VlWdH
f7R5NmjcOAyBMERFYTAENBAWZW2k08NOVdl50wwWX6mslAcUCakRhokTU253w9t8lcuJY/Zj64kZ
2FkFPZFCYQL1bEIuQ8jPjmsmmYl02ejoUPz27cAfcxLn7DIM/PSU/2U8UvUQC4E2uBWXH8qV/pig
AHpiSZNm5rmcw605zPxNtD8L8hY+H1qkcLarlJ/vL8whDdPdEmMfn96Gmyj6PmxM7KAqsyH/qsHg
MZEtUn4P+FexrFwDUJIVv4oN3NiWA79GL0PTd5ITWCd9RRsea59AdfEJ/NVl9HrNht8t0kX0DnHE
t/EFv/mUWQO/IaGJxTWiKMH6lvLBTwE4sMbLHg22Sf/bcKmTv3Y1M6aqT1cxZAOPKwlKQjIXNfGn
8o6GSllNAvrEzYYCRaoAVNA6g//1FxJJJOMM2lUZ9icbKljFS+VcGAt5DZTffR/0/OUUwADNhXto
gruSj/GOrZGT3ALsIXR9UzqOpjpRrJyuUPgR9Ik+pTMidN6JZS6k9Y+HlCbmdKeXEjoYygFynVXN
z5JWgmHeFTJJinrIMFci+HWZ8HSL0zZWLksg4OsOzO8BJBqkzHeTo45GZVlE90LpiLUYAiO7qsCb
q0Aengy7GNABRg9GHnVfKqZ+uQUOQRBqUUoor6s6TiQtkTD4upEVGgwLMxBzCfSY52CDxPGsERT2
/ky2t2hyQaAQwJZr09hdXRplqwkc+kAjLpQ7h+Fmyqoz/C1cFxnLwmwX30qYfdDPjZZLsZM7kF5+
rEW959E2fJ9G40jkWgUtYpsv5OUqrB4UbGnECrKbjcrfEIsZfuhiMTtyHj4MxEi2d4juDtBoXxrm
/VRTuQRZ4IrzdyeFu1sKR574dN+y6Ny9MS5fs6tfDWtMEWVrHS5W9aDJrcG72Zm/tTGQ0SATr5Xs
PG4nU5bUndihnxTlDiQmn9A0NP/mvCy0VuzTk5xAKK5PVfZIonr8C2QooylBVzt0oW7t8ftK3RRo
TizXrJlJVw6U/O5z7ZdoSsJeCGPEuaDCo1MKDUjoalc+WXa+Abg9oOqWyIIhV6qdrO/Ae7DLDz6p
SF1re6qpjWmb6VezMqPMsc4Vr+ULeTCAjlVcJeKZY8IzGG9jAa/CHGa/CjtjxIkncamQC3pfEufP
0N8OyWHGMaH/T9XLHHX2rLSC2a1IrbUI8e4FU2BC7LkaWHvoK/3+nW4DXrhBn2R2PSY0RPeEk/jx
TdoMR/vV/OEmSWMzb7Mm9A0SyFE/8veVCj5/9M7hLiUXvVNoYgS0QjsvTym16DGbDsbGi8oDgkO+
7MRLJMagUQQE9S4U+aw/jBguEH/kUEqP4tMF3ocLVOmj512j5o5pktwOOMMjGs7iyWyOQdlMBP3M
1TqenCBduxyDGyc+01IFMJK6PVGQ0vMl510ip/fNvj5mc3ffUD7ZzThC+qmvlFVKNaqfDPQIIRO3
GaG3yR/SwlL58YNgRYhxa0PDZ15biHmyZ3d0uN614NoxdGM/6ST4jqlq7mUQ/4V1XVspIoVdIuVg
0WGHACgkIN5HhzE8uzSVJIyGw6xsY3Kmsfq9bVWzskcPqMfPOak2UiPNEeH3z0/KGXvIsuZxgg4N
3mc5HD4KUUFf5nUvXzTMB1Q77HQcFnf+U4fPd30P8NZStgeiUY30K2th6IDlx38qc8ZzncUiuEwb
SY7mEPfhEdEyDcwOpfekytd0j5ykHVJ5mhIlxZZ8SxSA3aIK8JvqxOHljN27tIapN63JTYkKDyZA
PfOsPeRLblCaROB0pYDWs+/1AwnK4E+jzzmm0C2RAEBpjOpwMUzHeLNNskfTp37BTSIb2jRe2W7s
sJWCf62gI12VZUNogHCPHbcdXEMZXfvShfYgOONFEYTvQGm+gTdNBifS9StvFc5C5rdADt98Al5y
BTb0UVP7o6UpBBRBVlXmVU0t1nbWWN0iya5JOorihh9nrSeJMRMHjpyWkMMpa8zUHInzCai6oNwb
Mw07/n8/dbdEh4UgoY/CqPT9GdVvzEj+vph/8tqNUhTB8WtDgLyKqoLLsDKIUi0Thk9ezhJpssi/
ZuFHQx8g5Unzd0a34gG1qMpmMAPa3WA9Z4sxQnX2fxxlPCaxMzxCqdLiKGj1g5BP+HZZPPMIULMe
etUIb4j0daCF206v9r86jsmjCAoaybU8pFdg5GirItZg6qWMn6NmPHINYBtzUpeJ7Ao3k8B+hhgj
wIsLiqCoQxfQmGa9TGSw/6bVSeijdUrjNIN3UKYcJRwDarOVp9TKb3IN0JYAhoDPhNQ97lILLE9a
t+9ckdAATdUUbj+UNIGRjwOGqbT6BbPaspQdSqXNlK5DR88gWClXjyvy/SEbJ2goK2y0+QMLVhLG
Mk0XsePEKUeAiy+Cv7Fxe3ehW+ekP/yOhBP4U2+E799eLM7zTAJA2QGSOYGwGwey5nZrDMJfjTMU
DAI7Bc6fe+IHlxGR5TYE7DLCu2kcSSREvryKVFRFbrETLjUrocSpJqsFF1B96rnnFe9emzCP7TGt
xt/IvxK63BKxc6BxJaNzC55ohiPJcIJGGWyLzyyaHTXGfc/i+GwP5+Lc7L+qLR20zdhqxrH0eFeA
U/fD/l0olI1V0QIBAY7+29jHRINcxZ8AytjGGYHnTvCj37VQygL0AO81rs1/nhd0ETAjcvdQqOJW
7bcffcYuBeUdAqRo4FX7TFQanMFnlGfBTAufHaQ5PJ7b531cqPmucxnP1+CpMxuS3yUrfXONq5ho
WYpsRTReopw/L4yBNHJ8p9zlPdPdsMMWbGcHP8GO3fix/CXcbWSqwvoZvViOolqAUQtpYuNnBnR2
rsJyFvzBzF8xmiwoNoSSp/NyazZtg8oRHA8kOrLfUaAe4mSqNJHAUNq49Jt9vtNd7iEbnZZhuBo/
edB5q+ZKN+vJ8CVA2BrJKfARihPn410tQlaGDDvqJSrdWkbQK0DWPUlTUItWrpHb6cPkstnIVKih
5k+RVGlxDYaylqV3hqtbgOnaA41Fum7C8g2xEEcsuxKfpempxjXNTfusEVa/tBTCmcmd1CrRgLmn
WnCYRDh1h1XhrM6NcEx+JXiG53b4u/XDxoGpZzNCaeul/0CMdoQ1jbWRznBlvXKBjpSrVoy6N2ov
y2F9RNvD8HEwlpMA/6Phe5Xr8kH3to9I8uz56fMHckjjJCu5faJv/2XBnpvNzN3lggzQiGL9StCs
Icq9bP89r009jvV+/2t4EjElGLI5r2t5XL79irL0ZNuEM4g3/zRVxFpDFYsALQF299HM4e7012Hj
swDT5lfAmSCryqX1GR4AMWmW4a/PWIk5HZyI7tIHfXo/g+cpeWrXxhqLIvuZGxMsDip81u7bps2h
GAXc/ZYqMfD1WHFIPA9Z1kI60jSejoL/Z7PlP+BgZOtedBM/PmnBtkIXg7zplTHFDZTi1DMZp4bH
IfVrg8nyc2ARizmFvpfEI+fI9ntIHMPtdUXWIQiSzZOOam6CrtmBQshNjFa3UrSJNQutuVcWxQ/a
ZwrGYV6gqqWDqxu4U3wDjlSW5f+k43GVgjd496+ABqlLh1E+3tgP6Q5yPwMpFAE0SkshTw2Ne0ve
11w23in8Cjdy3CQfy8hGQHLYzKorywMFNJp33smTSFF10TVJxAVvMdb0CysXNv8sZGe8xl3GCaj3
mybR+LA6CXHKlrQ5aV3bHNlzqv55MvMRQM1dg7C+Akj4ehhoYdWu81GRvnoIIu0fCBB+w+ssW7tM
KsloUa6WvUhF+UZBzRstfUcEFmHPpt9LU+gSY1UuE7Xt4BcjrRLOgoGoQRGmwn24mo9+eWdJNJAd
Q+WSwehJrVG0pjG+YhpLsTzSNCTkl5lykLejW3M7uc+F7XSrAF5aaQJa8U+ojEm/5Sep81b9/Lji
29883R+oUkZBJARU+xyIfkOHx5xCxa0qTMj9qDv/rTRXEhZsOp5kP652pO46IpRcIhoOamdy0mtU
xzlsysax6p/dSzvQt16C3zX/RVBjOuMUdu5obzOuJ0xRe58eCtBMVLZVSubug5y5/Z5+fhot9f3c
iAJb86fpLQMxf96VdqTexz9QpTJ7NRKAvUSCWRBlKTBPqEHL9Dg+Jpk/MoykVHtM1Ki3Wjb1iRo4
Lozx2xN8R3+cN1VxK0lgee4duySk6LXiWwFhOf/FktONFqFRfmVkR0bx5WDPXHG3CtuYDTzpE3gl
u1Y8GSzpKS2IfazhLjGsOGEZYFNGVMKwIPdZovmRVpilA5GublTnW0Ooi/uKegJaigOQn/N4f1Ol
IsEBD8kdPqpqnmXRzxwtgWQ7fu/88wvAuNRvPX+8P2o7dfDlcJKa+aX47HMxGjlYvAV4gx1mUEYd
ZbS5vfAYJNlEJ3KRuQ1dcnspYy6anup4103J71SxH1kLzvqm6VwzzAFHmmAg5TRl15vB3Z6WjfYI
12qopj7DTSBu+RPZONdYB9sm42Sdix7H0tH2l1cB9bTvOrkide3MUDXdkthsy4mzSM731C7cGWVP
D4+g++U7vH2efoamaMJe6GhZzt5IGvzTpu8CmGfG3QUEaYTOq+lF8gzmOuLQrWvLoegUkXTevpGW
+zj8v+M7YS69Dbz2T8G4t197csgZ5vmUZL3qm6zqDnhFNtTIuwCOPYPLbxDwSEX396hJ7BLGOGQS
QBu86/i4oYlsRN4mBmJs/cgztO4izaHmCH0Y48gO9tAnlHRt4IcZa43KwFlZ49LSzKijLhfp8mG2
Cs7z3NPxeZPn0OgL3X3WSqljrXZBxMSzWV7xtCWFMYr1w7+VEO5eN6IaZai+OinIOPpxnJc6Y8LX
bHz03bR742cNLBs9kexKcbu29FrJWXR9OZYelhk1a8ATDhNj0qb7XDH/xmvOh4FzWKYVUX5rXc0h
L6C1XgzmllYnBfGKvMaidgw+0eQZtWdZrl/L/jzkMhCrF5YNwCMIXKB+TKfon+eTCNkULOC9yc2G
hdmnD+a5MzoHYhMu+QdQZeSygU8nPWnpnQqk9AVO7aMw5nmwSb+kwhkNRK8f7X1HJvr81HFtEkxi
6QIHK1u5o+e4st/1yGJMesdpI+1O8yr1lExHe5myxGMA++ajUygp0BrgCgPM8Zp6/fjHi2BUkopm
F2wasU4KfCOVVI4tIc+w+vNMxavD48Y2hUyS9lt1X2BzIvW5vDeQGmKPDGqzz08sDLaP3Kekb9kr
J8u3lE4zImUHRlZXygVkb9DJSzRpz6i7tgPhKWqxWEwJGjJ0sa4B11f5s2o5DyPtCDjubHg8PMK0
ghM92O6mV/LOh8OkobGajTQfg3z5ZbJF/nPHBWvgEiMPEbJXHMxqPMItcuOEeqzmPpP3SwZJOP3M
ZM1BOfjMeYwSKIzUnwTYVW5a5ptPtFL98lT17hhQk8Is/lfw7oKsrvs7chn+1Izyt1/a6wZ28SKj
xCYbwnp+4arORVEIDDlVgJ9LKHvmpUHa5DfMVTIJnMzhT/B9VQgSj2mbEKtxAjxDUpJKLA2EvDBN
3WGOwsZieXdE6BssXB2vtacJm3C4/2kr6xAGOYArxzs5+xkJNi6X3evfw2ZWg4+R09HCo1Q3OMrp
TOA5nSoVUqql46JtA0eKgtG87ZOeSgt3nxfr3WwmEs5v2tOug5zn2DsZvmzIzKKv3dw15b064O95
kOP5DxGLFRanIavnp3UH29O+oKV/+52IkmiXUCA2xVKIHL1B9LdYHxaWEJL8N2CPumt+lLfaW7n8
l+Um3rwx6S7oZqSgTGGl9LoGWqa60lZKyLRwkuUghz5rmKoFgIM3nNeXrLJa1x+LZHsi542oYPJD
NsARQK3FgN6B6pSFrGUkx1HjOCgmp/oVY2WQmxfyG0RWUu+TbDNETOO+cmVoWiRtdZ5OnSEeH1/D
glgeEnuI65Xtx+FnpWHDMNLwt1mqo9psaefX7ki1D4ceyUPzPRFmTRCZvLU3OLMDROMY2iGzAhQm
KrGyC+NZyqUd2Lhp7HxwvXceluH9agKC8Cei46N0EMUyuljwsymvKCw/fsGpT15xrMgTj21EphRU
X+4sTVF0ScWrxFDdFRKz1dJUKjNqZLLK6etZ/8gPYTqRKJSFjW1jcDvqrTkYmh0Oo6mJrluduiow
qFaEt3bG/FOnuZRpZeav5Elu0pH9HwgWJTRhhw22nOlIoSaPvRlsqwZYL/6nhqDdSMCJUUt84HSE
CSPsmAAnv7UAas9U14Korko+fjvEYE1NFhIfBxow0Xt0O4gV01+y2ycitogXurY4vpCvPTk7RHmd
yXRQF3P0KkNg9s4B3C+5YQCl355IsZYmP/yL+KerQPfS4TIZkw7WXX6U1sbtrwDehCr2CfcLK3y4
3RilPGXVkltPsnTWk8jQ2MP+TrfPN5C6FusLiMEIMy6eWvDx3mbmBEDMToyYgwYorjfT4+NGXuNs
y3TJu5ksRAosRwQPjDFKghEPD3EeK7Xh7eGHzOjzoZYe+kvoyJbzOoQz6/Nkm1bjjATcRcUqVn+0
nm/wTth31QacwF8LBJ2m4/Xmdr1JWf+qHb2tWNdjecfqmVtBtGRVUnqAqY3rrw1/OXIY1wSN9SfE
E7wyyV06CTY7fm7zzDDqOW+In55QGQF4kYJbwlpH2b2wnOuCkTX7Jb8NsHEV6xpxvF0tbBsdu0iU
8N5tnxEFJ15BOhmg8U0Tw09keGvSHRhBCp9FOsPE076cWI41OIASAutCs2n08BMXVzu1zNv7p91a
LKRJKKK5om3CdQ6jpuefjf6mKCyBWlzCAGqP/XJdmBWMP5INPOYFlUXbVoGF1qRIQVCD6JH9MU1p
tzM+xpqTcXkgatoOpAeSp1GzmV0MCtIyLywxgERvxBnj0HQV1SGKxP8iKXFFCclLu65AFymix5/J
xelafCkFj5QwdSKQLuPSv2+bCx0HIxCgCbGsvWdSVnr2lLl+egmXnKWrBBroDj8J6U0MhFpo/vwu
KNikGJkNjIlkuuLSFIaEv8Yo7zrhlnrmAwY9egmGBIbITksicQT4GkBlZaMWLZbBdzvlGu191sQi
1OKfvD6eprsNp+i7NxBQkU0CgVC7VgRuFqXBJ1cbStC5TniCrYtBuA731qX0WNpgQh4PUblQhPc1
7OuwCOnXHGBz0V9fLjscNetb7EbdHvUN+sTAILRtKPN18cIhkJJZ8iNdZfc7ksfBf4gY6bmCNBl6
tkfusmZ1kHI8ejMgF6Fm1uNTuGM75tECLSU+rv+kxfRQyNiODw4LCHQD00gy2RpD0l9HiR1aI0ZV
p0TjdwAXuFv3Y5VvRaOgWaFTj34fI5Cdlc6fA+j2411ntGu/fVUKunCVR4zzRCBjNGEohsrK+9U+
/ykg2hwxEqp8tr5dsqi1cTKaqirittTyg+KFcF1gGf5SABm6ksQ5EW9HvuR/REBT9aUMMas4RLgl
cGK7PSFkOK2ckx3RJN+eClGT1kuxHWSvMXYbRSZxtVkMl9/6nl29a9EAVs0JmT2Qf/yMXgWimmb0
3+Thm2SoY9Ra0U8YEFtGMq34P+y587Jj7fuM1cv14RqbHAJ36iG+AMygjCZYukIno4u36GJGDwLg
v/Qe/vfamjMkDxYvybv/gGHh5Kw1LG/Q6qeeLiHoIs2CBxObjDqOE9PAZYHjlWaALu3uJxP4QzZ3
HoeDDOx094ohjMIrrIRy4W4UDtg6wfvAzrpmHkckod0v+rncTUgMQZ8URLp1fCm+oxclLS4z0K3t
+62G8trEf0aj1qpbUUzgO0efI3hbl3xzDEjJHNbEqlyrH5WbbRTZNgbAEV0UyXg4ngLQLbPgAnKP
ueLKaI2svl6DhHZYlfHo8k9qV1xiOt4a0ewF17ZNUIYfgiNvn/4fT6y+DWol/7PMg2XheULgfEVH
pArpKEm8wojz0r2A1ywjmvnLoLRs8MfmOmGHzmMtzhABq3NQp1+bAvlNZdif+fT0u9HCOk9U9F0f
xtXpyqB7Tb5EweSYoYaYiaLoC6elm6j/AX/7aDdrwE+TyAYtht9C+Qrt+z1+R33RIzFNuuiBVUhh
CiyxtiPwvA6kEZnXSYj2iY6CM7E7NdHp59Vc6EHjjxfh7N1GbVCmPqd2KAZ1gI3xEXgvHCQvEOYQ
jjdkDIPFJ2iZnHJ0wGbyPekjfXT7DzjWfXrAkNwxqlQ33l9lbXF4QFbrR34+pMJpag4zj4Ou67Ek
jJbp92Dy4MGWyd+NjytCqmb8qeNmq4xz+SKwLuiTzDIkOhwiY34a3Qf4V6LlHBhYu0uQ7XlxldzO
b+XoWdmu7gjf/lBH4uOYW21Vf6PpBFFoSNg0IiPHyHqqOcGOtd0SPPRyYkktHT7vtJ7XLncv8GXl
yVb7IstwXx7/wu7RT3m/rDpRjK7bIkb/1BdxX60J4RI36K/gdnLoK8bPLZVJIuPaf+M3bzehzUYd
nRqajKVlnyzWpnoQCrrVoZlpRWMFjAwnTc/EFFJlSmI7hUWit3e0i8585mVtPq75LVBgwXkX27it
vGAUs/WkXHvNTjdJgXEC8SOf5pfC77pa5wDGZ2XDiUurzj1mT5X1li5Xm/M/l8K1dtqgJ4E8Z8uz
xRo0MVINIsnpiIeETjKDx3bjp85/OSypV29EaLopJZ/QkhIoVJAXdHS8a317tKZkz1oUCm1y6fjz
Y62zxG+3PiTyI4l8kY9+WnoxgAkPc/9oH2fGY13lgu3dn4ELWj2Ryra3HISeA8JAOJDcBZ0MVq2p
eNG8Kzi7LBM7+RTTIPwIiCH4YJFV5WSpeLwe0NzfF/MG7cpHjrcJH1fbVVlu+/lenh2R9iaMy1Eg
NMnVRUUiIEkYcvlxi+3wEvZWizljBVD8gd36Hie8zi1FZydtVz2TJLspwQgzATf8b1GTao2vKF7C
jm4BVxm+oxr8rPVNdQ2VQD8LDGd9doMsZqWGt+8HFMWMtkDvchyLUUI4Fg1DMhgo6X/2viVuFwOa
qPSz0CJ92YP2YzOTKl5tJdGOGnNyDFE9xoamfYP2afFB3kBq6w+1/eA2l+Z930rDx4QAU1mFlUvU
dGdSoygspIkLr2oovpXynPy4t3a+yavKLJDWfmYBb2Z2tvcLLxawkIeiWwjenHL02rxncljqN3vp
EP1WVIw9ApCpRXpt19XAf+oxWkbRQRzJutcEZFK1JID7YN0GCq3cr5z173v2c4KfbQlYGd2m7rWd
NEOPUloTAvEP1J/difuXaw5X9Lw8BLtVVArmId9D90wlRWFUjFoOpDVGeQf50sKY6y/aP2CmJhPn
s80HVODroLCo2KuYTtuFs437nIx6GfFhY6Du8QL+FXqc9nj+H1tBtrSivlmW/NHV+YynRnt101l7
sXlCgzVTCI850qiBb08p7gcmzN7QIrYz1xSeRJKIF/2PZQ6liABvx9AT1+tJiLh2vV8X/UKG4/y2
zVPeYMre9wsxk28tDjAtj4xGGQzHdp1baYL41R/I8JCnpkQnIZYKnUiTanlT7iJAaHvvMGL+KmMf
/D+ZVidCvXU+D5fmKaATlcE1oat4OLu39DG1xkRd3M2xgQZJuvdK5UsUgEn3Ixvh/Uru9jk7PMhm
OlxLSKkonqIhuAkvg7gCCusUNlqKrcFSv5nDPHU4ZM6Sm+9H/m0K0BjH2HKhKLZHRDm9tbSWhY4e
GPAId/Gr4O3xDjSFkVkXeveeQEeEo1iqjgGdOEc5IaWWROVAOLotOwgzC4T0QY97K4FlGmuHDukN
W5sOETPUAQ9eR79pMXDaeld1wp/WtCwvlmNYzVDd1xyvDy6K4bCjj4aPfiVkL3ynwSKSTcQH6Bdn
ttCt8vRV0CLRsmkeLtJJhNT4kOg3WInAg10rbOVLfYPFk/ImYtS6Mj0HLrV9ns/54b0/Pi0nX+Hw
90qJDrfIoCMDKngchghi0FMdPE9ui9fjA5n7UFL9zfI4LVRVkG6XWe/XQULhKcJUyWYoGn0vMhe0
Wv0CyOU8y+Oyscy6Zjl2Bfx5g/eVztShmIbNOvVle8BLangTXQ2HPDEAWs8y1KPjcl6w2IPoxKl4
XjbyTAWYQM5/WSDvrMt8AGIoJy1yEOnEiAWC+RHG9izu8o/LgPJI3aX9pwt5jmMqaqzDXA2oZbfT
hoinDRJexLTwDTbd0iiYvCV8tXkRk73ehDI93Dqzv5+5K8gNfn0vyL92gCPsssAF7ZTMZUNNbiuR
Qef8+VfdWI/KNcz/cXcRb+pEpbvWrIFabDTiFBhvCmm/z7dlo8CJQS/lUsVYJT6Tw3pr1zn5QpGE
5JbkFwQLC90NxfY7GiYGJ/3aU6I01hmqGMu2vT+62uuelBV0GikXqTNDN6LCM3Yg+KRrVetXaUdB
kAO9PAbYndlJDeIZFX+4GW8vuIbFtjNUSaQfL91RU1zkN3g6e3ys9NUjUTM3FIVtOfXQm5pMuZMK
oKYZUf43Wkie0OkQ/vzT8m4hBj43FSjnXLIpYpoQEyoN+kMYeHhTxk4gvSwMl1a4FOBqAyzXU2Pt
uxlDvDLNZPaXSLOzrgtwTDebau7RUh/3G8Wu0gXCLcgLyYyjif0LLsn2Db/cfnpdwb5ubWN4jXAH
9SCB1pVNx9O9vLnEkj3X7pel8Qa31o0ryj3RjjrgELnnJ9tLM5sdp/CiPd9YuMXixUgAzgiQ2znJ
Ef9jkyojO5/kO+fuuwtKAuJNF3W1mGp4xNcWFBR3vErHPkfg6x8VHmZ8hI/Zz2Gx38+MB3F3VT19
9k9iJLT7rrYYH222TdcSBFgxeCZuAtBWy3FF3PlMxp7Y2ofArrmRUG9vXv2H7sMb73gyxfbglt0t
FXd/b3rhcQbGjWMc3X0lbVUVo8ROk6yBL64TlWnBilgEJ4yu4FebbvNr/kTRwSBgKs5QdArGrCCf
OW3BFng7dGgZxBCy4Vy19E/pXncUM+DTGHxkDnZkSmXcWsgJUdX78izFzVGDbYa2cM/XV2IGgy14
p8EFiiq9mrzfWUeX9jttdt6poZZWybrv55/2Frmzca/fQ7ulHGbHp6Wb/RsyUjDqN7cty2JZF8FK
LaMIRj47En7SH3NfZy62RjaKY9MhlHVnDcHvoAFojntqUn4x24sOBDUMC2VGggDOIHyC1kKNN74A
Ps87THnDfqsrGHkXnSHmfeQLly6nAGZ+4aYSXr2eF4Vf6LXh+EMklDQAx077HrZ0OwoZJ+kkPjKp
fvKmjW0/PN3CFTrv6mmGeRRd0r27ycEQ+HOD596N3VbpoRFCuHwAOGp5c73zpqL46xmaXO/chqGu
heSVVw1s93Sns6gnc2hhc+3p0JNyVcORMnlT4ZCg6OPceNu4yc+lmfZnAhP779SlI9Bvjv0UKA0g
G1IZmFvQYN0T/iDIl7nviOQ6TBZk/Ifnipl523m+w0CZPKU409SJ72/TSRHNRWuc9W31xOdr1siH
uIq3Mb+jAhnRIJD1PM2fKtKrpe4TG0usoFWvKXAsFXs9gOfjs0MfEc35WscliiyP1S23YZQBldmc
FbOu9oOgJBgxjOssJC4aEMi1k0DGNbyT4xqE53m03XnqPZ25lFAmbLfJJj4oBmSEZpR07pgx1Hxx
cB75jXEMzjkm3uFmDdML5QIvuP1QUsMS5viLr67RKFL4bxz/vemwPnvWPH2DrfbqiOCkK98MwsIH
ITsW3wZqtOoY6SqK3hhTvfopDN7XcSDoOP3cf9koimv76j4yBt1Pk3K5raKeEbA7nqVZxpIbc9Vt
C2UPWgzNXAB13ykMoo/O/JV0ZGRLrdYOxotQjEkx3qPFmgoIDjBUQdSm/m11LtifKR/pC4MwODVN
LACvawTYCIrZSv7j9h0cFE1Y+0Bt90XqdhxpDWw9kyweMIoCjG6KuYl1fWyP01ACSN/PqH+mMiQQ
5cjnPnBFlkAE7jOXl5DTzeGsUdTf5gYY8OxM+UafzZRb43D608t/uVM9YXqeXxJ10QtvCMrvsVJW
FIf6AplRMNCoVfNVWVWwq+dAg30g6Uhqiwr2NdO0xANtCg67js/oqF6cqfimR3EpDyX6Gj+o4OWX
FRfraq0aaYwFwVQJVhW6TvkpvLEfBoeQGNy1rZJvfGUbcu7C9pyp/MTovtrlyvXUz6pPyYAmauO4
e0WlKczD0r7vykzrDxMyX84KEzGq11B05HCXFGwNuiv2jLfgtUDr8ASqHYdCQ/GcouGaWNfjQZ6I
Pz+CZBbqeEgXtdEHinhnfRtQ7nhYBtJYIyBYyhbPRH8tWO6+uGsluaXOUFHy9907CAERSwKhaufe
rJ5L7PJ3iZszwhkCRhJS5YuGMWGs+z8XwAiNOqPoMmT0iT3wvPVwZaGU6cLVVCHtLXR/vwMiFM1D
ZYibaHQNIv1USuZA+x0TTPywsRXnpkweByJbQzuH+Bn/T7qpucZKusw7sx9H8HNXjnTBHc5KazN2
FHuVBkUltGZNaOnTbW9z+sO8Mt9qtfJ0UguThXwaXF9NcWZrihztkehltWIqm8MDrVvMxBOKT968
XhYH2/jlboSls3+i4q2CEOvc3R0XLioHRBUmyrhpyAAGf2gpKedmpUu8t9jOZxlEMQRyI6WRRgVI
cpRb4NYdCrKRWuzFfr1ZctYMu5+ryxJaAbxxXbm/D5oaGHkjiQvfDZ1RfMUlHZJQXij5pQScHUyr
IUbNjbEoXxI7h1LKu4y04/6IzSfge++Cb0sI9Y7jgCZ5f6cxv+Wtte8l9WsDxOXVkuv3gJySBZ9Y
/ULWunp24L32MSfJrKF/dVPRtY5WcvD31bN3+tA3wDsA58l+fQZkLAbnXjKMBffegF5jhhu51CPJ
L1XzFrKluFNdK5yLM5k4CLRezNLIZbySFIt/4A3SPLOzCD11M4Q3kGzRGTSFFnr3xLoVUcALO9GY
PsVCwfaUxGfW1Cah/YjHYUC0SWu5A2SWceJ94hg6f/Xq3iCohLnVOc91uux64MzfZolyHoXKsUgr
sC88RqJJ9QxX1KhWHTdE0TJT/YArxonYEc79VqS3O8bDvCUxEchZgLKBoTW8p6Li87pYx+MKzrnw
J4wbXBvoUfDDqjv3GfJaJkTd5YrKCBy73kb3cU6kmbt+x9X6CwG+by0i/6xqHFcGsGPeM8dSACwy
rx8vxY2IcyAkTzpQMZBxR39olBasgJgbDklt6LH7+lq0txN4e8uASOgwfDF8JhooX95Y+MWlp0hs
tYHRBjEZ6aQ36j4KKXifoMTOGRgU2EiK3O/bjZresnedNBV9D0ObGGLTGG4AfgaEIUCwvBL9qJYR
2znIh47pGaKdWZQu21xPEsMc3/Q0US8Upu9NWehRnGr8JsTfW7MZaJRemHdbYDtfGVfhoN8OR2d1
1nbaP1x910sixeru3bxlCebwUgPEZ96yctqslJf+Kkq8dQzOc6goYzkyOa9Ym1kjXecmqGexHMU1
tFIZSZgQsgoozjGOQwdzsBC9xdZ/xAWM+S2FqqBfCdAG2Oa8JGMZbwbnLTXMU1uUAirMzeOeT6/s
xwowCoj5maC0/IETmvxTqfZah/1jrNcuJa2LzMMmx7WYUc/a/IJ25IZZUuMWzxJT+8LI6YGEWeJh
FMY/4/UAGVGVx/zk85jLKSeWyh5I8ZjQOMzovUbqCdbx32hnxOEYxvwR6b6+Ze2Mnso++p6RenOo
5yfAXuIj9zw6jtURJg2561BdFebIbPCg7ytYaqHufoXHf74AEgFOVmqqRRczXvV3J1W09JU7jxac
65qvHCxTDvHfx8p06zkpoQ2sOyQ3NMplGqF6p0PgJPCb9BRW6ls/vTRLeeEKr0JZrbHfY8KEQyje
BZNlW9TB9gNyBBhpre/zo2BNKYeIkW0j9IoqCUnsvZ+U8VvqMorXeDWz/+y/6CkHrgbElm28tniL
vKCj1lYPq2GGNdLle6dfxGzJU6m4F6ClfnoaiZtwBgBXiq/gO7/wDNcygTGDFKIZTZvPVyG62QOL
TvbAhRan3/M0EMNNQCienxCUtjSodfneVEEjktM2XAIF1j0KyeaYbU2RksYE6O1Zj9UQqJ3vZEyI
AY5/HRK8ULqUO6Wg4/uKfl/JyWsfnzdxWLjiCWq6VbJNyLti416F76dXkkgDcJPD4+TSFeKot6gs
GDBNWf5W8C8eddjDhbfxL9sqHBXsv1ZDmX139UGb8+4CX0+tXThiAAis06wrvkVdRM5heuMb4Vyd
bYJb1HVuN4AYJ58fqK7/wJCHy0K/zs5Avus4oyAoRF63cZNJy0kBdGoxLRzZL8twi2ar8AyIu9v5
Z3QUZHo8sP/8CX2riZf9fQ4z4O1l9JWIstKr7x6NGMgEdsEKk3uF0cQJIAX7j6qC5heQMjxNnVGK
KR0okcVZdSXv+CnweVjDtr4MYyDFPhCWGZOkGr382afTdNGHP1sZnVOU1ncJauV8IZMZ/MuUC1JB
Zq1pM49q8YnQSFMxd+rnDssuancgwhSarwWXIdrio3twex2lBQHQIFs0JCxK2waYgMlZBj7b8YE0
6eG7Fqsl7BDNKEyVNbhsC9r+oXXttTOpBPgO8mNCbYHApnTTgxgPF3EULEWqL1ZHzPByYZi1TkWK
cPFWZzT1d4G0Eq0IfzRQPHue28ZwX7nS9AR/ZVUvAFBLyew0/Yc3hbZ+fJb30dNo/T4+3sLVs+Ou
9P+Jq0Bf+Nls6QlbjgZewTd7x26shU5eA3JH7eXFkq219BJHSIa2Wp0d5Yk1jCMhr/uf8mU9Bj4Y
sM2S6oTgp67Kb37dWCZFnMnLKCoY3MhiV2Qa1UMKKe6Nb4dqm+R1iAzDWQsy2DNrL2rb5AHtqtQj
acabtK4xS1Kp0O5AoEp7FfMN65gRsu64VuGu9rJd/FNhq7R6m44m/Ub1QrjWLFsaz1JMf+BqhT2u
6YXLuI+xq1Nh/YynTShrEOLbnii/HKMskTdPNlzjY3E9yBPv3SdvqgMhT6LDjazFLHjhs4GtCRA9
fJxbjJkdzydcirr3CGm+vWIIGavj07FMw2eT4mdpbeihpoxFmQ6qbjaO26txbJSOaUChmEHfyDpj
laJbbp394RmlXnXzdk9uvbuw150M/mjAOnvPvQclJjQg0c6IG67077rdORCyNmcdHSQwpur6yg5B
gHe/cezIKRUpn+aX3INTurXmoG7+m2TEwAINqkklve2Rp/KBupENh5cMPX2mR33PoqgPfqbnYWAj
Ke84sGOrRAFUFjucpVdrRJ6blgMSrWocJA9v5+hUG3gFQYrSe+A4Ac4ctV2cUyL/Yt0ga16ZzieC
leNkJbRxmRt5UlxAEOaVI2XoNRoZJ6UkX5NsTkOiTUsTOU/T/AAq2jy1gUF2wOi+KbRLTOclAz7t
s6cSs8kGgZmrRfaD7NQbx6XwNzkRNIff/zxp01Khj1pJ4VR41bUKt9l2A7IjSwKZTH6GWE+oThCI
TFCdZL6tuLNvpnvqK0wg8Sbyk7UzlpMoQOsp0bkqDhfCWsn4coO/PQuYZvFIMPY23jldA3xSN5MB
e6xgZI0lqRdqq3SThUoxCV4Jc2FDdrzB42QZfFkUGgHQHIb64zSJ6Yh4F9Vm3LWFtUIzEjMNxXME
G+gKVF6ph9QQz8AK1pFVer85x3KXy+pHSxQPIUxRpUb1P49vZ8Xq1ThULJfXyBM3f3NVQy+4fepO
t8YKjKdINjgIMD2UOoNWZWhB+fhlhzJ6GzfHmP5azb/LZeNT/Y6s3TTjTd3k0Y/o2zo2R15C+f+m
ye0brFnjKkP7WxsxQWIKEM9fyOkw7dcT8fWnlXsvdugsmMLjUxS7PIS0av/vWBfoJ61LjLm8QcTE
hHFLJyuQE2ZxfttX/WNEirNTVzNQ6aPeIsIiVKaOYv3xd50a+dssc1Mk3Pi74TdkWJfIPCdXvq2g
BLdMsGoiFmV1DJlrqmOAkn2wkNv3gC5Dnn+YihAMq/Lv9ZCplFBrTTTTftPV+R81r+EEqIbRfRaF
a4BrsyyWw9EJK9PCWlu81LZPxtKrBz2h6pOTmjDe95BVinbML3Xr6JYg28hz8cw/XPWTvQ2w37ck
jEuYfd3lQL0P7hQGco9sL7YudwW8RIAMcSckGJEOaJgJVKLpXitvWRTpTIJrqpCS0tQ8MwzknIrW
KCXzdqHfetYhh7dAfZxjgEP5rJE0FkFvP7a6VHPlHJFXm0rXgIIP0VbcBSl9fJ04pr36F+84GiRs
Lq2R5YRKeZkut7hC7TIjpzQcwr55bXwhwwu+CSfl5NBRT0f8ELeLYuwZLlf4HkHHU/N08XNRzmew
oQyeUWPWOAG3sc/9sWCjTr8mr4ZWpaEr6KB06/KWUTbB4qGjJ3BxEk+zQfWKAno0Xw1MWEoeiOo1
wR8sUkdXWTPM5QUpAPsx5clO5M1bOF9tiGaeAh7SWl7h33/aAlSmJGNzIi85Zi2RW1qlhGpTtuwa
TpmKuYcBjhyRlt85ouPxJvckKRtWTh37gQQ+vzbVSL6WyyHyS+slmDvO+yxDZpOFOnnn8vZcru8o
pHkENHSYWNyk75j4wR/gP4IsNhz88gyTxa9WoFyu5x4dlrxHRfpWgNTvA0ihCSAGdRTD7kVcOhpb
/Dir/rDJ6/DRoqkcw3rf6l+NRGhgOwaGYija1gPiJL7NWlZiTP5Tj/CPHmMHsllS4u4hPe1ID/PE
/djXHd7NjQRoYxE/x4v1pYEl7uOY9hZj8g8Sq9mOEC+3Jqk9G/uBi6RTaB0TN97opNvkU4lvjPFh
NqA3HYz2wy+wt5sbFoHHpev/QDhhMun7mjFMrvPue/0y+QBR99nOQd7sUs2VziBO+rBvQ56Fzutd
rf3/1JatM8e1mQHyGIfp1J0ymuYLRVmEZawUhnPzjIqlYADAbY4HNEBa5r/lbZCfQzKdina+UOuq
RNRm/5xAqWBtiaW0Llx4cFON9aCkZ6YLbMH6rLUmxAD50z2uE7aGjsqhQrNUsS+dkj4g6UfGK75U
+kXx74rsAo7k+YBa+anY8Jl3ZjGio8GiuaXlgZF7ycrDf3vbgh01NQKxddLZiFbCjd/RM2HmuuwP
t0V6ZRKwSULPfKisUNwxE+GUEhOM3iEr4mTJzeQbapfNLb7gIroPBeQJqWDouhb2ZZOtxZGD5kYM
dOpGWoyohXmNnm7IAvQnFCPi2B8SNOrBEFZJtf2VjICORexAiUnZ+65G1mAlLwgnEAfy1FRU1Wrw
AJuYR/P0N9Zy8cfSV729mlEi6qZFVOI/KgisJSQ7lnVziGSmoQOUqaKCyZ3RXkTMYxVwyV1/yf8v
RwH/koEj36BGKLCVZnJl+cQnn1kDEQHQn0m/qFDf11vQ+SUfB2Bz5IrTEr70aYh5IDJHjn2IqXKK
NSgEj0dNSHFn0w4W4AHJrm0ZF0lzNsk69g89L2ydAzH1/JqBJRw2YqNuvq0Cz+ZirI1w2hOMPCX7
d0g+js5DesWSXaS7+DsUbinUORwGJwms/58fSIoc8k1la0Jzy2nX7Jx0H93ZHuPQXHd75tVo+ckv
KWBRMNlIy+DOOPrDfSMhBxEjn9nvRXLHVhwxH5z/bx0wWF9GkWyoVjZ/co6gyOTM3WtJG3u6R6Zr
1fDnsuxGoPKD7DCMCuyf2oRxWpBeTPNDmb9YRS0YCiscZf/acgPxAili5zf9wl4droWplhqW7f2b
166oU+XvZrV144CWYwJ0Swgf4zuUkLNqVD9ods4kHIJaeKYiw5YQUXy3Jj5NliU7cbENTLuEJtCd
GXo9Dkf1pf6T3QJx5oWb0cZJ6ehvCmd5XOiOd9fq4R0GZFu4K9MfDzpIsaoe0YZ1foNF8Fj9G266
qJ6APHqjB7YzkcqrMQD5VZs+kM4M2B3xg0nIsF3FyWzLnuoZDzl7OEJsA7hIw7CDr4rqlv5/QhUE
hNfnfE2T0HFmZY1HgaAqxOZD8XPMePaDLH4tsn+kcn4EUCEhna/60YFHFwyjvqMPt5C3R2o4yNfc
DxX4dp+Tb1rJQkTX1l7uctrb4uuHMG0SgRGTqKZ1kkBJIjTEmOJFag9acXGoibEsUBqMo5FZvKpn
U/5B++pD0is54bhpMew+6D0d8Pu3fOCywhDJ/IKcdwn8u5Y3EgeJRl6J0EZq3oiCLAhl7JylZYUo
mXlI91NABneJswBDmc79Rb2v+hwdrWtXuBLF3PVteYrrEZbiS0tHreNA5Wl/5cuc6MEtMYSwSRGf
1yx3Q46mmwLX6Ij0KxTFMSOHbgUdALJfuSOnFNQ5Kor0YAlXnkSqUbRe8fXrVxU9jompLuAJFWb3
JEgSuOMEGb7nA1MQOCfqPUXFG1c3G2kT4+hc8ELvfgAkic34faB+IB5J7USw6tI3Z704jY2JTTvG
wCnzTv0BRDGhSN3POxQtpqccJISvRvUePaXvY1ANCADurN1GubetRv3r8kDs2MamY0ztDpNoqRwU
J+QjYw7o3JSi/7JgunuHJWojdbZLMwkCVEcEEDPxpPeWbZ5JAGU8MZjjDlqD2sTMSy57BB0036hv
c4/dPi6cK8OYGqMpXv+6oklm7VL2PitrAPxNtUt+Wx0iLfxnqSlO1k72XAURR1XbD0gsZdv3aBK+
3dMvGb4DGV1e1+fylrAUEsACpbCq0d05srNCNX4dl1lr7rV2oFMln1RULQJeAv/qqrd4tyIe5L/1
FQJP0vKuE9wNTW6AWKtHY8JM1oAlj1KoZl/GerEWLkjFMh4my01c+SlWxL5MPxjhLNPQ1FRdaXme
iSTEimhpllZlDsmK+NZoSN7C495bLw0Af5XAk9Ia1n6wgynOEocnNBsFo4diGPCF9W45Ld+EUGaJ
DP4F2/fEbggZ+HxLfFWtDOp/jGAzOAYHpTs4+Q0RqYp00sThWFFlAdqk3OJEqljue6bYjvMQL6tF
WTmAlJ6BZjSHasDBt1DgjpQGr2iQxdvEO8jESOB14Gc96MeM5T1KWvqjY58OYgahgPvYeYrmSq8T
xmEd7eVNB5eA1aIN12aFtI6B/I+DYJsQ3auf103nZ8RpMZINn3xWRud0824HDLHg07S5wgb54hv1
zFwEeflxBnh84UViSV8k3eYNL07mvCvC3en0nl2ZuhevccufVacX0yW7kYAtyrA6Pu82Mamr3+cc
ZcqdGmpUsQBgjh4lhY31MVAFrQ/l9h4itdzBTrqrOf2Ywl+Fk8Xk1WvZqOvRP8eZ5BQXdWJlnGXF
kTXU2cJg7WofiK6jkI+UjMEJsB58kc96jt/68n0HpB1OCcnoTMjwI24VWcH/61I1W7FG8g/aS0dU
e8aSoqMNwF6gO69qAzZgQzVvCfb9hdUCPxj0dCrs43qHSgss24cTCl0pBnEh6GA+XUNTms5vE+qf
BE48K10xhdXcSnXj7FXlXEJPe5w1Vvytm9fWMUz93PP8KdGH0QNHWtmiwzNDTCx3FpZsiqhofVUu
6spO4gHPKF6rQu/H/9e6Q8lI8WAOsiKo1rssr88cfTp6drurgEgv/HQyEI4pYeMJ0yn+YASsdKqZ
SZgDB8puEAnyKmoTFhBsEwHOhqKuJpbJxVMqu1C0nH5k9iuLo4PA8aJEXbZ50wlArvlYdS+NJjOg
E8kvYDIpcAozbP7lKmXJ7MY6k9VeM4kOvJsjH7yGLvolYrQaQuQQbt+TgOD62YE+5qq9fv5Ndv/B
DNM+P7i31Kw7s+K0p/KG55ieb+nCAdiSBV9bJGjQmAdHeX3JCZmreFsHkbcom5jG1OMjy7NYzzEZ
HAOnfT4ST4TvXWyvj/TDaWgV+cn2yH1hqNZ6imisrAjg5MSGm1K7K8GfvDPwtyvVDkdS0+g3cUr2
1Et1fBi5EIGyf7TSs34A+AYrut7vCF8tNMvpjZjfQq25Ix1WrZXandEGNddl978630DuNEDHfV8j
XJssrO5Pi+NcJUDJ0bpYbn3GjrxPz1DZYNqB5J9vzNcGUEPMJXb3xst4tSMMI0yP3tA+PfZLFVp5
h90uMCDfAmC5NX30sZRKRpKfq95B5RbS2gEJbvJUjlP8eEvm/JkjVZqcKZLO427gJK18xKzDciDG
UmA3fhHaHPsnkJXZ2A+WQJgyB4pfaNacai64I6bHVV2RvtBff34jFGAJsAPzQABubV7LQsigs4Fl
RpUXB9OoZNluYYc/yCQjJ396WjeO9EUH0WIs7eO6Z204LqrxY3GCEJLERIYUILW9BI1mp+3Dtjti
i6Yvl9GwmB/ei6LAXQnhTkPNHp4LGJV6dtFYrtygyjDhVRGgRuSzDIhQlo7Ctm/nUtRNX3O8U2Cd
0Tq1V9fCB1J6C70GycovMMQ2VJCUk3iEXLbyAygPqlX0lTqVo/VrukEWooiG7aACWXTQkYe/T29a
8h8m0HuhZ1I/c002ATgEM7hhJiJi+o3bQUspOUxG5YFPAAAtc77wJNJNyIv9Lbib8Xy/yLKJIANK
XrJu79ueqUdtk8JPg38V2kGwXg2kVqQyWU6902JqCEVdQV5Erhl2UltO6GHjyYAhdl8vsFESDdCa
pqVyCqxmgJV/vJoNIzfs0YNVdrUh7QLFzq1XI8QcEP48liYqqtuHv8gRvKodk2a5ha9TtcM4zzrH
ENePEjVkSPr4OBar1/EOQjEMKICynt9/M15Cxgh8ljQ+r/ySOuVvKUGFWX+qcyRC7UpXoll6Cj0U
pSwGbNaJ1u+KxotGhqdJ2vkZEbB2QthNXfYYIOme+9EADnjY2IO8XA/QbQgx29GyYp1/EeCEh7fu
e0liI6HtpWtfuyVJ76OPNrMTD9CZMV/B3pmpTydfVhL5ASUjEpzRpCqH2ja942PJdkVBRi9j5V9U
9wMKYKoWedaddQ5b7Ad/Wk0uvFvwHd/Lz5I1Yn+YfO2xzwYi/iVgu/AwmkfFPg7f94L6K0l5/egz
O/fxnRf5zbG2dbUT4tF0hPcvgXI3toe611PZ/z6bUvO83SUspHY/dGYBoeBKu4WwXZbUv89IVOML
OCUym+HrQ9vBGrxHK+zfYzqQj0fBJinoZ64AucA2Vqz32PL1AWHM02iwNZZ5BWXuU1Mt2/mmoLlK
mA5uSMAnzD8oPt+pLzpr9kK0zcxxXRwpGrPvndKBuO5+SLtgLuk9gt2oLcZ8Arje/K4Wo1wOhoYv
EyfwzLzSFWnmnh5jIXJswzeq4G+ZRVBIbhkN+8FNi9A2A6BFtW/Z6uvxOoMbJdD6knaALvu6tpP6
yKPqYmJOibwzL/l3vWC9nIUhCaGLNADYNdUAZ4mlRUgi/7AEk8SkBtM6A3p/Yk/DPBWS5UvIdEKR
pBYxVyuVUbuhcdmYOm/HTxI7HN3tRVP7FaRcAAlfOAYwVMMkmMYnETLWwOvBlKqGvKSxO+EpmxsU
s+31xVdJLEjgrRaiUW320cqlXQrM1fpiprCWZKfHJqrKGLeiz7KmklcAhAJufN97SyE2X0xJaz1p
7VyLozaEtwdQxVAYWnGdsFz+Bv9mmjmkVTt/bGYkqmsQ8mlt4I4ySnCliMGNPRl7icW18udSEcGu
LmPJ6Y7JO/ebFC7dfyElQkbEDx04qlF8LCPqxp38q3ZdwBKl+1+Q+SdvwYN8bW5sv2jwumH+Kmy9
+PqP0dn/9iipEtx03/Yjypc+2gnosCMaFmzTMPFDZ5jIwO2H/QrdAjFNyEvAOR4ApRy6LhZMFq8B
ua6Vh9FfhV0IQ8s+CXy5jyN6z4c61POTWiMGt/SKuOj91B8sTJa5ZLGIcVO5ks/zYXXvBSB/v8BL
JUOSCtw+w8PspcqYlnOnfcr47pA/at+ZbcolAEFUUWX0mxST3VQ9UAQkxM2P9z87M0cLVTnnDXLO
Hcr2KInfLjlMVyuuXTxhuPDi5IRXAItzusKI0qdB7bG9VDEHEYO/5ledKnlqE+/NC3p01nnl/+QV
clwQNdBtyfmrEzKPfVfxjK9SmuT7ssYMORLFaxUnpOJFCZJK1lEq37wrg81Wnuyy9gVhkVnEyCPm
LyhFwUbPqdjwqbU3huOCoz6B+7qfgRCIs4O7BAbEglBwPm5ADN3UwWsfDfC5+YyhhGB8GRaxU815
hL242nrBqVOEanb3hC6BuEG084AQXiFp13v29y0wWdq0vF3SdJB077VFtYPtyHY59jAc1Nz6KB51
u9/2rc7eIM1Z+wWuuEvzoSMfFh2dl7TIBHYgti4ZaqCMj9RBiQB8r37lz1/yTkp48ZFBfV2MMygz
ph+0isK4NFd1aNrf7uMUFa1/xnLgpVbhZmaiblCDX9MFBjL9J+HCBASW+1e+cvVBhbbuNc615KOA
gdpfx8xjTGI3CgekFUihi/buVEKklVK1YMndwWciz1Am+DbAtkWrJXZeWMcaBGaGQOYOq/3Rtcne
8I74wA7MaQxp52i8mNhzFvwQ7UtimnKjyS3ZBgU3+8UbaYtZI9XQVvusPhzy/Yy5/0QMC/G9h9U3
hgx9hDGrw61BycuznWF7L+Iq4hVSj3Jz4FANor4uAinxciLArqjpkxrV6/c1sAaMFJ2CjKm4982r
hp0Q97HdxBu8tNhgxEP5t4H0+vkDq2RU7SMW1yeXjHWzdKtZIP3GtGLclpKnTiW0gI6UWuAmbd3s
y4rjTtlKZ907WRacwKM2Lw1L8p8jXHs0phnPB7gVQMIUh+ZN3lWRmAcFnAP50FhqbohkLP9WJxPE
ajUU4ZXh7h6vumQKkDFzOi62SLv/eq9jtsEBm9rdav/Aga+N+9wBmVz+0dHyG6OOMME3S6ndYWQw
3DAZdot+r7h97FG814kGNbfcD/POJvZ4Fy8hh+C2NeVKhPIX11jDMuODlU3fZHoIQbYzNcvmx1Wn
53g1IEUyVTIY+2sOMCaTauDsyne08Kesb6fyjjGkxTawMeBTKdjh+uP3VRnZNUdbidlWljCcHbhP
N83LfSf8wEBPGnmEW2xZVOmciE5Glkj4u+IVOD6u6M4lrxNxDnQSe9RkYkvBOflYzFhl9u5O1wyo
ClKm7zYuGK7PRCPyzlw/3RlTxpxe4ugSBl+fWZ5U7zaTqLSD9A8BcArGkcNpyqMo1UNdW75PMuoX
oTMOWGjbRvT+7ycZv+QaZbE+PVsyzJ5aX1O/Arsdk7OTlV//dUdGBV3Bdf2SP+X9jMlj8QSS0Pru
Tyt8WNp/TlA6N5x4R5qJno7cDWD2ObgRMQVlc0IoLwfp/2tGF/hTyILWM3P1EMWArnkOk0WyjfP5
cv6vYs1noaU18GnjZbXs9p63CG0v2ehsGqTKk9BqTufNXNNPO608d3HFq/+H4QQdQkFn89w0epIM
GeVije3jGBHFztsgHY9JUtgssSrCyMBy2VyhdFppdo4L4GF57RskdToRtiYiahN6zkC4MvcoNNzf
0CMt1IxjL74gGYnpYSU9kmfqEaGUh5dbI0po5qzaliMFmrScKliET/Hucxd/KU87dykdWUB/nUBI
XQnDnETWRrAzyA8UGrYIJQjw8koaYuvResYibfBPgoWtPg728xJL+lGE3WbxbfJnLjJhT2ee+zMQ
PvlFCi0QiwTXkOscsa3UGfWlg56ejU/4FKgGCEvAlNuupdMURcfXnr5jo6RpkluZY+RcZvSkTJA9
VlV4tgl14Os+EIp+AadEB1X19lzA7pS8UVuUKZ+Lzl2Pb7v38EeIH5kpFTvMv9WpVK0HdSj/9Ftz
fOaUK3D/Un7ggw88v1EAwwI0tBl7cDsOIcsmSmn5YxFRFypzZDF0rIzM4NJTW6WBxXECIIFe4wh1
cL+H9L+jFL7IhhJMJSdfmQX1Q0QVoOUSH9dgIVmLFEOAJ9OzYx0oHsQRrRzxtnlD1GpcAA9PM9w8
BDfIvWL66gRnQuvkBjgpATMyJXUA+tEP2KEencBkLJPnY7yVu6QUKkNorn/5Pxa6FZ+okz/h6/kN
TCH9JEaLYcQCo2Vha5rY6iU2Ft3uzWd6UBCnkHNV4ecetRLydORysAxRzNletLD6nzE4gtAyiYFB
XWZcXIsrGRQC/6nO5lNzihyMXTwCGJz1y82FQLVtTjQsYoPCSahZZqMeaxS/li7LPLNLd8q41Yih
0WvyWqdlCYpS3ZxMIy2oPizP+/3GtGOwK7wgj6aIDVXhhSghcHI8GXq3nIkFPLHVX7EShBsGe2Rt
58nz1SB78Qi4a+aM2UncZHUOF+fJef+Eikyfv8hgRXK0j6ndAKFTdGEgH8c0gnL1QpXN8QtA4pXr
fnS4o1uKASP7JJuH/8627MA2FTo/Y++fUItABPsgs98eg0/DP9wfkdyEGMOdfZ+yMyeEME2PaoDE
hXf3es+WCGb13IVALwiVZNIMTBwFSLarODnENmf7bO4brzZqO4SFosuDa+p24o90zDb64+9oiLh0
wTdxqtDMPbsFZ91hP+ucCsQJuPi3Zf1Lj5cl49a7bZgDBMghzd0YKXsA+aleeLR0TjBUzGppVIk2
TCresnBenRWLMfxIo+1r2fxNwKJA6fp3no4+aY9ugR/VpdSIEUiTeDD9l+wqt7BjGKfpWPwzRq3j
3ZxyrTnISfy0YFeXrylkU/SQGolpjN7+nPcwrywd4K5ccwZyauVhVunYlya04bP61QfoYvQtnzRQ
/2n57KXgc2OQxEZL+4/G5y+VveC2uXNuykz889GRodENewBF/vHu3KHhpIojlnjIf/S8hpdQez1z
sthwrxqAD85Wn8oFxY2jmgCS4iDeAtBq8zmmYA/R3+heS/poDiJPdnTuW00dfQX1zSxCOJtgTKZM
hfoPJvnJgRlNe0r0HDaNM1istzAtior9QBL3HZ8CSM4PTvj8MRls2ubPdVmFkQqkwV5yQoElvszI
n5d6P0Twj3pYAUlvh4UQhKd7WavJSRhMB9yxw6iSdqRZEPlI27pl3AkKRoce3lPSIiM5daXi56WQ
01DepHJczAhRhuwf06N3qYjzC2CX8maeNB/VJm0vcwdPZdwRZeWsunwymQvgYC0o289PKjENihzp
/OVTT2sG5FWII/4wZDlaAgTTK/WDmRJyj1H6orVD011opiZei+pr88G6lyB43RNBIrW8jZFpX+Ib
xYWpT5U4790U5miKTz4IWThwOvmg62hS8+DQ5uRjV0BYFi1nFMQ+pnqRpqJPbm9L9eW5up2mSEMl
Dy3X/snjwkMsbbVJSjNeIyjIAql6JrcGHeVc3OgERG0P741RYYoqUH+65bXmrzqA/l7OfVpapSsP
p5qkwd/oBUaZ2nJOva7wRVkMAd3W6tebuFvVA1qPPOZ7W1QdB/HrXzjzAbGUwmiPAoMWOJYu7VTx
m/jqVqrzTj4TPhdD7zwfklwmKcjuRF7EV8OwwHPPKmJ0yiKmheNOodkdQsgI2j5L619CoNQJBarX
mBEoVtXeVhftZKIZaotskvozYHLUJ7jGJ6Ah3zdnF4iRL+1X2rrLlzaRP57RHufmRhQ/xgaxy3mj
eY5q1mfQWAL2Dn0SU1UetRrAOYZdfPgFqvksxC1C1n+KNEDIxw44fgzl2adWsu0imksgiIRyPJrn
WTWTveRgB9+AeqEFnqP3eB8zohQv9+FMkrp1IgkzdscYM15Qn6o45gBRoc8+r3k323BDju7wABRf
Yshy+Fvz6cSlg4hhQKYbAv/nuj1Csai6EC9NhRyRFiC3pFKvXUD3QQ6nEYgkHg6V+8Dzz/r54a6c
FcfSJmbokwUmIsyI9sNXuKV3WVLHHFulxfsgfESpt98spOEYejnB6Y5f+YQ7hx2g2yF9DQIOoatw
3ZO1b7T0tdP6ByvvxC4ExzD1/m7nPYZ4baVWJ9IuRWMAAZ8/od4dh+fGIwBaJEdtmKK3wsx2D/Od
I2hAHkeKwMrragaAv+LAn+zmUADhAigJpGW8qth3dON5l+gAZNsb6Mw5wg8uh3OIxu/kP+fBMCly
adwIMOtbF/QG3oKBMCU0nxzNFdJ4EF9ubXvQuJAff2guJhOtwFlfDAq68nRh8Sdu7YxDr5gstEkb
KzfNvwn/2IBJ8DEi9IAh+8OXzHQUMdBqiCpqM0zjQdE6U1/5ylsD2Rf4Y4MquILKR8TvYrPuD7hf
BSF9bYsIy88f+Hw6A600Y5izbr77XJiOFX2rSOWsWKDrLdbMtH/Hgaz80eG9TWHO/ysf8zkjg3IA
PAZE8l0mUE20/WOhfe5mjZY9nPfBoEyDWHbAglBycvKdtLumxvBaF4ASl4ovI2SY0I3PLIoIXfV1
8X72tPwOKmjynL6l76OFxDcCG6oBJThgb7pqLGg1PAHcaqidtJqcejYo4driQGS1JJvLEdHo6IrL
0tqJZ6lTgoNSZlhIVWNPjeIs6lcI4zpkEGDt8vJ0HkFbYgU6Hk9N0IpRvE1lgiFs2abK1gqeMepT
M9VUH1iirX4jpoR5zJi7xlggWE5yCvPJ8lIDpIk6D7/E0ngsL6NdToItJ13Sree5HpbI6KyMKh6G
aKvIa8QU659e9Hw6NIsvQXBr/22ZSrNdEk3da/WqV+uNXfrH/UWspxKyHuZkdw0sl5nJM7cQ6dan
2GRFxlso0Hcr/1PSWYPUNtqDMP2TayqYVER4frHvvXtpVs2DiY98MN2gA9FfoadUxLaIkXgh4nVJ
vJL1zqrNO+khQ9D5eJnplaqCV8+L7M3gZq07UvYufqgBsva7Yo73b+hCt0qtGm/yMK+qNXanu4zd
ycziPX92K+8jDBNXY3fZLfT6f6MqSzFjb4CddlSKFiUy62skz/ag5AFnLkyMY5J+ScHK7i6Dt88J
qfrd4KuuWO7t5BBjJapZvN5jX+NXDV8rDNApnZc7mjxJkXh1VKBxZ/C+bzMupDVAwFkV2j4kIy+d
wjA60bDKmjSOzPDmJKW4xT0jlRir+RzlcPNIFd3+qT6IxMQyEjwL7D0KULeOdKCF4ZS9EQYPdNds
iP1shJt1CqFvm5nnf7LjqnpLet69o5kIuHxm6OBvf6SIdxJGqa7XnpO4ni44LECvqU7fyf/w5cdO
Te1vkkO9U/wknVynuLiVUituuOX6ltHjC4+YP6y2gaojaQNkebQRVsV+UfJ3LP7neNw3x4g3HWeV
dmxIEdLPAmdjrr7EIesI/aYNxf5kzT3MZhandiTecg9NsNosJipa/EWSmf8lD4LJrpnFSGDfvS1x
/1IXnXZysn67ZFm75UmRjCziL7jAM7JTGBO5QHJX29HDa+fVvUr6Q9JJ0N2Jm1ZG100NNY9+C2GB
nOvz3ndxHD67ne0XBtdFzzyygnl90MTQbPnkV/fFL+qu/rt/f2f1oa4jZA7I1gEr2KY7zyO6HUWl
IY00GbC3LZFkFtgxHyzYiSzb1EELdMioSmgzkfT19j4ZEByY+jd0+lVKYthpmxB+scutGy7OJl37
yIXwyAKpHm2pZzQ6bcpquO/1pZXmmadMr+BVS9MMS0SwQ102m8G7aGr1E1nnCvVPZUzMX7IQPzkC
QsuxtgRjsVqOJmGvKfxWeGjVGJOmF+OhxHgBdIlwSgMJQtKvyIixnEMhtCAdRUMxISlvr7v5sOGZ
ohUgP8Ghtohwc0GO96s9bAQfw9TdvfIkVjubSUNCnCtAiUeKVWHYu54S1XHjEJVrGg0lcAzt8WIA
z0/uz+GEhJZlL1gRbxP/yZeD9IdTi8fi5f8JgOBYTOfsLs/j6X8ep5wozMDOWo0wK+ZGQkCj8DDx
XO1BgjLwt50bXLoHMGaI91T0u2WcRzxUT5d2ke7P2aCYOiORIGbFV1qyKAqg/bQEe2cGVuhgIDtn
eGATb1BHXYVm03UGQfYtfkY/G1MVNKAQ3UdMfR1HyStE1rmM4lFWl8txk+jQu22uhjkeljDlkbg7
Mq5xqCNHQ2+7xM9NisT1/eb5mu0t7EtzqlY6ZPK1dT/Y+ycOgBKX4uRWBcXwJbTAWCN5R1FB9PTg
d2SaMbC+PD6YILCYpmYw5L6EAyAAk26ksH5T6bCx/6ojUfXzhJl6L5FF2vrCg1tkV0xbTsUCMPIO
aHAhnEIn6QbrTM5bZBrlrO7MNhQnQC+M+h5JpkqRdalvdgs/B59a+b/8yz+7RFMBpniAjtLLV9UU
0DI9RYQR5WZwy7NS3Bqc7IMIWdso2AjQELthJw6BIRO+RUsJT/LgvMupBvseW5ne6NmKenudOmNi
eHYGzPvExI3Eaiuh0bPmmqwX+hzUm4nq/a6IpOR59scHDqe7balxRXvCKsQt9r0RB13VKYxWntid
wF68D63tQVJQTjHnuC5qeOTYwLPo4+MSFk8J5oxSa+LXnxqhUGIXpIZa996UtHoMvWRlaCc+c+a6
v5cLCc8LGfENf6J1SOiRguw0giWpC/v1M+jEsw03Q+RvRs6lfVZM70x8LIuYj7CZkJZ13l7YJm4f
5SEYsaAFpoeJDak0YbfFiklxd27sR1szXoUhVsMb3hmaF+vx01LGZwuEB5Y6UD1vt1u6PQH2xkep
YiJ8fc6qgSPsZXa3qDn3gHqdcIr49c9AQldQ7bLdCX4rSD/PENXscMZ3shgt5CnLRFY3uUy28RFE
z2kC2xbaE/slNXJA45R+KLkx2met/7N9uVQ6nu6tN6cBdq3/mktupqxjT6M4AymHeJUdjf79ozMB
YJTePtCcBUWhOv0cgtob6B9VGSZJOkzRF4sH1z0qTKqiaJaRt/H4+Cxve/q8bZoHd9NrX/YhJeVe
YsZw6VW5OuhQNO1b1cp5nRw+vlDAp0QegiTUO38l3W2J4ScYloaBdHgGtQf1VIT8ytrN1Z7umXKt
eHb4a6ywzt9biQSVYsCnVUQE5wrdwajwlt4Nindtm+L553zYEL74rpHj/8zB4I8psh8pUlMfddyG
rRD0oQYeqD/V3fPQPCLLE/5+eHyybpF2kbuy3Fpl3aQO7QISKqEOyFrL5RybI/b/0AGZcRvnNsSu
Za0G5BbAO2+qQIrAqyb2Yn5DY1mSWeZaZ9KDYgVAVcAXNntbhSsElXQGxEmyCmvG1eG+gFQSPQeZ
CXINXg06KvBmPqGRNXlxSxBDKZQ8lm0aRBa0//ZbbdaktuX+02bWoY4rJiq8si76JayRcuSEHQU2
XcLZB1jpy14L73jcuNSt1XvSRKqAEDFf0Vd10U5sjB1c3qNW02vu89xf/m9eRLdEk+Xu1lBgbfpM
KdP4jPiL9pavQtiXEhT9eZVhzBoCuB7xESQrmuUhLTfHQm8nHrF8PppIol1yVY8MA0HDH1y88EeJ
ioRGlS9BYtcWrEe+AfJHLhSg17xgNtnM2DBG+YBzcYzs/6F20dazp340AsCL07ZKdgQjIsFMb1/z
sN5SMiAD43G+zVF6m5Fs/Oxh2SmDZXotXdrZX2D3p8C53o57XNfMY1dyskhnuaWyiAqRb8ZlZtBD
hVVCS3EutaFlysq/bZ8BUm7tRKfCqKEOgmzRXRr1KUcUtKLzck+5DyubJDKEJKRomH3+WLHNswiC
dF5T+CuZdyjc13kVglzpNDrkmGAXARJGpGo/RnqwK7M3s4/HCf94ITz8ZXQ3c70hncD2jDHnVWih
dLFhJjhOzpv+I4JWRACzGjQaHk7QXaxR3WgiuPVEAw7u/mMGom0DpqUSHO6faIGB4vFyJJnqovpE
3jU8isd+D+Zn1jkEmF3sYJBRRxh20tY7zNDC4Bo/ky4vqb9fm9T/MfsyP9aujJWXabAPDLmujjUL
e997Yi7+g8qxDzttRRB88oYzv79MF8F3kMMJYFM7kSC0xYuSZuO9Hxc/7xrsHoahriuCBYstctf4
irvV7pNfEGBKlIZ5ugsiRWsjLJ7f+rUNJJexHa+U8Z9XLCoZP7tDbiWcXI/ty6bFzaCnI5rZrIiq
VT8loBqtTEgZ50UzqgOXP2ay/lSqdg0Ilfs32XQAD/chDxqHtaS+P8ddd4dzQ0AM8rPmfkJ9DpNQ
JimdumGT4XJDPE+RfEF1fMJIyiemWLdDZN5WAYsygaBsfyGgxKRF5ZlC2sts41rsJ+bc8phmLZAf
2II1kA3vb/JEHi9MwVT7aR0guUR0QgfKOEf4evLOSsDVv0rWQ+lcb6YLeuOMkCCaKe5UrqrJ2X5P
gEZOLWW7dRGZc/6RkNsDAyviAqtXfPTJ+/Gy85idpctD3wU1X6IUOrpmAws1c0DJBtXaPaWevQmZ
MiPs7+A5dJXH5YptGIyy97BiC3fkOlY5R2/yEMklLbE+7Kj3hXtRyFQHLcEMfkmr3v39JBsc1Dcv
xwuBjlU+xbXyutVSpfAAbfBQgra6RO7pduvODkMCA7cy/t1pFPoxj2jdgwH3cfyIx5fut6UxAt5J
FzDmh7ErKK0M4jSMuM1GNr1YVgA5EieVKAo+uNuIDNdVmTxHIZdf2VT34E5u4bR8Wre4GJUpfZx3
AW2skiAy+AzfVTtEOcPPO9Hx+x9jWRIyICm5a4XTCv6zS1R9V4uBr4cUZADTAdGW+c+LUDmjURtX
NpG4TAb3mOd8WV1fn2gE848R63MNg64AcFMn7FLrWPJOKcE4QW2n1nLPimYgUBTvAZGLBsV+IyJD
d0ai96YMjplvM2UZnXE4MRgIYhV3qqwjyNJtzagrgzwCLs8dUbDJdK5EifWcxxagkBR/WPj+tXdY
0vyso11KUgIrlKOHu4Dt39N7c2mKQIN3qy5is1g3AvkK+e9MSlKmVxL/25DUq1GwwuD4Db9FdqPF
Ngn8ZTnIpjE0A5qsA6MERDdUyFiQNOQUBnpNpCoGHZKq9TxBJV6xBtzSsEodf6Zdde4JMTza/TYM
+RqJrZFVymI+0NVOr+u1oycDBljf/fwz2X3DvH0gwHOIu7wvQgLTU25U6P2FWuC/n4oqIojGjVdb
jXHXg7cd6HdwKqeDDfgh/FRK8CGJOHqAse+99QcbdueDKYdcWvT7DfEjwIXxZkllFrjpqZBb0MXc
r/ylf4kYwZrgiK9xoO3F9dzPMGbBt2z/j36jgs03jZvD9JdRKFWzgxB9/emfRJVr8WunufORUIjB
mFOWGujC4l4GaCGEvJqOzj+PMxFVYx2oNp7ArNvTQH2CrMGQesCoJA63DbSny2PRXQD3Tl4FqlYP
iwVbCNacttpONsisPK8vDP4DIIWXLOJxEUd1NW9p/aPSDBcnqKLsBzR3ZSmFg0VmKLpQ74l2fck5
I0umBbUFBMOeSG5BeBWu6+bP31FqYYplDGdTqEPTHmrNO2Mrjc2YmFhMvEuAkjzUF5DgN4KwSwcM
+q+0D8R/+pZAKtDafqFcY1wEcJuhxUfVc20OdZxW9HX7MM4hrqhnYvYM6bDO2l4ICOiGu3MaNXcJ
ZisbRGTeeFpGg02cwAZxheSyDecm6/lVjYIF6G4vbSeGyJ9KREV+4RVW/qp0Kj3VNFv/NDisyqmo
vCzh8BRzjtFHAZQQAEQylyImeGhFFfHXCpXFL9C1kVxTUSSBpkfNHD3K9GJZQ7OqBY4hqUJ7lnMd
pEZLrwqTii9C5y0Xi0Urohy6eLdm/DeQyvTjBRunucRu328PtXRPSlyyqoNMasDsE6StYyRYFFOF
/c1GZXIy3QgkaVBsVm8mJvlK1hPhHpIOSKpgJYX4yhtelm8lGrbZBlhSh/N1gDny1K5WZKnJ2cZO
isloJi7SKDZMZ7TTewbKsbyh1JD6wElG6qZ4RRlX/3zxFCH9DF38agv0C6t3sH47vnKsbzbV/C6a
B74dP4C6eliD8Q7xOyEwLqXoZv89Bwplqb26YO1q8uJHzf6CKSc3McyaPCY3l5FjT8kI2Y9sqig3
3ArZdTvUzr0yrdCmeezBzzbUl7chBR7zsO0qp4ORAzjfTiwVWLWJC2vFuZViySdKJ1MFqYf5c3Zr
pi9Ynxg+DBdK1TPAAEju3Z9POgeXuS8A8zOaFrhLsaNgfrDtptjJTHeT/FlL6CpoQqQ1zph0WWq8
Az+jUNrME0c/wrCOBbLRr9aZGzbpmYac2sKdIicHvRQzgv1MXf6lu1x3Uy54rMGyRzxtnEGslCeK
dWvZN4GCM7RvqjkiYyUhG9L0y4/7OSjO4S67i1dIYrwP+nu5caUNYLMMb++0C1MyAQKTNZ3pL/Fp
CaEPZ6h0EcuI+yBTC/592COKLHA7mtsEZ2If/Qld13V+5kVYDYXyopdHvvW5DbR5I7Mek3kcE4kN
p0gjQNsmiSjuu8DvTq8R7dx3g7EkmMwnuqgLrLKD3unM4vVhR09TIIGZnPHKLQULj2Cdi6NhPB2Z
XfJ/zmg0VRVIOD8D6c/Lnic31ojXQjxH95VbJ+s/8oqU94FoPeIT2plqdTIxXxuuZFAl64r3Uenv
M9l9f70NSOCYx17/Hn5JbM8ZWKMaY0MPIq5UD+qHQIAUJZWgaEqJ2+hfCwg1PlbhjtfWr4Z4ki/1
fVjF4WL5tJEKGIxugNdqjADxINmVVKF6pOVQeuO+LWSqPL8hBVZpMmexabe82LhEPIOyJpR2ZuNJ
aUBiA2UeKlJhNSYUJ9wPhgQJgX6Ft2rYgvXGxmT/LMcS20SacTeOiahyh/vmhwQvtTIhQLegFY8q
NDu6Yo7pp69M+BPJT4UgvgsHgcC2+jbZurpEfdTFJy/MFPlnKrYbaoFdftdDGpPsxyVZ0NVslCGR
NVKvhTuRL8mODmaD98YNt8XVQCMD3VClqzYgbRVAeJFMfh89FYdOPwXKGYpAG9kxQNgwlAPParjK
k8DyGzaz86qV63xcwDo4GTe/Xd0Hyx2vqZhxVCYhmuDwbP+H2NRXGGIpVmFv6JyqHmmW2zeOUgXq
lO51Z6+jCDm1rJ7a8mbR2jMqBnM/4ZXpZPqT8D2Bx5JQMrrz7erp+8i/jwdpsBWATainy74o4SdY
iGY5JDm5JCLIoDEtuzGJY5Rrzd0fYWRPLIt8uBcaDGm6EuwaGZPGlLD6wH0ltls8KROWMoA54ASC
MWDwJ7ZQwvq36J5R6UrGeqlQ6VRRBy50XVMUV0VGotODwno8Fo/Mt4km65Q3HSXQZIxdHxA7U6le
qyfPAjFW3c8w54zrNOkE4h6dCz4CrwAN1/UDZGHH3S0pK/wtzdgU08I3yRmhanKRZDnLwATAkeNc
6DvWF9aj9+FvGNxRdUC7YzMyfPIwSOnTBe1PWVshhWKuLjrIPBLJNP0l3uswqSOoEzrSXefshhEJ
DYvpHkcQuKwO5FAlSC0FzBq4EtsWp0szr3fb824+USRO30QH2ISRF66HYMYi/t7dQAdV+XtQP6yD
XJFW58XHamgNCaKQHj7oJ0eUUpraon7sG2unEZrmmCscck8bPRllzF7A7xDKH03tUhPM2xFtFNvZ
1kYVWMFzsBxCAWzW04NKXchKip078+cvAAzRj4ccAZtap0cDDDQWacBSDZKq5h0f4AZCeiGND9mR
WZhW6N/dqTTquenN/EoF3DmLESx+DcpVx5svjzlhRXQ55eP3jpNUGuL1fIE4s9n+ofu3hY1QDhDw
lWM9GmWu7DasXtOZCxlH0gNmXpH7uFa8sJmZJij9mFTXVM+VnmSWaKS0TK3LDlHfHXysiZgIVUTv
r4Aam5eshIBmjLRTyV1UMEY1vf7BFjRIT8XSBseYGm4Ea6TMkLg1c6+OtLW1dbTUZ42KW/srxTI/
zjQzR/0IzfN2Z7d6vkStoN9Ygn+k4MeL+TweZGg42cqw967vrm5OdKOE6LAmFRCrIISJanmYtWK1
BQ7uoYd7aBVQpNQQYkQQTVc9PL7rH8lb8U/kjzgXuuUmI4lqlLOLA+55/KWhKtAAiF1LB1YdC/Nj
lPrihdI0Apq/2dQoWSMX8jAkmO7qxg4AfyeR/I7F4YfSbr0pAjr255a9wVert5f4icxU687RwAGL
Rx+ydskA4Qn1yykjzHFhWmtpsg+LlqeE33h5eUokGpRzdWCv2KYVraBET+9sAa0U0O4cmmgMiNtF
Rcqqb6C8hUFPQyjnU4ATffxV6U0H6Wse4psKpgY0HJwhYpUjqZq10+VzpuruUdo50F2RWF1kv9CT
64yVZsJxsyyj7rY89c6Yo+MK2X+kOExgF4V5LfssHuAcFcY/tTMb6rB/XzI5eJuHRECx6UeXUqnm
N9PKyXUv3LBXHerMjHLqsECKKp+ZT/podrDIPc2sTu5aLdce+Tqan6ARsy+m6YvOUU/848PQUht8
mX3k+zvVo+dmIQ4NVRbA55kpJ7eskd3qZfbuyxpCT4HvFSD3pLzZ825sYaZI+MzUPK/XgI+wBvpJ
YRSxOzKu7qH6RM74rWBbFqrFwKo9zjV8r20FHMr1yEJlJvksGFo9+geC+38Ex0oyQX/c5BAz11yW
5kGG8dgMw9AdBTUp+qylDkphdJAQX5Hogkmap2qe5cMHlcJIDKjJv1YCvdsqi612YMwMJUuSG08i
WeCFyoFIl7bpdQFma3I/6QNFO1wrNnDrFzN3ZE5LQPmwXcukAPR+lYjx3kr64383zq2oi/7NeXQV
LgLuBsQVPGL3ot+deAWu4VWJmtmE5ZGHhjMpQ9F6339i3ta9XcEov0CINsgMT0T3jLI9yvj21E14
YLU7dUQ7UmlCMFBFDWPFPiXvtskSpGnJpJWOk0hJm4ojcVN1e0o/SsAz68KQVS7+LIvp2IZH3hF7
WdDug+doCx53E1ZXSetoP//Lbs0r82Q/Wv6ALV0B/KodUYowLmx7vOcFkOOMidencJy56JwsRa7X
er1f+uoYsXZKEzQCZ4t2IoAM3zqEUwgFb+w9BDn5yaQpqERSK16KneHYNrdv+/gesrL4CF0oJ6DV
ylimVM9zUR8cJArYnIf4u+Tc+6tLyleydN9nnw9LlAThgafr+l00UaIjBAlFRE84olaWWmdyaU5N
pDdSADwsumPtv6vUA9pXVTz1jyfszckXASBkVWCoyzfsRfvIm1IXTp/07qrX2n2ASBE2IHMR03k3
xj2w8IJFqnv400XTdl7Ka7s/+2GtfgsqV27fXk4R9Mm35E4r+ZKECID8H6L6XAnCt8HuToVTcaJI
pyPTbQVh/rlMR59U06HT/XKn2eojckk6Sod5W2U3bi6sJfERwOfZwkGxxcuK6j4pKfpbCyLk153g
90OlClPq1YzQZUkNz8FUtVyO+tstkWICX46XKAlVlJSlvf01X7dJOFbMDOwlVXvl3udr9q6xQts7
N61O+87qdSJ7rSA1Tv4xxKfQDpT062f3gLYAqLdEuPK9reTmJ261ow5OXC0eD/VTv08cAGQrVjBE
YY3yXNx579xINTkU58S1m4qy8j0lQTg9RhRzmpOCwj4XuumPWPRKOldbtDQRdajCxe5L0CARRV/d
jYOqk9U0wbkgHNoK3j4yy1J6HVXqTXta0xN6pu2Ph7UKHKxvUF84BXqNbcBYButVcUtAVZ8oPfgY
dzYg004BKY49CmyidiYOLKWejXMqlVu1zbgcvo5rBfitzfl7qgZM0rRyqwqgdDemEPtwN1NtiuJX
AjtAMWJ6ALX2ieQHSlLbySNBzVEd5IwSGMF5p/Vul6yjKlge/9SWyh26xRQ5mFHuzoE0fGRxtfZs
h9L+QO9dgCm7jlFwEHEy+76CS+KScJX0EnntY40TVOzTVYa+RLEkc2fbNHtExCv95FGEs4ZNl7pk
w8MZWPTTaAUeLuVFx9z2DcEQh3FT94tNz1mTcbxQIDbOgD1TmTJjOIV/lK1fZBo/LIEnBvtvG01W
KWkrLboinr0tuhBPYeCWrvlag30R72/Yt+l0ibYytBe9GUB61JE0t70X758BCKZ+YmOB/ORwvozf
tw+gvycPQeUl7M6hMrbCaYZ1W3YwoOoI+QQyfI/DISGwqTJB+Hm3FluOqSvJlnxNufVnpvrCqmQX
7s93hP3LG4PZe/vyssIJARqgtWaKPuLHUw48xbgDjeBjmvsY6Q3LNLDudJbIutN5kiXFWKMIrI/6
PDWfkHPZaehOUIWgyJoU/WZW4DNBrXqMqAbBfQ40duJTVUNJNGqHx03aoDX0NkEBKLpf6z7deU2C
8KES+L3N9WnHClqpxF+zKQJMzce+9skidcKCzAdYuxoFJpTzynkxeJtd7MLswVploUj5/Tse+s4b
ctHlFmGUU3XTC94Ivy0aSN14zFmPpPf/u2YPqdtIL9epevU70nvRBfZsWKT3bxcQH6C+zMX05rEb
XYu1/p75TuwZPLeHYIt3Wa0U+z863zUQVRq1n0AOMyVsV48wTgdCc80f0K8TTwdw7hOPQR6oChcx
1hcpfIzzCYlLFZMvHTy5fz33zocS5Y+T71JqVdjvgK9NTqvf3F+qikS0riKG7eFc2Mh/z0iZ/+Ka
XlrwkyfF/4UkqM4fBmbwxHsfWz0POLks6a7BtB2nEGSbItMJ7Xc0z/ceB/DRovw/GvlglJYawVuV
ECtriSuRGnXkV32SrC49z/5H/Wp8s/pG8Ck/XqXU3PEJsEvWt3xLAHuPKY4wAo2XEKQiJExctBXw
87Gl7HXH1mANbh1KyqaYmVMPoBJvx2haupnQxue5eUB8GROvXxwrv5MtXJ9Sm4DG/17akdVf802b
83u1wf0jV7WF4J/ivTcj2V7WVo0hwGk6STQiSvPM1iEWS+sx5FRWXsHqh98ZZyGG1kPS24l2d6i9
Sd99jUvmVhLZHDhT2E/5sWW0XUnqqHWdjtZ3Y/9FLMw/5Iu9aycixf55kghTvEqFHsYp3gnbrvS8
R23t2/58/IDYwV2FkE/6JysJuPgn3P2unUniyc3oL1EArEGkTBaRT7E5yK6b5F4vKE6nyhogMnud
i32vdGKDNnv/c5kOwHjVXPt3CXmWrhqu4DTMZ4HezLPskqraa+8wyF820FUej4p18thSHAhqLrGv
i844azIZIe4gM6K9zuN8+y1PBNcVpz2PN6HNeDZQ6RCrWTAVMzVA2pTyQcStkXTrK48aBzMAXFqW
y6aZ0+prfr+4g5zLIL+aWALSVBAbclCyg0dw9U/h2qO7BpkJEqpffgEYaXB3PEIuLPQMp3PIX/Ti
3dNR1SmOmvd5NLTrUYGjlGVobTnFolrJ2wMmwBUr6+Ls4VDZ5qOLGrehuy1tercffcf6/8Rhlb0X
OhV6g++BwCnJ88ekuremky1bi6/Y3TRgvUUIy/Z5AwVHOBFra7tvXEHa/Dy6pWBMU+j9JgsIr9iv
uxbYS3JTtoVPk+MjKiS+JInl9DCuzhe8RwuNJhYTtOQ127p1cLpeo3XzzyyQ7iV+rOd5cyYpJi8I
Jkh+Yz+9UR2ehLbvvgCph/Opw3RrjyRyE/2WZeBCFDnPKAQn4TeTOVSyaBvvochZ/manTBoOY8Ms
VoDKGNcloZCTiHshnby5tvPMDRMYQuSEZ6cw1rZHP0VRgzfrTcGYxZX0pfWf5+Z2szLeQZfDZDOn
2Le+o+jE6jdUNu60Ap1Mv3v0WDxZDghAhiGZMUYtPBIqQhuv7qB4MEvIcaSp8xPktqJqQqeN6etf
Ofu9KOCLWa/g7BXYELR+XYJXY47NsxgkDP5LDgNnCTBRIzAHO+DiFC3zcj602wBOShANyVClmU8q
W7MT8lBA2aSEkPjchn04ovpGZABt58dqRGcIViJ9GuT7wB2H7QSRHklkVqbUd7JLgQwiauQwZ/8e
+bDR8zNb/GaJlgOMdkka8rE7J6ZvbUiFwYkVLFPVNgxFnyMpgEQlAutJKBn/aoDeQgaayKZXDxs7
3yoYoChJYzpj1G9OaWCKf9QkeFEay4qJ1kHg0Gw3yF9wiSrNGpNfn/SLkNb9mCRMBYDciD1Xkwgb
wDeHYxmBV4CvkTchm8cAqLXjo5tIgUr28iB7M38NVH4YDEczANFkw1I/K503g9oha01vttGjqtwO
aUwy7j1dmgo0tJM1Xs74ubbz2t1e4j0S0WP+Qmr/E64pIM+84EgeMxxfBZptW8M9Pi4Y7Z0AbWoj
FKveAwEqVFdfkbvSuud8z6PKiwPRFhgPcechwp6J/Lh5AraZJfSQbQDAy27ziW6XzpUYNHLoEjhY
JV4CINobH8KZ1cjvnLdnjTY65Oxf4KfWkbjj8DiZkqE5zaSnoByicxWry2rEj2/ApUMRHGiNhyAq
aSHKwvWrkV9I25nmL3Pl6ZEfOJWhU1fkmoSvXU0Mx3QUNhWzixYtYGQxJGF4SMI6QlWf4rQDFPXL
RACwzEPNeglAzFfIBUpbN80EfUF2/0G4Jb9NSBZWEJGQZcrO79xr3xrfVS+HebSdUXO2RQVnjdCT
pDKT2MQSuosb1MmdlUBzn+tYYDr/sVUYIQSuDZx0e+qzSnxeSAIqLJfQLL1A70oq3U5krkbrsalO
L9m4UlwzsJU3L63j1YJ6jrovonNA0wa10vHpJscGf5BaMzpnCSJnXT/vm1c3J12aY5huIqvv5BLn
7ynyGH3iM1gx6aTha/PmdUAYenS4ksO49C8sXdM9gdjlJD8qEyIXFaLM+jiLEilCUYtt4X8N+3n0
KVtoVWWaWZbf+TG9jIx26W1R7LzaErRqnDWOr/q4SiDf4lC51wmvSYbcnWF0smX7FkPpFDW8w54Y
BbEQwCepCwZWE3vdQUq+VHXXhQDur2Ag3rdN1vO5459oeRbSkjPKzLOB0NVShIFpRWlIiyw2TtGS
d23PYM3jqzIxv6isCaC0BMotbr+bI4opCWgSLNI+azj/E1YTYyGwSAmG5gh4k0S0nl4+7XRHT3yd
3qZnDG5j5bXe++Xme2TRbNyDf0TWppFEuyj7VIQDK+HBNqUO2PSQ0OFq5TPgvUEfV0AF8BzmkcHr
mfUIXgEBaYYSQt34I9ZwyLmPmTp2/xMuGpx+G4vyu7owxbqK2eK5Y+CEsuXJDWXLPfTNNg3QfMfq
ge8HiWN95WqwxSdD1EVNlpxNkQ+GF1jVr/2GnZL49Zmz8B6qkxFJqg7na1D9nUtHN93wt+URzj4S
Pqg/YfWYysPOtuKcz/GSG1rqZEWvlqkSARBruURm3oX2TkwkluDSPaHu+PChsAioBkIyM6imFG4+
xRcuNlqWe+JLScHwDolkzeMiTzcNULhD5bb+FgLBFwFK4ky5t9B9W+ZNBuBy43vpW5c3LxTfkX0t
W26vjMUWKYgCeQgABBfNjvlzHCFg1aCsc3dbgxuNF9ovjlHmZYCz1K4UFutjkLHBKDsByiFqpqLi
FiD0vuOLxPIqlNkm8P4i3hP6DnIYH1PjA0d9SrwXurUljI1EAs8UZRUv5pNa1i51fDmtb+HAI7cU
naTbXI2wPbjfbCM3nYQOWeuGgz0078pHuTKsW/Y8imIg+GzacA0YbYfm8bWFzckP5lS74yUQuTEd
RyAVU7y53PCVfLRE0xMeyY1IYBAh2UnlZuwMhkjS6YxM3Q7qvqxdywxVHEifzbYa0qGVHIsMibd/
ZWQ+A8G8C9SB/8T1vzDQC7a06vfz8udOnlz7cXRWa6xLU8vGcuiNZ+98kPdmmN6suiCITzgt33Bj
9vLPmniLnFe7SCUGsgcL2+EyC06NU+RE2j0bQfOT3TPHmPDvDiePoX1spgIV61g4dVA+hKF0lzSn
TOiEMpfm9S5emONNM7dp2SlnqXMEFAnm/5x/VU4XaKklADDrR0IsJt6JtFWQNQ8hXXojWES1aYuJ
lzwyAjci0j/HnamZO4W2y2obqeag8OkUKtEEvWWkyI8FDq0l6IW+TesOoGRIeNdJ+sj/YiWQjeG7
z/WF+Lo+f7h9xe6WwKtuk0f6TzZYgXogNiV5ayyIux2ypIQBCe1YBmw7NmqDgVjULEtXv7UxzaNw
4LqLCw4F9eJladdN5KEtAgyMVwcVLoOUenoYMNlA+L83oBb0NY4BVdm3KzSSc6szEA98Gkoangyg
Yf4wPFfXI30IeKEaYbmAQc8HizZyH3h1GtmGOGqABQiakOQ+m+dVi6oi8FSUqVVQA5+lKkH7oZjy
Or1lgWB6o4PYDNTsa41dVUt194jM2JemBMYw1bqZEUnuFw4PsUcnWH6vX5hpe4fMF5rbJ151aTb7
l7F7sMOdnWelOsZWZdfMLxbIY0fqI9oO1q8rQko9bQqC1JRbksNAAHx5Zi9w4pMZWd8QYi5AM9Oe
uulvurDX8jl5klFv8HhrhXD6Rwka6A2upUIY6SLLXBgFMfqtiWNvLTw6siuxRP1GkIkFHsUQYzww
SalAoO31gWyUewkxmTK3+9HiIkbF9EmLT+0uAkHnRXCfuMeOFcmDzBNMUaNrVGSDgtuv/pcrATVZ
2SJ6mz7GZCnykx5kItLlx4F8TAiCupJgnRc6ZFuGHU37FiE3iIfJ6vJDKBo3FZFEPTPuLGxPRIsl
jqgXxpHCm/Z/KN++bIc8KwWALp8N+3Rcoz4VFFvmPSmo5CpDTZg/LAhC+KjN3qwQldGGY2G8fYZQ
WU+X00IwxYAb/vhKUVe+ZlYigieZspGXlx/PfYAtHWK0YJ2c/HPKUkYquou3q+Py0fYXuMsDg2KE
oZMHJYvDN+lW3dpFQFAfD+pV6+iH9qC2mFcsMuFloz7+kt6T/is6XvlqrmGV7co8sacXVcW+/aZ7
GMSfCEboyfZyoVWYUeAzmwp8nB7oP1zvLDbjj1GM8yRLIfX6x1KYwruv2JnMeyEIlm6TOu6UKAKn
qOxJix1Xu+MlbQW24Dn9PGM+99/sOYCq2U6VMuXFLFPVR8I9SDycoc0naKj5pGDf1vaP+ReZokz7
J7LP95wL6PBVIzxE6avhpEtuXyV7eWw7jS6XvvdBLqgXvCUYpxnu/wJIoMmLVexuxbj1nrpl9opb
mCcBa038+Psu8qXLwmrR1glkP2azdhXzsmE+1MZNf8r3QFKNjplztsfUiaOEyyPxi4Q3H+EMarGZ
q5Is+nthOrafTYj1Bupeb8MyxEFrN9+JNJnWA1PL1rT+KrbpS4uom+bgCAyXvgkdUbXjsO5z9zsF
CACQD/RKzv6famr1VdwcdHaTvz09r7bciDhZNGC0kdxrNL8CGV0dNZckkDs9aPrkfGxICBQL7JSj
GAsms1btOUQT8/nD7epI0R8YJ+8j4+I3UOvFlPT9bPB+sM/W6G2KjyXwkKXNTTj6hC5RLhZtvzeV
uWyDHVGlKOMgsfhfRayEnrfGMhftaCEeceCK7QuAqLWYq41eQkmhc9h2ZbvtUkB3G8dIOYhd/Z2F
Fzhc0isfU5MPy0qAdft4vT9NosFnx6kvypFt6f0X6jLrK/G0Hz/l+qe7dE6NjwmZraXKQ7vu6sw4
0c1I6K4C837YEXWKoV72xcfWCBujNKxR038qcqynUBG5eKJgyOBAJSkzkf8hctqmYH9GLXDfpk6c
Z88Ot1nBtUYNBMFCkKcmd5/G6xzrZmXrfmxOCU5Tz4UsTUG1PmpKv7BDdQPf8H4gJVkUkPvgQNkk
EG8GsQLg+0VNhvfOu6V+NoYymz0OGKurWtv7eyJJkjbiOroTiZmGn8r4w7dvQlBmJj1f3xa+OUkk
O+CimdBF0MxxORmaqOqlwU4SYrPdjoRRxsMCC+FKFDCXX5YFzXL4Ystw1hL28rlEcYHXajbj1L9y
w6V43c+ag4pycUSfqXg2fjVIaHswoYXGcpxfRADz6T4U2Sd9XcDZ92pZLHzffOjF+6BTJoEzogxk
NABtqgYGpQyKuj5DbMmbx6hdCXlME9WNxf209SDIjUP7zCVYD7SwMqQH4n3kYKtGF1qJALV5x/gy
jQY8VEYvMIJCVQlnctByIYAoZz2alerp6KfKEiZhgAKPMoenPqdlGOMBF+f50/XD3DP6+rCPPzz+
k/B6PIFz8QyeaA93xKirzMz0EfY8cBdc+iAyp4io93Sw5vKZMnm/dG9kAVbd/CCBsybwcYXLm5NC
kwv5Cv6t5uMzT2vQxjh+2pq3LAoQ2vkl9BRVMKKoj1VJNDUZL53sYiRCHq1q+ghfzxDi4KbaYUQv
qr4CYG0IdpLXSJtsHtZRK5jTpVqcorDi0MQKU6t0gdu7wolXrh7S5e/24DHT7Qr146io1YhP+jXr
1Re10vw7sKmnJ+uOUjMoqiAsjguXjzxuJyCR0GEmk04ydA6d7dnRyWZ1yXaweSQfGvpaeqCqooYe
XIv6XCjogleVNiuowzDXgxtMrHWgnVPZd80AELLs25IsZ7rFSbGXuK7eUMxJMUH8gZajnSkpU2Om
GngdymGAliojuhQtLjejUHFG6SuzQSvkCgPzZH2MdqDiyrdWQ/a4+94W+CURogKB5fEH0pWj1tht
eKP9P8za140kp9H/DDu9oCQRij3HH41S6SnQoX5k8ljRG3VUe5n2wMGq1mfdqtb0gA3oybuef2Mw
hTkP6wrC2y0M9+KHy/aUHydPD1mOKasRAgPX9TIL/RG8huucHa97E7JlFe79Pw0dEe2Okxh635x6
4hgNpHywW/lmFNivYIqMPJ6zsszo3bxYHU2Q/old98rW0P673fAe+OCq17Q7Vws/tdGf+4t15veM
GZJ9LNY8XNUf+tj49F01b9JHtcippPERt50lOqg//vjPstZQhoUNU4hZXSvksEZVYCLozm6mdH3v
JZI8SU8VHxxkATh7ZkQ+/3AqH96d5FtD/r1Q4JR2wzYoXGXU6p25XBgU03yZXb47xazThGUxjVvx
fa0pKMZyU25V6JFte9Sq8849+Iyv6b5BFGIZ3vOMkqmGDPZUg2fdwNKxJAeRFwfivHZ8Gf8Qvzol
9K0xphhrv7Wvy9tn00WTh9LbFWQxSnTJe6P4nlQMztKva/EU2n8kfJJlCTD2hmKkZMl/s5nJs4Zs
DLY/vsngeTqUuOzcTciN6ivsPKthB07GhBo5xvIsiG3/YJhpN7TN/8jzj+fWlgQQIvp0YBiDNoND
eaNge1e0mDYOrfhC3fPDGR+ZvincQVTGnP7VNzJLfAezuzzbf2YPvbOxkqQ24rbtDfC08/xyqyYD
+Bi/w8d/n6MMjzTnv1cwcwbrTHGlxtkUcvYug8mjV+Bfw1e4SieA4jduFHS8UDLZ5nGy15+10EHg
L6fWsZg47yMP4wJGfnEHpQ7F/Ac4QnwaoC4DzPJPlIiz8yS+NkaLKx3ENYpjwo/b0W02JI62nEfz
q8z7zxapvH9o9LDr9XkYSLYEJzezq5yhVr0vZRRZMqgFwdZbxd6FGs34oHuWbelSjjCMc3aEDxKq
PF0VZLjlUHjxYZABt+hl8XSAy6d0EXuDqFZKNWdjbXlbinJwFRAZ535cDFatm0q+r2t7vcQm3QY/
rk/8bMKj/rMkNHwsDimpDbvAQnovF1h0udnYhlATmAgeiy8NJ9nre4BH9osi995VQB59cI9eW3Ms
t1JEjF5s7vYI0qC6fuYV1D8Nkwgzc8f072Fa2k2gJFIWzo0mB3gQroT/1mqzj5v1ixo8QxHyucqK
op+QQHcmzhXPib6mc5peLQIXp2UxMaDReeDN/4DXUk40M1DovcOFPs0vIbrwLlS5PZx9Euta+4RA
yUaCho5xdN/MfRTug2PyRX5meWaDhHk0vvV+AZJeFB+8pFLqVgFKpqeui0UuBLxaWUIEpggSQWeY
nfa2Vuil6fkRgW/geinAyA2l9WnkkOW5a9PHK4cB8m+du0l486gp78nn5oYG7BmCBq2/zmTwOyu9
V7jKBjbehYQvavclzH3lMlPKoN/1/IlGR8wPzAXNzg4VOGVpqGlG1hYIoXpiM5DsCKgQE//c+4OC
cCQWuKS+znBtztlmOvDQQGuY3W6mwL5+KTrVs7wpcTIGj79qOzebK2m/61YrOaMEMlKnX2ymGKcy
tMp5svCMvVUOrMzALEDRWTlzCfWCgSeuqryGfOJqKxpxYNENvKJb4dTcgZnJIe08ez7QLrBzPkxY
k6xGqUOEnmWkFaNvpBuB3Ktwv7VvtFp5t7Z1kWjzQfcpTmyABdHJgq1Cwo6Ad4VF6uSTmtXSr08s
JSi7mUAKTkgbRD8RGH3XmYrhRyHtiLBpYN9gHorNjNuuwnuTCCigwK+N8Fx7MX9iwuJ6Lg+8XGFI
7uvaBQ8xhL8ryFzw+CvHpAE7ONHH/wWy4LOg2XAacv0Vz84Dvpje7vKycO3Wg0XudKajRgNtju6U
2MwylNjaSXZgUywvehgYhoM+7b0Nw1DxXOB/S7rIPgYlKaOC0eciW1qF+/AxrsxAWYAGran5nra4
1V1Wla9xFaqmrOOWzfOog5RtJM98GmZVXx0izd75hyxKyuvK92IP9tziLy5O3ZNBC0AdAfwhKrTX
BKx157bZ226lNmeFllfaWUpWyeVahVmdJdOflFwqwxxAlK91yQNZVwh/OOnNMo0crcDwt1N1o22P
3jnQL7Zj5Mh2CvxV99J5CJMpBRY9y8KynZ4dlCgYaGPTX1pjGMtmTkpu8I3Qk3eLZbmmlWCVMk2Z
BFTwBllWs/EF6HEHHvhVJvjBFa2NcardbDUfweM2j6JCAELLUGt/RkqYe3+so/5+4h2Nu0Lwm8QO
ZzuCLuD2cCS0PxiCFSjau9cyEX1bqF1d1QHps5galacHHHYZVqxCQa+gDJ7IfTBCn3r+EmTevM4F
Rv3mBuA2fxBFG9Gnh+B6Qwk/aXjNFEmRDW786G7M6mOIrFm4goDTplvds66Ewg2xYsGxE4NUG68H
TcE234vCu+tk7DlaEgWAiL0BcOU01zCKrQUY8PVwjs1+ysG5Gba4lDLk/0CaUTOtqTUnDxeLVTB+
p1d9+DmWLuZUxK8WWQu62KI0Hc+D9wD3ZYwCEK2EJ0KPG9oYzZuf4TmZEogiPdnqzQvaNilR1sFv
718zH98E5wTe1sVKgpWNQi+nCF5RaAuuyuxSH3VMjQAypvDhiZn1e3/vsMEfekITP51WpfNRlzVb
r8lP0mxLs7EhuPq/B6QySsoGQbRD283+Ptmu2c3uJG1n5BR8BVvYm6Pxa9Qh7i4nMF9JXIVHz477
ySFHIlWfiyK5hrl8q66zLpRmFk9rjDoRDB3mOzcO2kxOyUV2x/1nr9NEd34ziX8hbf5lKFxw60jo
Gpbz5y2o7F6ToWhxb+RAoKdJ3RNw0d2LVnmzjzg4dx19Lbqj1PENld7U3UldUVcB1QmHkABBxwNr
1PQcfMDWXGw2ZRU6Sezvs763JqaOwXn+K5C5DdK1IHdtYvxuYxuA900wHOMPPzzlevsPALPXZSmX
RmgIjG5sshvJ7tcIuyG+FJqmkuUoEVVlnng/UfY2hY6SnxRFhNH0Db5zjgM0s5jyCidBpkh0e/ab
E8OjT2p/+AOH0RocuNHTUmBQ7uKP7dJ68wC7U03VUjV/P8lJPPmImVY73M6ARS9ImXd1pG/6keBY
Me+PmYxg1yxDQv1uQlxcUDDz8rnkoKUz0QpAZm+yfjqZicJpjnh1Odwt9rSQrO9dlwi6akxo5Rdg
T/EV3s02wusR7L8WEnFbjMtuEjLXUSY+bDum0Fec7Rj5nTV+fa4d1PTAA8bo5WzGvbi6s3XbhEEY
jQUga3+l180+mXIQV/vVySEJrexCv6bxwzFW/RUOe6YIQTTGBU0XMm01cRf/lcqRbvtYl7TQ0oFx
rcluCOV2xZX2mtBom/ZuHernjW11qxhqAQ4MIqpEZMbj7s83NtaaZRVHPfxg7VkmSrEZ9/jmR+1s
TXF32X4qi+7WEOL8UPGHF7ESNhEwTPTq/R9gdUMHaZ/q/2d2KAr9YHtLZYxrLHFoFM3qUoUMtC58
Jr6eE5xwF/ThYqzk5zlUe/u8AcIuu/7SX1J/+AFITAZq10Vgw1l9UT6tto6MV+YFXVYiG+0c6Hwd
xkMnAPw2Ppdh/xuyMjwLnuaVeFhC0hlyQ7XjFg/pBx9/nLc7Blxrfbun1HsabDiBD4G4GXehZxPN
pwvUyhwp0QI9HtrRRTm4HRi9ZuJ53hFRiYPhjuBJABAsbfOkumHLdHdHLkJwKlBtsfGItprg+Ms8
uMkzyDVAAA/pAAI5AU3ZQySSBq/nflWqqO5cfNN+NJPbMq3fybHhrf7Z5Qvfz49PAlLcDLQoOhPk
EBRuEFHK7Xf0G1mkXyYaSgrcB3WQ6vndFgLBOqeJZta5TlzGcLoTDv1HTXqSOmtgrPLwycGggf9q
BybvypRRx6glTPMzH7C9OpTQidvzTcFTgwbovkw7M9EbRn+ZJ/wKelnSSKBOwkPgUVcG+V5uckbI
Hv+/gNYezMkAH/HJP6cm/BC4rR1IbUZt1hoFLp+SBMRi3pZMgu2Ev8yGv1i4RulA5kwzOz9qHMjf
wlt/LYTJAe/994EJBPoMm01N7Ria6X6czQ3GhQwPV2Jq3/eH++8zdguI2Jdflt16FYYqpZjZOYgp
dgdEO6e+dmgAJudlVH4uGNPA2ZyN7/4Bb4JuKA+bHZU1HkVf85FPl1fjhEInD7gqPKLdUSsk3XEG
sgO/Qn54CgMap72PHlX2w0wtS6hfSvVO7ofKX6XxzsBErtegArHmf0IVUn0C6ms0IiEzI4KO5w5p
W4j+SXn/1O0lw9HaffvkONhr6SSVKY/7i2TWouVqmv0SivIbTX7BJnl2U+7SiGGNtdTpICo53CJr
owkXU1ADTZj1CCqWS1l59n9SSM6G7i0G00erthL+rnaooSGzrlEjE4l2NYFkENYkQ7Rrm6er+DLM
vqdNrBV+aKHuuOtTOuz5KK5aCrcLuokwm0edypoG6VnUO3S8W5Y7yMBp0hMROHzkcLMKU2vx5x/f
ND32ZI2z1jzlquJbfpgj9kri8OqFJXjgxOfRSdibbGoJ4HBq17n5DEodPouMQqUJGrfuHzXDXH1V
UYFsz5AGUFnuh1T85IE3745fphuAQ/KGaZiGZutEhU/HCiyr6QuQkZ//Q0VZVmnIkht1CkkZrpLm
W9vz+57rRkoeBV4Hd2ywoLKQe85kIs1UuZg1XtRQQqWMhftFBeD3ezhkRb8smRq8TZVNE7+aRuVu
Vf+3d5LbQctXRLD/wXlXMbeBopsVW7xwBR7LoFwfqAkn5SfcIoskFeK1PvEY80PtMzykzUmQSD8b
AEw/IW0gG7SwBXxEF8e+jny2QT7h2yKo/VP3O8e+7my/T3MffxYJgAAsfcMkhRv7HAnFJs1aTR+M
Zdeh8GSxI9hB/KFuE8Ww+9aear0zsCkUoNt2wZlTFbRym1dMsomWVZR4c/fHaO9m4Q/FDk1SpArq
xYqcaex08TEB7iOQwcJisOugkg+rKvIMwnj67ClTXE+V2r9sMSKyGHCNIXjq9v2/2uY+OW7rspqh
4I2tsFZiPFRzU8iECDMqG5yiOrcw5TUrK7BPtmXhJfhXBrl5J57LsnbtQCeYo7jbQZI8eMMwxrgr
JBrqrO0kdj7+Fn4yv911hJ0H4fNbOlnPxSCv/7E2fk/J5lh5eA0DZj8TkVjjBC4OBsqA6xPgCCr1
bWIMZ4WUTg9XJqvpSzlBBojqB3rT7vVouzz3Ml3vTBYlbXKuIhO33LuG1DBlBVbMAKhtnWsTgKQx
sA5KU5rVGDk7gneVLdBbaqY9cTna7S1D8eUdcxko/VrE4BwodTfEEdaqdWKNrEiW59cz49dhKsfb
x9O/Qn5KaF2r1iiIct9NXyErDI2dRJ1qImsfhhKZrGCQrmtp95T2LEugG4DDW8f+8Huh8eHk+NQY
YzXopVvLOxl71ucqLoUlrLo5NPoXOWrjT1XMtDJlGgB4U8nhBTsyumtbhzyqJvhGg0njFMjBJz6z
qrYUgZL33iPk4K8GukYTaqoEBkzaf/46C3NWJ0W9SKsFWtz0iapHOfYUD029HkMF6ARzQPZQJYBW
b87OczA9GrQS/HUps0va+SEElvx9LZryWhwQXGoVse5Q/Fo+HlxAmCO0WXjKUp2tXH8dhm77JJzV
t0l1QIpyy5FGH2pCVokkXUx6u2aq6MwZUf+xyQq5xfU/nclryi+T58P6tWM/AwTDwOPRRI5VakgF
LPTtNWM16EivxSmG5mNS/mlh2dJZyOlJSMMKPpKUobuuImc3BITgTrCuouqLmSJrkZYTuRC9FOWM
WLv7Von/lOOtuKQbUg6L1Cf1K9eshE18yB3OzqwsBOkY7zAUaokP+9Rs7lBXZZESkO19BZLwvBnT
axUbpv9/km/czMA02+h3Ru5pqSx6Wk5XZKJMaetfVn1TSSwIwce5DSym1pLSmSjCbGKE/VuOUryF
FVmwPRL8l2CKWwYdGW8pSEYvXN9O18voo8TJLVWkkElkE0UUhY4wwumesrr5djQrxNFlgSIM/hva
5QB57LWUipV9CXUvR+FWSStyb9+7EJWq+QnEER9gkTAcW93aF04gbSzFLxX0CsGJZpowh5BY+fpq
bEfnoK2Bxb9RTeOq2ddJmZR4R5IWclYf1X/liSbZZM3LNsSLZ7D+fAsCw0xtdA9gaJ/yiIWBm+Hi
kfnf0fQBuouEKolr6Nswg7N3N36ysCLr5Fq+zuXS5hdqMO5vUATvwPu03AI7CTFWIh4/99HCU61a
UC5yag8cTrG/gT/TOIQDQL3T6RGjQm6A/4V+72gAKpNvOw92PwbZlN3+x51r8DQDFCsE39v5PXeS
9NSskZDCyAt+ry2K2ipEIZZj0VPowYDdhTnwlR+vxn1qGw04SXKlyOdtUET1LcBIdfgL9l0AF5gH
YaMtAklK/IsBf833zqo08muEmWc8YY5A0SeH2WuKddYi+1TQdl8I1Xanuf83au4HVyz6jtE6n2UI
c9SAj98YcrFxjctjKsZhqkMUZugagHy6b1HmaeGLHml4nZhRyFQHhGSWRVCqsU30MKe4BvCv6Qtx
iyceLkMo9Z1tOMIYO8szq+OVoy6V3m9XNNvDfgYiWOAv/zMIVICUmJnk07cY6PfZqWyVrmaMi3Zi
ehOxaCuU4cAEuIOsq7rAqJEYEgK115Cdf5iRZnV3i9TV+FNgn7NWtWl904T0XkEa2HNur+wMIS6J
eONxtYdqMENRa27uVVA5uElNGSceqwJ+cmNc0hXnlFHm5/U1DyS3zRxY+S3nS+r+vvMXgD1klC4w
oB4PRdEGMKcaK4qwwwSD4b7cWT/+LG5k/1kUd/vyG9kCxwpPdOz2W5b3Ak3oyT/1soiduOQ9VhLg
xH6RWwJ1ZbJz9wDL0eF5FvIaA+IwDe7Cnzl/2o6peUNo50+v/PbWiWk38qeaozpuBccjYNyBaDsC
YygtEvQQeaHQvszcc8v1qD2jdTZL370PGbh3U7cwgqz0C8Xof3zM78eXyDMPvz1Ih2VU1BxSy0fT
PKG7ef6soeLubslZhRo5MWBKI+sKTdnrA1kYmelo3MTcYj2Nx31l6+Iue+c2fGKtUS6d1sT69QpJ
cw0Smef8WbY6AuCIznTWJMh46sxce95Utx+sOqlFrBiHL9vJdl2EnkvWSruxJBEwfiUc87+Lv7Am
O16VGMiaCJk9nGzgsfyMhdiy1Q9Yi0rBalAlMFA7k8vwXdBGIlmfGZAvPKom7EE9s9NzDoS6Eovl
ziFP5k82hlHcr4E693wpG/464XxRNDrgBIfMXwRU+evL23mVMhl9r7pRt59mMIISdFs8lmR+VQcH
Yy/s45WmkIg58HLEyVSq39GQ0z1ntiI+lMQexXNmbFOKWhfzUapOohmyzF6ErcVlLEaJb17i1Onl
N+nky7LFBO8vWC+nvKPefCNjaijvxVxgAcT1zhYUy6cIzcqThoBKQRzRkFnpWC1Uh0i3ndEtjkrA
1n43WjwGWU7piitz8GbSb5UDPB4hdJBMXqTOVGByWqHaVkqkqDqOzsOhvi2qK2GQ6Nytj6HcUOan
qISqu96dp9l5GO8RmlzEwA7c7xeI5BGeHVKoAsY85/hBw7SIqJmjI1X9gJYgXRB+ZC30/SxGvMoc
z37CVFihHi5G/amqtlJgLG6VMU54QflDwzy9E+CrwfdGvpmFYFFGp8KkE9iycWeTOLbGbLeEoU0u
O+SjEQkTh9yRuax8VnA2t5XYo0Wtn9ahWCNP98clgK5tXsaU8ZnyAL3hIcpVVbZk2BM4QBY7J9TQ
8ZUDP8ro+MEEC2/I/doGKpJHRVKe9zf2F6Dq3JilRkr5TLG76rmh6ItZY6sxxXC3a5I58NeWPf+c
DLcuJsZQaEW04TjsTS9zwIdrNZoOsB5Mgh29R808rxJMMjkMF0usx/bRNoy2tCUMeK8AJfq1GpL0
D+BQtB4+O8TaLWMAxsKBltHXMDld7JfP+A83t0PGdP/GBjk1dDc12AqVRZVNHVhg+2L9WDVj/mSt
LkpPyqY5sZmYQhq68auDhMfyP5dIoZ/z1Bp6L7wgBPAoQxUJ+1Tll2yRREY8MK6sGN23t3JkmjDH
FI5Kd9R20hjvoGbiCxTcaKIMRQZtrE4wxavgBYeTlDaKmdy+otbcPHpB4BMTqTHnDGhaUPJaGsOD
2pvka5kYyQYSmFPDdi9Ac2iEFMcttNi7k7gsTE2DvlRVEbyGasQusI08rJtTtORsETb7MIwvQ1j0
jzrdaIqxrhJyG7wBKOA3pqEFoHlnqnwYT4LJcIWIGxS/vtEJtyS11KQLp7L1gXmvTwxFA3xPgOqP
bTsqozQL+5diCSzEBxukzqdlXCEWJpmURbT7DEqJC+lN/r4rvSElPpcNKNca1pxMzhT2hfldVI+a
llvcxa1YCuDd7GUWxa9DJGp6RdGwXykKJgyLdAuwfWUE1AtCIeEpbI/UE3fi447Nm/5zzjYyxVJR
8orD3uqT+22donHt89m6v1UpAetfPvOk4qiVB1LCKBYuKgVTPmwL6bSe4c5spmYchKZBbX09Bcxp
kl8c5frJaPHKrSJWtV+6SXYq6j4Gmtf6tF9TrdMRzXbW7z92K8cG6ikr3jumsIGO38d1gU9R42P3
nKT4kFAnpmVnn3XOlTWzb2YCnf45k76sp2LmDy1SETp9J5hjhSoC6ImgDZtoH7Erw9eGMYbDtYZK
+jWrMFkYj6ZH764hp+SXRxO/U+I0NtWlx0IPIcQcqBTEfXhjTWmgOKeUwTpJjyifcIeaG5QanJYW
K3F9UauKpos8fPKQuSv42frrDhqPBrgiyhA6y7IVXJZSGoJyGM/lo90wlM03IPlT038KzwObKhfO
uqJbNxJUif10mXsd6mg80CcEFXunnWNf33gm8CcMU6I2noN5pScAzcpxNjOtsjAkTKpCDQrH11Ar
+we10HjcGJG3DDCs7k3BNdGiNbbQlw0muOpXjPVKGPRl5uL/un317jWO9w7858OcDIMqY/7d0ZlU
sNlJBCk17DyET6tTeVpuDlYnoMCqIEjo5H+hQMImtUm4J2ByEeSVW41/D3IffsRMgqYRGYi5ljYH
NkJjpvlwaIABqryAgYPB8DMJgO6zzmTtPxkTbskJ7KmfbUqDEnIBDxj+d3h0E+UEes/HSs3x1zQZ
gUTf8wsyvxiNQFUQS5Fw91il8b5N3s6AJUsqTdI7EwDIgaCYHea0WW/Wni/i855bmlF4ZuV7zIwP
WmAA/jM+H5MXO58skvpefc+lkVDRPBqcykfZFuy3FHDzjlQ4sdvPbVTkbgzRw4fGTLrKe52ErRsu
klH2FRjKgaoIcSIE7YulhRGhmp1XxBvJXgRkgvgkiSro2b/bqL+DSrM830fodQxlR+XU9CTg/iy2
Ao+2dy4H208MFXmZ9rz8jHtjWfxBXb5/P9JVN5/I/bQTwgKaWD83HKihozIS3Y2jYQKuRQIa1gSZ
S27rTcZneqSkEYWW7BZ168OSfNcJjjuo+neFr3LAH2D+HNLIStiyF9KsnR6oYeXD3oD19ARvW3pu
FFs29Uz65eC/A0vvfjh6RLAvFB0UVTPzKREMJBePz4B8tZAyhzkL91pCX8OldE59DttUclOhRg4E
vAP/ZUSVnZW8j6ccfhG65xdZpBn+NqN29HxjqqZbdCKp/2EljxxLz7iuNcEbwuKnQ1COFVi+sb3z
dnU0aj33u/qOaoTrbQ3gkE3CKASoW1XIjKc7FVA8elQe3AjdygxBjWTbfdm40jGTlqHsFJgga41R
VXRrz73kkEyKu2higkDYG2Op/BG+/QadDwgCnZ6tQ517d87hdvG6IKK1EgdcM7P7bwacEDSXwTjA
ad7Gj154YXEZjHdquDmDJW1ecQPwt3arZQzIG8/KwFHlvd6r45vnkz9YhW4Y5vhgCOZR650+t9da
gKXNp+KppDx8ulTNY/os+rWQU0/0DLaIiOfzwIg6HvyJdsY8JlciQwO291+SD0nBuHHZ8FKTZKUB
S+gJi69P4566qqHyrIBU5k8U6epqXOUKNZ6rx9hIWYeUn8C6yQJc7OKwfKy3uZXSKkA2QCy3UfYq
asXoPkN6OMhpeYMKbk8VYgAW3Gi4bCOIZRQTKKA29IgSobjqb/OILDQwLQV5srMb1cUecCZRG0Y5
IHsifbkKHOUdA4D8L5c1KhXR7NEF3G5NA47vzOx8NRm2jvq2nFR33388wChpa5yD8j1atW3uOxiL
CZfxW5fQO/odQ05f49Oc9uFU1e+t9P8NJ8bcz29cuqNdNPEWoI/xg1o3zudBptpZ+Z2IIkcUTbC8
wTZeLs1s0T3/WRek19JX9TSMyDn9xuVlyFWwVvfJU7YBCC3CoFWn9sW4irDuZJsT7tkEiOCX0mYq
JuHwV2ZGyGJG/sj5V0gYIJ0Ffi/T0CU5xy0MQR9YuwunCnC+S7a6HM4CBCaGfrkr4fBSRznrTrN6
HTEOabnH1seIi2e+DAe1854E0wZmUA/GPlbw9OyIl02Mz8Fcf8ecwbQoV4Fr4IwSYMh9osWFlzIy
ZK+dC1550su4itp+YVcybNK4bXpXWGkQ6AN+kc0wMD/ilzCM1+5yMTOwOr1jXLXJ0752nMAUmreg
PGrbS/tyzjUkLuCvRyJFXcToSY32Q1jj74/0a8ekNol+ozBrSsLYqL28DEhnhM1VQc6b2ii7+awN
EU+UyJx+05AfDWqjjK0y/gfATehI/tXiD5uaKYVrmJIxGQ2qCEoNW2IlS/X84YDh1F4vDEWAroTK
PGlhy70IG0yfG3M5ep6vD7zHr0dUAAzjen+u8OSVwWw7fXmIG1ri1Hf1kMiR3AerI72ybBSEuFTD
1XxN/YfF+Lb7/q8lbntwlwlolA9wdqp/VFOjH7VdU2UCuJLslHc+FVaO6EwZTRhnxZZxweHIDbCU
xRe4V6mezQ/x5YellvjNsH4SJIvXxPAtteZsd/zMih3UnRanJVCZSF/kZccI7OaMXwSqbUCtKkup
emx+jrGDucep6JMVZZjifpYweLm+WnNUU0OO5qWpeVLaYmpYaN+8pioEvoaIxZZu2i6Pkb3O9Vsp
jfStG35XaeciBvNWO9Otz1lLqBO9j720uH/S5+1eao/lQjQr3bamrg7D20cNgX/3WxF64gzs242J
i06V46pIkvHsRwWE9cHh9rgNLP5kELhax0gjbYNJVkGKjXKiO3AYEgj3/HKn9O+HEZytdT5zPSNl
k4Z4SCXUsDr/NoA1qIjqxczakmPbvjaDdttY1t7YT6/BEjhlSKXwI7SUxo+u9YEsQVa/cYTUJifw
AKpBMSjcoTdu7JC5RAsAG+J2i/Ql8AfD2EgMteImzbnAhn3hw0wcaAFi1WaTDq6edAoTgg5X889w
71GS8+cKdv7p3jggI7yGmETE139BhryY4/JmqI+Mu3bw9bEZkcSK991GZE1r/KScCNE4kvqNYBeA
2+0QFlV2Lgn3uApwAsshfN3LoV8mvFaafMIqXpFKTVAW5+M2nD2BkZrQEsQqfX1cQANnFwGp9Mti
ha3/Pcsm/x/d9+UEajPn4EDFZxQwx6pFBAw6CaSoi92Edloz7JElTD8l0HVoCJ0Ctx7CkzdRVypD
2K5hIiPgbYnBwbdH5PL0bW4N3Qp85Jz0ShBZVWPzpdqXN8+Eb2Oprf+drmvSJrKWAAtVUqCGjg8H
tEfvzktf+acbaCdIVfbXM5frdcqOw6uKitqmB63KZXutpHyeQqE+fFkU/uVD5qaqfp0Ty/US8KGp
mV+7Oy0N/n09EOCFSgHDAqp3Z8622Le8yze07SjkpDJDppuhKmDFqX2k/Sn2Aa0vhp/z3+8j0ZME
M8iDApgxRTxeyQ5vcl67pa+laJ8JefLg2m1HGiuZrzB6HlTA/IsJjw1a/onjXIgFZU5u8K92rV2s
mAIEiTfzltvqV9FbCEYOHwiQ0DcxI9IXJs6P8ARj/OXQytlu/g5QTEqL3J8hcnlZBCen6ijUkpip
WixJyv4kEUzf1gubnEiTr9/egrrEbPH/MONcx8P7gIYZKVy0LcmLUxNjEf6xHFvTurJvwzrJTNBA
IE/RLR2G+yO90UtgWS0eccDQffetCCNBTclWXDZvbit6PQblV+NXg6YA3h1968tZHFodY9675CeC
HoqCJO85RMK3zuk9AZi1jNJv2l0/P+jTlcd+KA+N4xH6+Zl8moIk8ufaCWLtsn121NhA5GviE2ow
X8tdBouvrsM12GZ+yweIkOdjQw4l6gStNx1Xf+PdSHTJG06dJZvavoc+sRdBRDfCTcH7BGfD2VgI
O33AVcjpNgT7OVU7jvOobERytMZHKTVEyrl6SwcNjSi2ItxIMStMceJSyJqx049L+7hP/1/8hN/6
kmEeRmddcP8NAqS89grNAgkhWdPGozhwrnDpg/U63i4yVefj+X/Nub15CJjj6jaC1VpBU1OAsmoK
bGqnEOj0LT9wTZlDBJgrCXjmtHv/cbgqr2X76/e6BKf0FhmHiB3DnSwjeDM//0U20xNkHyLy9TuS
HDyv+DlVkAx2EVF8Lk4maTYQh/WsLuf7a3iatJWk7gEi9oPGtwwAQvcPtJtpl/GmxHcdhjmV79U5
vjyPV3DSZWw2UpP/7CYBI8v6ay0nNyV35lLbh8oIMA4mNL/5gT8y+UJJ3y+5nSm+UvCCyofkGqZj
v9kYsoiMqyablegmGzGy3aPJINg7PNFVgx+ft2ZsJfk+UvK4xbyKTaR+3FIORe9kD+9+NLmyp7wg
S/bbcnsdTE3Bs3FbnB5lC8fmzGZ8MOtBa95AI4PfcRRS8hLoH4i+5DHtmFNt2s1GJhGbLGHun2LF
P1q4lvuVa6XT01rvdLG4O95r3OWVs9OXY0cc1CEIssrehW7Ho+UJUUYHUBslJ0SR5Qy3TzmcajBE
IeolB0XfUw23SJj8KFkO0OYrCEImKotZp+Gyxk1Ex5oFiTccjeix8AtSRAFg4kaETHBudpLjmfj4
3Xyu898dM/3YCeHqCnecFWN3F85idN6KKDvWNdsmH/NkcdJMMx5KP8ir5OTMyZ+iBqQoP4OKR592
ceUbp+g9KY/MWgr7U3MacIraQ2AE4qcRJkhOPYi8ZoDj8BpuME8VelZgDhdixlAqsBWEwXx7LQXs
tzBxqvi2kRK0fW6A97Y7c4mQTNNBSZWXoY9BfMWvhXwOkaaRKNOe+bodJPCaAK4FotSewnpSxLMY
MX3a5+3oU0OxjV+QUEgnrOYtqfT7xkcAROgguoPu/7Di452e+yoHnWbMuiO5GGIOw9D4/fAC3OGQ
5O8QYtKR2jRRTE9kPk03aIlZprz2frB33/kbVr2SJM/tljmVlsUdZSxGboDIknzHpLmsVImAhBWq
8Gkik3FE+Mqhb13NR74sHh2r6874uicUiTpFFLiJc+8Xqc5lSASDMtGaA0ooce4t/ym83OcXC3nC
kXl2aKx5FHX9Ctww3nWcUEHeObehSrcbr6apZFai+Nzx1ln9FNjD5a75xZB84NfKqdppJfgk/428
mHRS7ZaiFBRIQXmqlF6mre9MWjlhCruyG4Hx/CFDmN+hbjKKKWGtbyBp8fM7SWGLJCPrkhNvS1Sh
4WSkEIRLmbu4VChBLJuLIaoLTfcfwi5pq8QBRUEp8x1P/PQs1ZHUvEsJD+senrOrwLJh3nOC1vkH
FPAwk1Q9ge4CtCPhX1QToKX1i4y1u8eI8m0o8YtUNmGFj2Wa6Nsx2FWK0IvuMtvMA1ZNWYbhh1Hr
/OwbVYIXgr+xmEI+rwYFltF2+D//Mm6IVSe3tF07JFBX5jlH7JjlAW49o4NIvvY6sa70elcgNW59
Eko7D8ETjERmiL+vL4SZUDdUuA3lNyQNZRJbiSqxxIntQXmbNSh8BE63JMRw0YYNpIk990cqCz2P
2YvnPe0CR1W/usoiG4zDzzX52m41vEdQMLj2bhisSxWX93xE2pCPFAZ/WZKF1Y4H3Os3WiaU03zE
dG3tuW+VwI3SYTHnOgoM2OOkJIUwDEM3+/ogE82g7VPoVXlkC7XbTBRflVlTv8Ik2v2d2rfKTrWG
4aNujNo9QS5hZ6OT9WPOgbcgHJuN1IthRfcCYI4JMkKrof4hfX2K7kcgYG5IHIyIs8w1gVLLsMNv
ytmLdBSxx5GdLKo3obLlOA3p81k6DZ8hpvWJ/vF9QssW8Bh2GjaVkwb1B5/fELCmSwXLBJYaMhbf
OmVcX/1uGbPxbwO62l/BJ+7TR+pdwq65hxwXz6rRc/atRnKyOSxV5MF1G/KUQsxELKkSqHnkcIOA
02cUHR37WwJYko6ZuYukxCnlUT0oqqeq9HCzN/ieQpQrM5K4cduCVYIc9vMLwq0NvfIAbYg7tEfn
6kx2uNqHYWWNTcvT8BeEQAJ4Ja8JkGTBtn65RPYT7y5Z0BfAUC21Dz5bgSe9Eil7FAoigFvvjprr
pZfuZwbPKK7ILMxXJW81S1vk4wMOM32RmqVQsR0CMd8Ng93VmlY+XxEomzubUrya+uaSnuxGYD6l
N3vcPsiqOPJOFwO+DtDRGrwBwx5xNQK8FrpHw3a8dJ1PJJdiagSuUKbs11dm/thv1bC6cOnPZcmi
24vEiatMN6w9ce7jwPGbBBma2vQs/GofhMb5AQ3/TNHsEd5XW5uowyNFnXpHSOSt0PMODhpbAsqs
5CFokpmRWvLaSzX5yrQXGudwVEGrVBXTtxaZ8Y8/nNqmhHytu6bUI3Zu22d6cHhFQ4NLrXvjCrKE
EO197AkLgYw/Od1bkilElT8DVp8xbQGYhnctCjebjzSESxfpl/tq23m3CHe6Q1cpKOOohP2sMayr
bDiPua1bs06o0mSd9aVFPXSE+GCml86gQ0Zv770xk3+OKH9DtVRcvkwbaJCDEfP7HFJBmvYtOSyV
bZ08+Q3gbZIk3v3tF5M0gWYzgsYFAPKJkMcGwq9OyX2tT99qYzKStDmcs1FFPjM9bhNqf64+OIrL
UzsS8g/TRSV+Jo0z4IgWj0H0vCjYsGkyYvYiYzzROwfkS3KbPw4xYv2eaw43dcaFPH8BAF0WRJyM
qZQrzDWKMO9Tj+0k2CmljIEtVX/SDonk5VIevQMLWMFQjQH9R1jY4THMPdJxmTbyblL+6sUeIZp2
pPaE0c4ZTz1a0PXRDIJNNV+VkkPJiRZqVHI4Ihv5EMEDJSxi0f+Gpeu9EWpAgZQGMfp8FnMT2/k4
d/hKkfBYAaqBbWq610HJcmHB3A+9LI9x7XdnZw9pFTIOcDj10vsd8nnPwpkGnZJd6Gz0FNEqkzQy
Ur9RE/jztl146LvsVce1ZWnnQA161ZcW4cFRgWfZSwRBkEHHUtFemWbyFWiwqPN2g4wYHQZ8PVWJ
XGoDuiYTz1KubdUH0PLvcFnDgG4IUveB0QtbJztOXQxwMjoq9PgInQKkxLIvmrv32RXU2ENpFOjF
u/Ma4zSmVc3SnICLNB3Y9/8IssLNJqk8gEbp3TpEc+41McocGWfd63locaIK1wOjDvOR8dtrMUPr
kK89bjwYl+UYzGcU5Sj2gKRzOh5bnpXLCmXz7ZLt6flsCd7bfeL5hPipnl3p39kV3oMz3ubOW89R
96r4hLK0JIBB5qOVvOiseZJxRkCDhMkHKq4Bou6A0ee1RkuiYTG4jw+CWvmRKlC/NlIhcrCHqTSK
eXHSbBFUW3/abm8gARfbnBj7f+KTUVHw7Kcke9dJbd5/sROOfE9+l6Q+AjDglkXcVOUXB/JKfvQb
N5ddP2ml0UiLLK0sMM3Ao/02ak0qgy119UWO7Ds1WzIQ3lEIUE0C5U9BJH+bgNu/GFjZU2OPg6YU
iaaebGu/QvyVkJ2gh//228Pd+AAqGN8GA6k+J4h4crCZn+NMEMn/NmPLXrzpS4VvOykK0e4cFh1w
EIivKolBco88vzNdjSeQzw7qSiMNiYjuKLv8L7hBIzM0v2+uDC7QrKg4aczBdVhU7XLO1mhWj904
YKpGTb/4uanIYPE6JP46t26VpVUol6fW/BSIh9TTzQiVaHLjUXStrZgOpfRbVZpuuqBGQrAtosNf
2a2Np+eCXVDur7Q5C+eD0ZJfYgSMFMmtDiHp9VCG0qENfLEqbtWMnx+n07/ZTy5hAkNmI/k1bs9b
qMX8vWfwraajDTQJKrd2Tza9rr3ImzZ5yYkpWesAiPEPCuJLHNEylssqsra/sWLJHUuR3gYT6CaH
lR+mJQrIQ3az5BcPvnGfna+OHRsomq9g+RjOt49TyQMZlXkl4ViUrtElb9ae45toJeoi1x7nHIE1
UKRyXXAkw8AP7GTqZvK6jg4/jT2O6l2HQPEbLb2XFblJTsmubJOrXMjia4oz65UNaS8wahThY+Cn
EofUjOP3hvrHvrHFlQPFrDPG07j0+38twLKHKQwSQoILe5yQgC7we0uXyyUK7nmY++hRXa7hOBs5
rQ9gaYAdWZ+CbodLWuAsmJe4Cu3qBtGRq0Rt7hvmDLKzl0poZmELBXaPV8IhR+9Qfv1AYygWwuAC
Ni5A4KLGJR1pZ+RKqf/F8JqZmjlYGbGYHhunqo69gV4uxgvk7QENs4KeXGX6aUNS3AvNRC7NNMpo
GQNK0sXDC2HTcEHhN+sYNn0gQyxsTyJM8kb7pes6o3JoqCLalHSI44LfB7+AUSwxxj/PRRPGPCjG
AM5S75iiGjnzBTCEERCnBmMIWDgKCX/bx9Yz1jRdFKm3tcF/97b8fNsDFayMrQucu1O7J51xd0JH
9e0bRvlz3+9dLGJQbBLk41rdGueDfIRUezn9yclzUq4KrVgExMOgdArWrr6xDyNSqaxA8UfyEK/c
+pPTL69UxsPYBR3kwLvDUh0GhvoCuVACt74BgFCnPgQPbq88jKqQMN9j9WKLIh/zbyI6tcfBg4Ss
y0oR3cSC2jsPyEGZZy63vcro/vWPwzVsAm6SykwNt4HYKuy0UUGTRPeRtezCrToH0tQF1MdGFV8G
aC8VKo3Llqzf1c0+GNFNu6VH1CY/vVFVsM0jyKRupKxyvpKOIyZGAaQki6+Cu/leADM0AbFql11r
Lpmx3OqcmuQ6omjsUb5B/6P6DxfksyOR9Ir9VlNkq1D6N9EZy+t0L7koIaKdIH4R+I0MHlA8kEvr
CuiboWAiJa3illfjYhUVDZymxZ0Dryeo20WD560jSRtyf+dsPBTtynifSG6Ixd5yv3kSqbjWotH5
qVLA0hjPqT0CDT98pGNqKmkhIBRd9BuDcPK3Kcr5dx5AfFIBPhNEfunJRM6uTZVieBGbZRvOGkpd
fwqlZQF9y4SkywDnDpm1vrapN/ZVVcyCdLE8I/kl/u7OSFt7mLPemaIMm5F2uNlIDZGzUz1bgciq
LK3YCneLwJS07lLEwkO1fPQhO1HpQ2vosAACjq3MO1oIMrEB3XR8uqa0fbL1VSCIVTR7G14HukVJ
yH9z0ujDIORc+wPFigaMTGXq9+YNFWaNM1FNcm4srZJavpS2xB1aXNg+4/HgylbfzXMi9PkYXC79
KAeY3DjCH5dIYX92NmVaXueLmAWS9NeM/fPBuNQNVtc+7ZK/ukv/RM4VNJgWze4B3JArWtyR+VJn
pcD+/PEBVDSc0cJ2NgVwxKp19x22cPVRwlQzVk289n/vaA5wpjqctnGrZyZZd/JQL27GDHI4h8KQ
uzNoMeEGdEvsHm3CMFCN/g+uFtCYxTFMYrMXO6YPr+SmqYlL7up7seOIwthfBPoB8IW1pCqRyBt6
tj9K568Ymov9qKVa5Qyxd/+Pqul8OKvYkvWr8ullXYffkqK64+PuPjYamSn9iZBsGehF7j1fPx2/
9XTN9YZk47+EYpWxBZ6jTYWMUnkj4stZn381Y9ZPBk94l1FNO6rW8ERUSIJNMqu562Mx4n5cDgGG
u2OSAQVD71sSJOyTkW2bE6PPlp5sF4f142aN+LCo50Cedc22Qg4D4GGiI2/dFfEVeMreTyGtOF3t
hPOIG0tsxN3SAgQgQB+3ODBebs6hfwzuwij//wiyLFE3bTVWihuB7lRxrAI2NXJDGVFfyxv4gMsr
pf73LCylA0yMRoGOh9LdSO+dqUj0FmPLYnQYpEKzr0FWUXK1enfk9EIht+0ObKNniX1PBLESBsgC
grrrQwahxwnRAFOO+1koSWh+zZqSIidHPghpP+XGjQWw44lFvt0pL6q6EXzY0Y0vkZ+L79rBeO5v
oKS9tZehPK6a4mCMbI5n7BuyR3zdRKnoOPCKi9AQdhTUKzwUEuQ+PinuhgefmBCkg/c8uJB2/+26
Q0WwcP4PBsve1wZT9qp324KPcz4jxRCnrvv2tMbUNVzh3thW1fRzjtD7sSNgBoPFZ4ymaoMHeuzM
Ua9drqZTmiwwWXis3JNvTktjzv7Q0tMDE05oxyrJNGGX7HEFJ7bKm8KZWCBXCJJZbxh9Nfzd2/jk
/5+pk9j/4mQBVduZp5YQWeNFe7p3RM61R8djf3D5B8BmKtrns8glzw8BQgwXJCFAi36sV8kVUeRS
ehNGC5iW4EBnQAAkxLa/gMq3psrJgjFu4houTENr7hobOIIrrrHjW/GVD089dsmJ3Z0njkdUdKtf
xCe1v2TU/N1LwMUuSKecyshGSnq54/7TJVOQtOlhjWw0Gb7NkS9BbEb2Sx0gqfZrGeGFbPsL9ClX
Vd6S9FrCLhnxCGmDfb3t0XppitaAh23vktSFgHyIFdS5E+gRphrHGzGn7bpZB7wZHJQWWqbf0JuC
BrDyLP4RwSuzkh5G5BaeH15fkyfOPsJv/F0w1rAuf5hGlxm3zx1f75XJtWRPD/xCRr2vGQCC6K9q
zyNsvs784lAZVPsSNLIVjWWsAnRyJrb6ivzFv8CqhV4kvGm9mitjSvFrSliaY1/G93byP8sAbFUi
uqyjnfualyL2mtfiUy7AAwAdZivV/cNPk0NVfE9yskDmbZDZKXAk3Y5AleWfEJDKP8XYiMkTYZUn
oO4hb9HkJlF7IoijSE+woC40tK1pphoShjDX5Ngf9/VorPNrXNgwLhH0VIS03MsXqSQNxOc+gGsq
mmxrSZEPwySHCkV6x1k7himIvUAZ78njf4xSjFPwe/O6s+akMZRPJt3l8q86+N3yaY7ESVjjhiUb
4m9fCEamfLSFjJQ+OEj+xymSHUjZF8qANVJtE6n4DpMr+NNHI/BUtAJwZ2SisqRyRuLNZqFdxlqN
qfTPHlroSTq4+WDKOJ3YEqJgit3So92umsCGEpxyxOLjN7K1wVHlv6pVOL3sSD3aZjpC5+eXGdoo
RuWE9qMwbI3UQJZLK8FDbI6EJgqDXwkn9QyUAT1HQP6heCxLU9UyqDOufBPYKP3KENOH/GFBBwS9
ZoS7/1c36AEyVjDXdL/ZIkd0B4Wv9z/GJ2oDkD8JhEy6wc/jJS6x9P6TMZQS72I3onYknTGknBTI
76rTZLyhgh4zg7/a9kx2b2aHvCbhOYcPTTdBEPANYhjv1vr6sB1JrdZkHmM4aRn/xrMnnTaxQ0lv
GLC+U3apD1mEyt908NEgMEozgW88KEyYLksrlKZQZjd0Qg5XwbXAz8e/SVYmoBW8emxeZWhzYY0f
8r2IefEo86hqCpse9TI+X1jDUB4Pct5WuQg5ifudgMoFQXT3BGa1hrAm7cHmPzMm+FEBeB5yDpfu
bZOAr+MK5buSzjy+DiZbcs2MFjKlR4q+Czfe2KQ157G9FFgZSYzoRcQaehEHTBzHkIddHrY9jISY
VJn6p/K3BNg4b8dumQvdEMMSpnIsAFjmYt8VNNYKBIm7dMQpactZaVmNLWtMU63q2DVVBWomiJPI
Vi5kUfRXUvB9oEyiwZR3w5PDmgBfOgBV13CXjLCb2ZUfRwQwJBbMmv8vyhwISYigFNyUKneeIEkS
D/VxtCB4VloNej9VY1ITJPc/YWZ5dqfw96cCbRCmcW5kPvNiUW6FsBzh//hBpk9B6sDS0WUoQc6l
SBDDSB2P2eKTqcqmfwP5CXouTRJ9t8Bu33lLDyXOzT+NaceI8EmfciZrMovJlX/tRA5XhM80tSuf
ElL4Z+76dN6wTwMhsvyQg7Vr+QUyKNPdo67gzO4UgUilM68Ig5pFR+67lgrZnMLhxcuMLSNmZaGX
vqWeo45o9yu3/0KunlI/PA2b7QBw8jrjgrm8ytfOJLLCng5omTd8IyHoh7AOvbw+Rqz7a4YitTDQ
mnM0BLCwjOWP/4fhEohBzj+MKBp3XbrT3Mzv+S3K0j7R065fzXOdNn8uKP44CIqehgyOKRHUUS7d
Iy3ewIzFn3aAzXzUkJSRNsmhzBh2iVjJrUeAhB2pMYWI+u5Q3egM+hUIgZxhDLU7KLNZRPN5G/CJ
2folWWB2I5b3RGvsRsyl+QpfHg655KJQz+lUirgFrSjyKSFRrmtEZwt04fjCNirtrehk+jrPqk6F
v3n/Nm3i7NwKJiRT0+o95BN4Zfl6RuOuYfJLM76MX9uFk1MW/16+kPgy0MMnuYggnX2YVJ4mn7WC
3ELH+g7+d/W5c08iVjmJNcsaRUHhPf4Eumt6j4a+14sd1XGIeIkVhQaWEq/XU7xTJPjKBW46xwI3
HrGAQ9mgZfF+7Cy91Odd26geIkV24ItFjG94xc85pq8nNFX7mLSgiSQq11uI4Ur2CO7+Zlr/vS7T
BHd37ONQMEK2UCROvaMj3N9g1jarNpp7EzwocB78l99NP9XWZcvJ0rqJgUVFFgjNNjlY/aeyTbLZ
xRPNgx6kpJLiLq2CgFNzQh7Ap7Ww24/0KIBDdxElECyZ7SaUysA8hajRuUzqoNgthgHt0xvT08TT
G2rjsb29AigkNf4cV6gyou7a+6249X59QzNlp5HUcJfNv8LDCkhGRruJH5aWOIjpIVvTELrz2znI
O165AqQqyw74hXZxZeMtlkS/zJMTm01TRf1KRe1aJItMIBJPOYdWnkXfCiTgWWsdHGXANh5xzMds
tYIWjwJdLGjVpa7nrtlvv7oqDcdL1AyVHrsO4IuSuBEPMXPMpb2KXblNrtoeSnEVvxVlowWH6HNX
y40PpvcrAwwVB6PLKeVKRJbDPICSWc0oHg2m85QVqLvYGfPaAtWuCv7IAKLHAb9WD+cd/hLB5HVw
6cQ7GhCxDptsBWnLuSZzZif76v2gBG+huXKWpGAuXDWaS5qxLT4oPwALaUK5Xl+nxtPHJERW9FQz
75UmxB/Wjt7GEeijhe5+0zOzlwXyYo2ttxIyoAl7ewbeLurgP5YXh7VuVxISOssunnG3DJEOBZHf
UWLg4sHYzSBaVQIDQxlYy7Yp2zzdKZDmENZ7qByKR7Kk62uMpNWCBV87F8Nz4T/6FbvBW6M6/RMe
ZPQO0b/GEhqS7JqHM6liaIqCfDt0Dnvq4FgtwmjvtB5OjJ1DVhJKfpoTk/wSXJ870Cz+Zu+ybr4E
Pe+C4UrUVYYwPCDpbi8Y0KeIgj5HtmAdNfGHCstqYYDZygoaV6sjXinqiIIElliL+tcRqwB2+X+m
nT2hjWB1ow7fXOjFnD652y1CcK18h9+/WEW+pbrHsE0KwBo+WpM2AXyIafD8YyOXcIiZ+QxTyQY5
p83O0NkAQv+DcRrVLxfEshme4z3irqygZ85enW5U8cEeZpZ91u1VAY/52B6Sgcb0mj0h7aFMsOos
wTrQaSZPdJi5YYPiWjZ1faakzJG219/QaIo55KESUKume+wLJa/2DJ0ui0GB9iOcT8s3yQSM8mf1
P3k3SiDn7tm2elsQnw5IkaUiPsPEtGqr3b0X1c8G6uxMmUeTbcfSkOpSXnnymdqjYNqg6ECOjfEB
/bCmkqowjEMTmE/6ROp3R3KO0gPgfxEVGwMWoG7ZlcDVYEA7xbGdBLAx4FQlux1dqjwCmnNJw3OR
w1zlYNUj69i2KwclPUy99Dk0ideQl4Yt8rxtxaybF9YL21f7qNY+wn0TN0vYe8k+BdFYkHdsfvFL
4HqMmY/cL8K0frplSauwdTxoLfHn7sOZK7cuupvrhDzwPtLTrb8kslwBgcUsxc8jpooy4wWIXqxk
KBVO44hT7Rx6oNOr/fH0Ww7La8Qa6VV9HR+83AczhQ4KsKsd/QsvsCiiQqtV8Gb6BdfLpS4/nbLK
qcBRTi0KxnZE4Y+YU+dI76SWbNOLsRgBJQLrd5lL9RjWq2I/XNYTUFG5mFBc57glNIVos8c/X3pH
1o00Cs5S7ZCXDw9468d2uwONAbXrdmD87f3Z1JhJuRGaSCzU+eVxsx8FI71TvEQ4IcaP/g8qF7JK
H5KnJqZYui4eHmJFKQdAR+re8KLR6XCH+Cwijlf7FwEN3dHmEpwgazN6O5U4LKwR+o+OjDbHyUf3
jyng50scSS5b38ba0ftONOzRb6j3N42AvSnmpDPIRJpNFomfbkAFAjleaqwm57P0qK9XvJBgqw4W
gDTMAvnqwpVflBLXeOo7BGzrZSDrq5VBDuLGN1ke/G0qckiEqYbd48mwaYxgcZWmQvbVclPkw/0y
GiYFblYmbpHmXiPKAvGDQ4IJLfP/uLPcZ37YSZl5i8DEdy9D/4Qk9avwQZYOBf4y+EycRk3zdS14
EyWXha0DuGLn9FPp5/M6SfP6nqlJvxCRBgmsneU1t/miJ8nO61E9DA6OuOIifVCvalADnEkbrOC8
bQYG6cmyHzl5pDRVqVsgyfEqzWGgVEHjHZxqctPv638+9KpR4T89Lz3sa8VsFzddS/MWn0eJ6CD/
QTCg8Smt/XIoaSmv1/R00p4R28MHA3lYXbzHDlZKJEj8lYhLDa5mXQOhNDn+I6rCaaYPaHcQN1lW
yT9XLW3lQyJzFR01EiAoyvbqePH7ASJvn8NyTA9BCg2uLfNI2BYCuZ5txFUoiSsMY0HAFIiz+ZOA
Af8LuMeetAzJEUCU3aTH9VNKj1snp5m09YzEpwVtP0sJKKkVS5nww7N0TjMmDQH0ioG+LT6cDrG9
bOhTg1BaU/oCXwUTyr/+cCsLbO0+6WOumqn4YCelnOgCv3l5g2POYrSf4RaEKyoC32yLF+r0tBsl
J3rs1KHvkMAsGqGPdYLSNZ6wqFKr5hZSyZxcTGNM3+u8b1ZpdnA5p8q5DbeQqR7iRFnrdR3TxQB5
cug/lTj4b7QozngG2/zVPIqBddIGhzlDO0msopg1c7cW0n6CO87FoRYi2tQpF88jJ+uVWcSuZoaJ
BwXNOlRSeB3Dk4b55IfAPQRCleSkq9bQkS/S8xSygF0GsjrbSY+/82JQyqnzqHhgFJCaWaY8bY06
nK1AcERyeg4eXrzYpaBhzM2lzFLIVkauU/OJnpWZSmv1X9bQQiGA2JaHvptY/uGg1eDfQfy6UDeX
1VG8EIk+ZWRNHy8R5mM5DQ8Sq7Z625CZPCEkU30bqJ7evaLdGGNi3O0eQTfERifWOrjMxSPXclL2
MJQKfXFaEjPMqPs0NsCjcrWpd1MprvwIayIf1Wgpibk/o2mXgcFafxsVGkwLRO7wvgQ8syoLhbTg
4J3YQZ6zML+i55nUuwTGgDyZQMg0ZTJAE2K4cdZKlYuVCSRt8UniAdGig/hD/AvCeWWO9HFbXdsO
KRgB+oNMCbINQNkHgoipxO/LRP7PehHVrgJ9gFRHUGamCamvUt+32YoabJPZgpGlqV6beJRWdhYP
9ZKYAUoeQlX6ZWEKHAfXCDnJkESlfiuTOzNNBpsguPFrSIihLVYYdB+OrRaS5zOwnbflXBiGuQIO
UU/1c3UuCKMDTCgpEYmmL/fPoLX+hYICku1pqa4kY10vuRo8b9b8ojRUHrgD0Ym3UimC7G88ZXNV
9LThliXr8hGpkWXVD4+lKdk+1WmbYkpyJ08KZ71eExLUBx2EiioSGxePDAaTaEHfBTpGTmrf7yH8
GLeMAvOi1IfZAdqW2IcEi/ODcYEzTFE/BLItQw1tjZawuwMTMM5rSn/CWeYi71ZUYWBefcOBYIuN
+FxLD01KotUWZwmHKppWr/Ng4PI55v4haXRwgF9grHYTTbYAcppHb1/YsmsRLcL68ZlYpsxScFEK
noph21d1RmrmDh0ucILTmI6h5o4/b3MzUKEd43oy5nRhIxCRPmwRhb/4LaeJ/LExrolYJalDIWjv
OET3NbbDYweZWDbNDPIO76e9yQeemCE7DHnwTqJmX9Vj1bN52gewDYqZShFal1O9rGPw9H9DxzJD
6jfDKevk+/zq7A8xgOLrrBqV9SBwz91fcV93eSL8xa2Syfcd0/qJekmvaiFdGInM0dUsdcamWhnv
ieD99jzp+L3CUXK7FqmFphEx8ghEpRsV/C0JUcTqi6X/7SUlGAn56y+qhnKx5oSHUq2PFCkuoqWZ
eSEiKjB767ujnE9kilZGpUqRzigHVVZx+r+EAko8APtijKoEPwPPCSyHJS4ZJ37YTN+HM8o250pu
uhx6sagN+eDB6YzXIpA6Bx2oYbzLxwoJI/0oWFr4aNHnL54gKzZG8pWxYdPlxdANVkFzYa27QT00
CwE8jjJVcNKS3058Jn2mnKauyJlsvuUqpc/hbN0+mrjuzflZgU6N9MuRj252JfsHUej0hz53+hvs
UuCdAJ7xzAvutHNl9a9HNRfNMA/+yDPRJBRG1TGydEgUxc7SsskFh5DIAsIHI38MpbLajgSNb9b3
2fAOXSL4/0NyXg3appWU4nOimSR2XHMfXjdsR6uztXZUEWI8SoK6q1gsdSi+sZAAZKkzlBzl1032
eUjR2FZwF0c5nP7gQxMl6NXhHAo9SVBnoae24n8Hnq4a5h3bXMdrlBJpNbcPacGmBO5jTE1lJ/mp
9sDPEgJ/iqOIxLFL4J6dcjiu7S0MoZUsMss5uSF01Yhc+KTbkLM0ryRcziafhsEBur/wno31UMPw
w0lmMbytLFd3A8/zMYjCuRhpRHfJSQ94Hn0ULZoFCH33H8st9DFs2VesgvSL+evp8X4zlAED+TfF
OHmhXRJ2wBgvB8AdHU2IaFhgujgf2+fwS0SAe6MnsO/ZD1ftctF+1YzSSALKy+fZNDVgDFWpOx07
gPPsqjZEeEm2uwfgaKFsMQ5DM8Qsm9PLiOYynEgUcFBdslftkeb7qoWD95SF2dv+WsjFxpCJYWt2
4OUUw6djuNAdDoRnqVCas45VXgCcVCmndgGjkozrvCrfr6MP4g8m9uWRsHcd96uYIgKhrZA1941r
/2APn28VvDpDHJhlUgQ9hg1PliNBcVmgYwzQEyRudVWgns8pMRK7+sbvEajxfHjwgJaPq5ngRpzq
g0C8I4fOpcYjfdO8P42sq2skMZOF9nWR1MGFK/yoqxuZK1MuuNRJdSEdJVlx8Y116Z4dO7vcz0QF
RQl8DapTrwe/Z1a+xqlNAm6cu9Ww1s6z2rBdAiLrqkjC+vJ5IS3Cu0IFSQUkM5SFEDDir3Wo1M39
nmiK3UfMRy944vyDICoDN4lgShz3exprLesg3DOLuOVfKxtF1t9LXdT5QJF8P76Um+PyTAvZdD4s
k4jnXiMr2A/Ar3Yg0kTVwLB0G+qQxkc0YAJAt+fOV69pYC/TEcMLOafB6oj25TFEXXAPr8GHFaUG
QumZWSpskrWa6tmO2BqDpyi4SIRNCIDg2D86L2JHdc957u/rhjYQcjaErxXQ76EW2O5NNaJu/CtF
suGaiOluQ+5ZAo0DKBggeCTmSyIb6Y1RlTcpQNcDU4/CX+LC1s3QYeX6xEbBCNe3PXVBgmcMehFR
6zV2VC4MTHVU77G9JlvA8t+pM0BTWmZHewOzxByyDuQDKq5mWVTfTpea5vlIGivSoPLolrp87PXg
sctQ1qOFWmyRmZc8orvkpc/ocKp8R9KkufFywYs7xsM4vilR6eKFSHlxTtMRMZyh0cGh1LxM6JvL
QT9jiAnYY47PJL6H7TXEbo4DmdSTzP9uQvx6uPmvMMMfh0l6b3sM9NaL4wqBU2A8Jv0uOjxul8Tv
hXSdOzojAhej08U0MGmz+v2zDbhe1hssf7J9lZNRpPQXAuuSVRHLghlszgVFWfKIpsh4FWf7ziaK
B0+sW2zoVKI1b18oQ5XrzlXq+w6LWgvg9K3nYgtz2oPUq6ed/NM9zks2Cv6wdF5tBWH3MpCq71gT
NAKTK/+LSAfNjNtkOEdqzl4bqGLjsTMHc9qM0LWx07IcSjoLv3UISMz3TRbzkkPE1XFnaMYBBytO
BRMVNhB7GH2DtSJSMsa88G3rUeVkIclsO9gV/BWzTndZAHiaiz3+Q9qyqLCxWZLnQkwxmkG0XVBV
WUVdJUBBxjuI+iAKfJwra1DSikp0D9qtb4PPMbnCEL+Dy0bAdddkbYKI7cyrAWfeg1UV3zEONvXq
hYR8H0JydurZWXHDPXoAM/zeuS+ggw1IQyoW0KPUrXREZs8uvoaNTMa7fPXOo+LJ6uyyEnTDLdAf
VeoLJ6rdmJQd+G08aXnE4Lyo/6dQUQGaxV9Kl7j1fMSrx2GrN/rG7fAXbeN8oB4Fn0bYhY1FehPX
d7xnIRoprva9ZVLOTtakQH/du5WA4hEoIQkge7YzvTe0H0iPJrJ/thw3y2gJWY7H5LuIYGUiAp0u
yF8Z+k6zuei+0zuvCUrnMW6V96PYNYmT2VBINv4Qx7I4s8CvQaTmYJEOvZ55lmYxFIy1sgGChS7J
peMEibkwjw88/HbUYGfiOm57BcUArXbaL0HLRb+5AlzoQxUbdbvbD5YYcLoqQEcBr8Tj6EGgFDqT
GhHTcXIjex/T+fbMxlnryqFjDvS4n9roG/5/gWlFX2DJLJ32cl1V/ZmI+IiFgSzgEA3WnzOOFWEe
t5dQanJKc1fUWSJPqb6zr6RV/sgp/0Vq5tanPK6o/YtaMiI3U0SKb+cmVb79f5L4ktTsi9K4haVQ
Fbhf6yMrwm/8D3QytUh4MiJCysxaR0SbrYJbrpeoK35bDSeSWwF/H3tB+fEraIlO1p6CZWVFNykb
EcPyDqq2+BB7w3OB/1KEsEcahqR+yoKkmxZkBtvuYnDMtgvkj9urJE3iB8NB3Ri0/cXuqJpXPAnm
4r4xNX6vViLbEFhY5C/FT/f5P6ffe9EJLsS88mzDjHNlF5jE9uWduNu5/8mbRCvA/z09K1FPsPX9
xwqOVXDmCt/UH67NA6AB6xOvT1CzbRT86x1gaO6DXUwiLOrVw0oWPLN6T/m2uMFMMu+hzI2sPXTN
u51c2e2txRSmHtjywOE0IW0tj6tbrxCGhrpL7qMhRaRgKJc8fSsd5aJQuVG0a9H+SjT1sw/MzFMD
3iBHfthrbtz/Q2hSei74IZDwkJ4xdxrIrHD7bQwtf5NDRs5JECPZve6dbK2jXblLmq39SlkD+Cd4
IMX5DiGwRkD9VYcftZIJIYafnAtiD6MgHFqDZKqhZL+p7BxLorTzzBjNx8iYLWbSy/ZHZepjmX3J
hbzRlmV79lvkWo6XJecQxNWyL60Mcv2CW9JJm5aODv2ezOJC9lJ5TSpJWY7ojBoXUiYdT55DgFDe
ULzHlO2nRBbqiHsdrh7cTVGDEMrHqh8yHwc8zw6srglqCllU5Xwry+AF1ZvNALzhLxiLlZD5Sp5Z
9ARkY35O7Q7RPBLSXjuV6XiUxK46fuZCl5aFFt2Tdt4btNTQRz+Y0WuZ9e9LdEApW0ZPgKnNWrOn
ymQmlxNbAonzNlao42QAGs+4nB1ufwAphSx74XQoT6jR9LziW7RbIfFrC3OVQFIuvgq5WJIJj3Rt
ddEcQ/LCGJge9+JxsYHqeeoJyh2TcNUKia2zJnxoYO+ZDlumUXaUADpyYG35mxMOCqr1MCi7tWYF
gP3lDQN1IhoUQsbUqhy/GQtg8QT9y40JMskLDZ4U8UI7Tzm+H9E7syqLkGZW/hD589xHJ/vE+Ept
TTCe/J9IDWtQeI0Vfgnd8Dtjb9pIZQqF2TjzhZOKl/zAZA100AsuPCgGhEbYAeYsHKkJvaU9Yo7x
cZwSkl1aXf8rVJPlKgLbnGXpwqGZbkn8hMqUjd43E+L2VY07XHjn7dEi8x+NloyPXHvFupmm4C/A
m/9aQIY2SP5kHJPTxl8cNRt+P9Z8job6p///SlIDORxi3tot6JHWmYBOYX99oMb7SVap2TB9TVQg
KHb6waBVjvBfxTNJAbJ/J7DIfZ8bljTfkindiPjs2Sdv5h626iLSi+sHjrCvbNZ95wC8WemeieqC
PUbBrwCRHlgk+7y0fwJHPKTxJSm7fAwXlSztsoF2jIauCMQGzyuj7965olndC8iCihp8RBc390vv
EX1SnK8ud3nvjpQIvRMHX8YizUaHxohLR6WUkKsUqTbkIl6DEXZKGlq3A+KA63h7+0Kgv6BeWBi0
A2zKGM4tw40LCZShZPa75c0167SWczE8A7B1ixZpnD2z0Imo/jL1QODFi4c+cHy0klONMTLqnNgC
bn4bG6oyqGX/dS3D86MW0vHVA/GNdjCRW7OvwjRAM0w0ziDJ7BxhJ7pLvA9GtIo4lIMHPmHy0API
pbbsGma5BBz612WUGzHzuOn74liI+H+xsEWQdf7/QFCY+JastZa5Tjr83LRVaDHChwxTfBQLmmiH
DhrbrrrccU32WsGXoX4UTGgWuetU5VggP21JiBW5NrpdYoxs/TX+9rojcU8/aeacq1WqlA62BqBy
sPei5i5M9pexlBqi9IO2maDOI41+3ZC4Nn9bNELjz6PE++qR6j/aMSwmHsyfsQV5DQJGr13tLAFR
h/PgUtl/krSb5Q6v9KjoXLJgEcdy3Yeie6mwSuaIN9RWixI7WrOLti0Wh0UVEpk0SLZVTwvrJgKy
WziSFvT+VYnRXS7LeiqtSDfe0GO7cuqmtVlObXcVJZ33BSxHey75bzBb5ClYH4j4wUwc3IS8T4PD
/zBdsjhMeSV84C2XvNGGHNZbrI8TGrnsTF2GFTJpdOPumZy6tra3eggdO9OEnRbvICEQSwVeqOyM
HwxFEZJjI8lwZEj7pDO+Aohqbl+LzUzqz7Vc9lOEo8rBLnyVYkPGnZmSOcQlhDVk6GK0MxF+wcfO
cpnOXo5DlavNzLb3P7J+WC2ytAjNUEy2VoiWg57VExMKBBNrMpxf18SWtU//rYf3h6hC85UarxuG
WSJ96SRcrk/0C8PudVmdhWw8SFvi/8XIesSJxHu4PAoyj5exZ/zw58moFnYlN6ZUvIIo19Q7XSCw
+4JqDCLz7lzwLg+5CCA4idR5tLujVDo2Hl7W+7gTzrhoaRXDTNShKwmFXSFtHampxn7aoQkbHelM
v4Rzvs5ONDRSMd+7XoPivonX9ik86mfGh/ZJCuWgALOdc77pEoWbelNnQV3gTDpXTd3wFje60BvT
tDMUx1m14vt2V+itW/INnl404ITCkdzm+9EeAglXf2xxk5YcfOme22fcWzVWywk3Q0l/oMUGa2Xv
6mvS4fe7mUofeImJneQTQgxzj1LQHP5F38xeur63QHD9JPIK3zgcK4Yps2oZrF9HP8Uh2y7Fp+QO
LbGC41stROkFnuaf0OEP+3Khc4yl1Gvtdv+B6B78vWf8QyvX/8pIaTcIGH5+xVAAAB0l2hLdBM9p
oYwHhnVZfN88ZqHj+/eF5En4fgENjTcPXFlM9vT+U7Zg6ugt/AgeKfAWnWPFMNhidh30rQmKDr5b
oQ/SpSBR8hawzfdAjXNrqB/aDN3bAQ72BXv2qHPnDQkYUB3OjRemvurS/d+H5axSoFOyTCPPisxv
+AYoa5q2SNAVkyLaQ8bVhMsxtwSRRnEur2wZVFq5IqxAjuMoAfA3qt4ON8IyAkz/rwNTBvmeSuVx
v80XrfUMIIsHzDT2xp/Q304O3G32Pz2D3dUvs1ycuE/QLlR84AeUug0wC5vJjiGxZHjBJxqiMrhC
/uxiXeExnV+1X6dwsQUgsyJfVSwoS991azjA4U54zmPojJ6CNcDbEMaxayefP8ZaMjIgL+jM9qUD
Z9HgfcckoMvp+hNGj/+wTl+bxPMWW3v2/xst+i4Q0AzM8GS8/LssDqJWY2Yle+oK6pIU9QSEvuXg
++evy1b4ly8GD+OA+XvlabOBoJRs/eJ6xdXopeCKfyXhq7JPEQiqMWEh/LgDgJbvMHPdfshYkArm
30SWVBeACl4ZfXbNJZBq6wvpTM3fwXd75m+IGpJEHs6Zo89B5UvZvuBGrqBkxp7rkwuPzm5pA234
+fvN9EihhpfyfUF+Gv6vxsfgSDB6iKHvgyvUoFoeNnJgBF2ufMTDXZdSIIBlZecmpa4NS3iLryhA
wdZp0IpA29+89LOlxJ0u7Kq1ZdxcgQ+ltORLju9g2VtmvN6dh/nPQIneL5Ly6yVW+qJCmfZl9Oi0
OOpCCoFNCOTIs0nG44Hu7Mv4C0Wny1VxXZgRsMvs75YnZq2jfp8+yEay+KUSp0o+CLkjVQ6/Ivg+
/nOOwnl3+eHp1PtJ/iB6/8+avm7AkjyLNtepiUnmPAHPoNEoYDa95n34xXJHsgcX4iV2po1/8jPA
T8kBfI+SB/8UPQ8hy1bNVGPOfdKoHWnoFTx92O+jLEededNSedfNzivHmOT8PfNcWSHv8olwZsup
J7kF+r7mg0sufWvZvkb6FiZoBVuDnSG1ZxnH9tC9JEj21Oqync1pu28Wjdf+5TItPAUGm6dkHoW2
e0uqynDZVKOK7E1tgsM2jUkh+KO++kdLqppHqrXQVAUnLlTQUZos0CnmDtXKRPjbRhv9faYPew9S
131ElXPcym/kkT8dVQ5pt4/LyPETVFuTTwYvebiq3buYREbZt1TR14IfAjDLoyxAbu84gcKI5jWd
9FZ8EC9rPOWdyUy422mZ/VB5Ugedfnn5ee+QdDftgxVI/C+KzGlKU0d+QIfxSy6mfS4eXqOswHVC
cvcNQmH6j29Ax8F8DeN+As876345BCP6l8q4z8D1rDHV/9w9dB8UlDphVKK9SWzQ6gHs5ODvcqz4
cztYKKnfhOdTQeUGy+yIXXMA1PukjVpiYbrrDW0qGFizWuU7MJHOFbJJy70QGF381jbCA2JgE55C
BuTfyZqjyKUc76OOJSpqS0+I9Mgl6vd2pgk2nnlNcNeLzut1m7IsJMMLJF8433VSHwrZtdTsOFEi
tLYTEj7IgKeQgzrF4D7EXJVYi9Xy7Dvuyuc6RLOvImgUtRFSkgeV8URcDHed+qXU6Zxy/zQLFqX8
GkY3/vAvO/PYsQvZOs2cwUyGx5VXCgBmdsywEhM4QfJnC4JBTR0gXFUVQoyQd/34ioZbFWY7RNw6
AD49iS/rJj7I8pK10buB6JCjYDCPS6yq9NHBJnupig/jg/8fuOTTELumQDOYek0iw9OGEpchAfPK
vAJKOzUTY7jMvjRmEexyRb7+6AXn12xWC6Uj/IWSlIGWOsNzV7wIdj9y/KsXiJskJJke9BMhfNgZ
w5tjhPj6ahPvDtsHqs7p1329KKDhXMczCaItzHT3FRV1iZFeFaMDaTgLasAbQ4QdA6ezhzLCOtGc
qEkN9tHAdhA3f921FqY9KHhBaQVeZVAZa0hBuxZr1kFSsC9/o8nAbthg8U5xAQHQgjId+1rhfaUV
1//J4uVXIsezpmKdnCUOOylM3HQbiMuzvf8wOiS3z0xj+IECt06e8aVrX+523xeYghrjakIA2Avq
9sgKSVXQKPnQIbmUbdNXiFA3scqupnJ1qrQJFEeAeK3jUJiKubafX6eLg26Qq98oFpSm5lHk2BvI
p9acS17Z1TN9eRqrDSvS/jsdS4ZoLnO+16UPdASa27W76Ny4mELKb4fyu//E6gJeFkAu67YxrURD
KEi7uwn+/R8ZaZaj62roRO8xoKRZX9EwtOBgf2eDYcLCGmZtXyXt4X/faffTQ68I1iBU0aj69iJu
3RXAFNos2LPCSVo7W8mR/X7ugWsbEEEPr+TS8SxdG+4SgyDnJnyv8F3uPPqZFj3PizdoGYitzTW7
bdKUN3qRVthYW++fpf9axqHeXEdJ8HmY1HIKT1exBEogPLA+4xdf9RKGP0YRPMf6OKsvppcYUrgj
dZn22y5ws3YCVHxxM2kCvtJHCLFDEy7k5ZuuF104V/aVKMt9R4fK6IUPO+aVFS3C7IYAKbQ7NsZY
TUNMu9wsNVS7kJEfuR58U91JgLZnwkWZTq1zbr1bJS76d3z6tw3hWqwPtfMr1Wew7bhDrLCgSPCc
YxrkpAzI9fj4EnKMoSDYwg6qnw3tu6qNrR58SoJsRgCK6bgRXi1cXgX3bifJAjyxWji/6jQJxSJI
MKRQl9+jUWjuFK7FxodybbT0KlF/NKMzaLJnjd726cGINHftPrbDFgiLiKSO5fsU6g2knheViFaR
8dMpNKTSZfHlFkLW3//CZImIUiM20Nr0Vwlp7p3tBdUofI44vhn8u8ZCduqwF7UtwmnNnd00kgUG
miDgQpbebulpY1xh5kR0cYO3YHCLINAC7NXtbRLO4u9yC0Fk0yr9bOnfU354vquDN4/WXl3OepD/
JgIFPnE+VXWjO2yW3Zg81erJPEtWnNfPKhspSNqRCdkBt9FRQXUVUyAs0xPGCSGYMi3vVux7bZgy
Q6nv8zvXdPDBJrl7J+dYTn6pptyw1ANhOTd6zARAZ51BGef3lBp8quzr4LAzK2jGWJIkznlbd3b7
XAYTGfwb00IgeitKo62+ql318hqzJM29yn5ONrSzXLGvgFakqB6N6eWh4hDJZYU77TlMLiTFBfBr
Tfkmb5wRAnZUitoWBdlN6zAOGewNMp2TtNRrf8hHGJsDp54TCEfixiEkm86nKcs67bmkP+rJRr83
ZkbOLhXnMZ1lWla5QHqmjkLuzFlLrr0JMifDqt0GkXRcjQXIxstPmyGWv/gtrj7vkCuFIxxqfTyb
OxiPOQLiiGQblZfdXG+OcF95dg2WNqu+bjM3lx94Lb66HMQkasll83Rd9Kp0wm3jmN4Sdndn1TJi
mpJTn9wOP+NBEO4BdLh2C5sb6GuIXW6L3vF83eH4N6uV/UytosNb9C7e7RcLdHSghwDDidkOg5dj
WxqyZLOU86dO31wg64YiBSjy8Pt0iEkNEAA7cUzCsf7gMHHuMilYndnDTw0gl7Chqo73bK/hO+df
iH8b6233uKStEa89/ajVaTMMaKWhxr7HvWGAaU2hcS+mWW5Z6btwxM7v3dPBouxxaEUGhmZI8CQc
CuuAjaZYx58iJGM4wbiTmqGGLuhzlBlzznc/xiYw1vl1x1MXzOKayIVDNCS4pDHVOLAGYABEtJ6b
e/VLnRKZEgBk65yU5e3gKAYDbntoT2+/wiKgGzpkDIXMeDuwtTJrAKp4IOqB1EEvlgPxD2XYhFQ1
HGqn8c3BZSYc5o28Qa+3tUp+OpMGqoi0parSHMLo0aA0Fpcva/pKBLmMXMKaA18fedza/OvK9sDx
pQ+LXldyL5GzRpglnqJfAz5jaUvoaTlpWRnj3ik0x+H+wLC1Kdoyt5GlZJ1HcHj+Af/PugGEperq
weD0Xd2Qwuz4okx5kx80dNxf0mhMx9gxzJSuMGh8bhPB1gFUuI1efnar0MbQA8Xf6oMGnU+I+kaD
NpkE36J3H5en1cu5zUEkIm9EhdahkjBq4R+T+jDbzIwAAu1ka4GWzIj8W4sPxS93DVApoPnIGwKy
4uZ6ApHDmbYZpCjminbLtjLv6PfIMXTO0xrAsL5aEswunxURdU9glnGxhltvjd/07p0i/oBHGedJ
DSej4W0sr21/8yK3wk86jY0i1uOEy34zk+DxSSeJA7nSy4uBJi4Llya1ecwKPqzTACz/oie59AO7
mKlstIUtv2sO5/oe9H5OD1C9E2BeNy2c4gQuzUJCKCPg4QQ7SiwryY45Ah+r1TmLl7VmsZ6ah8Md
m15PkpEKrqW4F2iFHsnLJ7eY7jQol6v1xH8Q4IVYHZpO0PKrRsHY0eu/Z1COvNzzG6ElDeBVnIzX
BKJko5eISNJTtPqcKRQ7VHrXNukhoA5Se5ZW5Zq8vg3rgz12W5WtAUzXNseGUeOlFPC+8f1pmjam
4C2C+R7YkNVuqFtJmtWGSpEnhW80YnCmW46T0vrbox4y58/jQq0YK6dDP5ndUK8oEjpE4KSNrKoO
LJmRu7y23sjczx4PMQcDOoeyPIfAqhmHJ6OssUtZ1Of/htw9NGT5+hYHNSPSXh9u7Oj0R5Gt3PYR
U3IE1NPzVWKua6d7lj/ch8GmXUu14yChtwJHpJPRTN1Yuj3Sj7GOsNxQFoYjYROyKbItcEB6seoq
X+B6bdgyUqDikztCqyCuHRBLoo4QxInGwHDNrP2ccMGaof0s34ZnmMsadKr67VngsZD8WeR5zgqd
mfJVf+GUc4NIz2mpSC2Y1U23x6SJFInrFDa1hYGLDsxM9jzyTS/6LbLS/XB3E5d2voyGpyxfIdSE
GEEp5IMPrUr3+082K9IIMIl425jqGzC7+fuWH4ROD2vfr7ma22B8T5m/cxlo7Coq9dbZkopSegnF
iAsEGBMDmefwYiaWvRfwcvT2bUvn2FNxIcL/+awL1HBKWpbYgQF9t0uYZhIAGHWNua1nNpTDpHHH
Iz00ARDu6F+qJK2PfXg+BZW4A6knzfZjRvMI7DHZNeAf4jVC1ww0QPNbTbyAkY0lX0sewKfsHz3l
zGYLe21BeQnGKurN+YfvInw8PYe1EgYmZCzrej2NGgPbz/1W0dndHE/I6UQnOpnr6RZiq0/zL6wW
jfhjKZ8lckbVXp3LX2qhAz7yhp9rwAunaLnVNq+tLQKKlJ2IKUcj87oVfCIg+P100Lah58omOEY0
zOq6/8MshZ9i712yVAkw3p82+EMcKmv2dlesQPIz7UKpSxwwMGdD1Fy0RX5bP309GlPm5HlB8vtP
ndnxn7udrrWAJz+7NfQz4oKHsLybqfD/GuIqHUJBjSdWBXUUVUvqNVtkL+aRz/LvaFj4KcjfHW1R
Y/LHduqM58Z6Rcxhg8dM/q95mno0mur2WRA0qYB756q7INsr1VQ83FFZqvU9sF3JLWvXzOZhj/dG
abu4mgbhe/OGBJo76gPM8TG/juaHXgTr17f5nDa/46S6YRyJzMUGjD3gHaVof5oLsinUiKSLFsex
cED/+QyNE0Z72KNFM0FypOMC2LpckGNhQ2kkvW1OLtNXfkZszEm1P35NkTL0vD2gW2X4WSO2SZ72
gE6Tbk2BVkIcV39CqANJtfORZmreCIVW7vteQCNxFg7qvTV02bGc+4LkcHWS+tLbx0qor0V28XrL
1QY9DWTPB7adwWl0VWRiLbmhhEKLoQkZReKP8KWfyD+XZoLoRldb685AT1HhexchBYtQD2Koyrzc
5uSp2Mk+mbBpcxL4kW5rMZXKH1ipxbTGZUAmSXAgQlB5A5HAuLqJFAwx/GdXzrED+CdLbYYK6Pjt
VoUTNZuejkEEFS+tXlIXQrj8Yes7CMeuPhNnKfwB0abgyDh0BHgai0NU66Au7u6YlTMNqTUudF4i
PfUZrXWPn8DPNodV+LgrsGDLLJEgXltMybb3rpy5hlidiIaUUZlCoRekjhfmvXohnZdKslVBg417
ItEQZKnXppHqbWdAUc8TYKVOftnG/dfObrNT6QLSIRSBqbCDN8EM3Ghu5/7YqibzrCciBHF55sPl
S+AwbQGuE+TErSqudkoM08XlriAID3e9nvbhZfXlsGH+GRXyPde+WhLikP+ARQ0JgSnr0HhW8aZv
QFL8QlyTVlJ7iboKNhwD8Chwbpr+H/HuWproE6GjJSmKVr8t3r07HKmVyItsjX8lcb81KpodqZcr
a/FIAI/YOE3BtWw5bs+/NN5XjmbK5bn7nEoZ/YGCZlvmRgGnMDbGlqsVJ1WifJnDBCBUDQ8h/x2n
BQOQdML2lMHXP9tuAvZO4fDkWoLbNB1L3GiZNZZ0vrLpxVhXtFvB15j6ue0gxccZJlgWNKVJ2wGH
N2oY2RhSqRJsx4aVZdqQ8LaNskyuozRSi0WeiImdA/3fpHcqvnTqZKvxO67Rm0Ray5B+bX6sRqAO
i5/ChS1MAj2wS1oiC8jpiIYNRA/LyaX/W3hIg1E9WLLH/FVD6cvQ9V1AkyiKaIgpXldSEMKjJXWn
PGmJG9I6bYygM4Nm/ObB7YYNqGoYiIIpHRc0c35w4EyCASNZcMYceotRUyPJ+8aNGJupxE6VYTMa
ERf8/dl8+PZab/rP52msKvrQ9LUTD2h0458Qh4T0o3TvZqnWIvXPGfTNH8WtpFd4kIpRvCu5gTKM
X0nZPS1X5eh0Hjnavu4aHE98W0F1kUL4lFekZuwWf80nAd0hMUSkiD+pQlF2Q7TISqZCXc3qGNZE
lt8dRSQCWzh/U3DfNI6uEyD+wQwOOKnLe5E9amcPlAm3nCUii+DvYEjsIPSsUZRte5vkk53TDhu5
2wSORtE5jVzS62LNRd6T4AkJAw8BaTIZXBHgKRB3G3PbuTArsXCR5F2oQbPAfRbi9W09cHP4ExpS
cqGnp2rTAhg29csj6N5GvTwfTFUH1maCJpwfcPsp6Tu5yq7yXUPrlHWCYPZ2o7jRRdvOkH1Yy045
1MlKmM1nB+aHwbPyh4H88v14HlOcjXrm6/xOASVpJKr1Oe6RBMCatHpYY0OEJX/MS3a5NdS+jARE
0R0uS9fMy6guP7QZWj0QzK0bPIfTBJLnocrLetFCSQkctn2m13BvCniMBMT4OOuKsiRd7u5PhVK7
p0GOgzXtycvnD+K/ttlY6hMVsFKKLqQ88imUuILu4HI0DcfUp/TVD90yIYf8j2iPb25yob26gocH
XzRn7BAgiylzCFCo2aPNDPSltwbAWe09u7aGGPxb9F/joE+h6Me2Q8dpPvFMd95YugcRIXDBGSu8
tEy0+khOaEhZ6b8rr016M3b2K3X38fMaydF/S2Wquhy30wT8D77wKwijV73UMYwPJDLG8kX+Yf+k
j9G7mPw/ggcBW1o4SJLP+Zue2tLW/gvMNRAGyXuk0mO9xE19e2AKlK9+1FhgGwamPzJ6z+N0TYnh
uBQmMh05R9ITIJx1hMIAs40ruAesGbuRL+E0BqFxmpHiT2a8GZY8aZc/CF1c6tfEO/V3tUeblcvo
O4yfQNAiIrzizTs3wL4oye1ftyYRULbGy6fCCo6MRl1q/kR4qVLI06z8oAmgcKO3X4RQuMr3Ckd/
XcXXqDuhKAHJMPE477QFOuXYuOtYowtgwczavvco5O18wSpRY0fNp/gDmw9PsbBQYtmUXhG4vH0A
SMqdA/YUZr3gcAsoSGPxI4nANSJIxps+U0lphZuyRLvGH8hrEOj/dSWYKJLkPteJNIV3ickhGnbu
7pCfYo+IuVNtk/0Ls2nAAHreHxXvgHd6zCCHgYYLI4blt/ziJfIxQVOrUpn0LjqaLez9yC1t4ie+
zeBgnTPWixqFRS7MocqOTwRAUX/kQhjGNirypf3/td3bVOVxTC7TCkvPIJyB+XkcN4/3Z3lQ1ULG
TXUM2AWE7CzIXgVBnzq3B07WzC9Et1l2ijBvHzQpDnDUEkqQLqb+m9lzFMW+zQkb2KmNtjHapPFI
kKuwPyqH5R3VChAld9diIietvEw9ZZDJ4GRI1NDaB9dIl1QxwWwHdN1AC9Fb+oHt7XBwfwtCVj+6
UM0KjLrgFxCcml+jSfOT5ONxzUQuB3I77jUzi5JxQfwzuBbEfHIJkkIp4SzlHMErsW+lQbvWCaBg
cMIpRNkp/lyDXjdQuLtL8NzF3E+kG2ORI/j7ZF4tLYSDI3LBDLMtclZnFeyCX7M/lP1ZoZr3PG/D
hVKo6WgLpeAtgUQVZ4A/s4np3Yxhq+DY1bKMMEhsQ/R+JLVzgQm+dWTiucOVN94Ym7ExF7OC61tI
2QmUX+exiuMncevTc2e6FR96j1wV2LPzMxbgxOt8he0nKcFP7ZdnOlifjgLIMp6nsfUwWuT9BD01
/zgsf9zhvWbPz8oTMvP3/nJjhwu0k3Qi5r/GxkAduri07te+s3tIZNgx4CXIhUdqeCb7RhozRavH
9zK0mWz8pFpCco6o/QG+Zl++c0f3+iZmKlusa3VjBLXvoaTZPdLhmYAhE0fE1Ewn3e3x31iGbIKA
UyntE84eDpQhI0dtYI7EQnURbmS0pkx8bTbxrM1Xo/r7OJMeEYMpq9e4JMENlLprUVci/XbJ7Ils
oG+npZAX6Ziw0VneWoviB8peXg5aH66zOfVm22I3BswuVmGCGvwvlp9EU5tOAV4XG+BJjsRYmy50
/UXCN2C/bkaxn0to7CExAcqSecrr8zCmepYrzjQe4386J9M+2EKvONGYwy5w5jkg64adW6TDpIZs
3OIVG/ON/r4IBU9mzz/5IUAYJOjMPEoBJNGbbNoebG5SyDSs56xxnjjUJWsUta4Kiwyd4L32iKgW
sNJE0knguLDeCI560v627xzkkIhEdRUhinyQ/p1kDy2gdlp1XPD+k2jpvFcpaO/n2mzAn65FfDwf
7zbEAJrn9tbyYea72B71Qu2IAzD1x+Suh/T9KpbQN70I7u58laOAutwjqpGxKIiLxBp8M/QHjvFH
03qu2nDMfwQ2V4g921hLizjsFGMaPbLDtxc/XYDdA5GEAIvm4IzsS2UezObn2gId7nfygtRLC6nF
hev3YCTLxtEexE296R8rUqQZVBrE8QAkyPSa6yrbogeBm3Xnmf4Z3gcGOofMj4YbVx/5lFattslc
8fIAPvNANWmYQasFJu+66e/epxwqqK71PDCb3yck2fO4YnjAvOUqMFCbsHJ85hltbTNXRWdplnZ8
ovL0FYbuR/3GWoZ9l594Ho3UbU/ROLUB+cIu7crByctAsG2G4JwL5WHUZ6Ov+ABii0f20wGsouYx
fTiUdFisAmk0iwxJ+Oi3+XeD+OcCBFPZiA2qaCnL/itnkNUJ/tlZ5yWxR5UbXXsqtXnNUtoUgQNI
wbq5O9/bSS6se+uDJWMU/Mt68hOP+9Gnf7kzjBsgcZ0uRcQs+8ZElNscqS/CV/D7Hu6cF2DTONT4
ZidcbkDpqqD7kFe7sAD9EghMqBG4bvVOcu07m3TJ34wIa1OjwZRAigiCRYOC7m84gjyUlVWsDE5L
T+1ouUf8gMUaq0fsc15xRUzMoDX+B0wVzN8izmCm+tSCSM9aOlVtXI8L+YGAwtfRt7oqgKaSjGDS
y7F/BRMEnDwBSMiiL8mu/Gy+rYIgI5i9lRiiy8GoxiGIQusSuWVilfiwSwi1oh1/ZcoQ7JRSSfm1
Grgnxa3GrFHZRj3s/prmBKqLVf3g695T8Ew6QqzgCdM0T/b0g9iQ1mRXhxJR78Us5Kvhs2mSsg66
5Yy+PdtOhqPE0tHUFnvAtRMdx0h+fs5uAMiExrNbL0/6lN+aBn8UK1isfJkK2P48GpbYQSAcfPHC
0Oqo1EhjfV/f4D1Gfk8BMIR6gsZPwU/HXSe6XFI6bCqghG0nizmkw0RQxZtyU6sfI5jxC3MRi35T
PMLeEXCNePYDqjjgZvCXwVIlH/039e6q4WgbeRvI4gr3BEEfihUaDoxdEqER2le0FYGZkdI/TZd8
m3Pxnf2DMW/SwsDBSkLek7wbHtdy+B5bafTRug5CO31UdeqLD8fFZuHspSEkRLGYPvZw/GvHzxAi
PbuNO67n3GrwhTku3fH4cMHqoQGtb3PPZyn6XOLmfFngt6OcgMumoLvniAPh1dM8grVOvwiYXTwu
KN6+pYXvYqvtuccta09BUgbrn5MbsefHGvRBlmSGRyLrowNjC1HGYL/+AU3/WetWMdIxXpCVs2mp
q58jvNsySDaDW37TbFp57Dg5Y+ov9cYNWhZ82IM4S+BdL/C3Pr4/UULJKqch96L8aXzO/kA8mx9k
dFE2zseCT9DWyLWa9VBj0FE6HwzYjif/KWVMj+6vxlM5W4mrEFzcPFPUryb+C+FOZgWCDfDY5ZfV
z53wo/3ajsAowJTEkh3rWZnQAhaDwIGLGKQWABF0rOtH8PfS6LjIE9+G97P3KH4+HooyJwdwyEh1
kThWV/BqqlhUXTaqyDCiNvsOMGwJ/dgOcuBF3D69Pa7uhq+DGzswBipCe7WG6VsP8STlKkrnqaBP
V8dwKLkkyCSUYglmcr1V/klTlLRFfkC39zIPnZ2aWvSlpxof4Hio3XjFShsyfe6ufRoUui/mBYWW
DiTdZF2rqp6zxaEkkv3fzUpLkEK5g6XmcuvVaOwGSBZMsqVbLDCiaMsw8KfkKBBvcqCUbRW1mt9e
T5bJxxVxi/yqcKp9bpPtN6LfG6eJmebDpw3Rr2W5D01EvPSzdzayEVAwudbhx71uQZsdpn3z1a2h
84n9uV/Zv6f85cV8CeO+O/YKwvddR53CvIVsE7tvxQ8ACthVOaFMGM1AZGGbXXOkRUwzdjCnpgI5
yYQKSYSNcIO8aRt17ym9q7vqnziMNdxNDjwr3MF8pHKii07hN2IVcF+S4cLgQBfK9VQhJIjQJle2
/pVULOo7T4uyRyG/VAVStZsYfiCjB25/L1sBCYmkDV67JcGkVOq3+bCbMovyt1Blj0CUQPJn+JyD
ump0pKhSdcLDGu/lMtumTTDielbCn5krHiRwDgbLj+XFTg9xR0cB1BSSHGjDIrxpldBQNSweVufZ
JaeHUjjoOYWSthOZuZ4JMim0ZjpP2YpNaYvMy09z13R1ZCPJFWJSRMD749dPwsxBlk4XK6W6iD0E
ziOLVdUpSpUqGAVXw5k/ty7SDjxG5C2aEwGJ82TVrnE2SYpLRVNSxv0PnW3PPR1eIeZ1D54SFnZp
hlVO28ofpZhHxX4IknFc8UJT7VA7oxzUYoX//fARdHas+o2V9jofGlj1gEhuMn9TCBHKRmppOjHe
d+YcnMoBFagjfgznjKU/XJPNPfdzBcr50VI+++jTjNbgp6/liRuZoTcHNcsMddtqoOoedgZ6gZtH
UGALkvP4naMHuATxAZQJ6d6pLlQWZ9S9+u+W83/QNctDurMxMK/V4M+qJC+Urf2enMOwZrAagxUX
9mpP1sTcAkFeN7F+NptO6GORa21KY/UIpsWr0yGijasroLyg3LHovj3/ODaLFcGMSUx1k0LsFq3C
+YVJiHB5YxTJSMgiVpAEio/Jcmo0JKJ2sPIBra/BtFhe/Hjw3YevJBL4sY0uVIfcxxp4c0pPgSLS
TtexuNs93EBji3EhzSjyUoNFhrVFrBXP+sOwxg1Zw682dmop8ZeS4iv6i6ILJJy3OcjCQOI4bVgQ
Rc9wIYah/CdD+6F45xu2K0/hX/Ro4iIhi6M3ylU/rTC7r8sYMw+a+DoozjkPGblIfii2GaEbewl9
QKbKrO1jWgo4+L+7KH4fxRJemjZEybLeDbsNtIc+t40E4B8MZ4fSpI/5jSuCA+P44KV5ijPM4++O
2wB1RZk2n6aR24qbqh9wm3BDo7jfBRFc/Wt1qL7LgX8uLuSCk5sv6TT3ipYu/Q8t9BjlKXabtXCL
kAyqD/yoKs3recymd215Xor1lQngveRRVebEXzuUXohdX3ccKEvkioIysX92yvo6wwo76sW/EhH0
HY3lw9AVpoVi5330hB4C5iw3aA0b2rrnSqMn8UszBYPMjSGuXCmkVNY90GOhqIQzjYkYV1PbBoRm
Tih1+ET6MEyc/2ypZA0KYNKg39hxPkeWiOV/3QNw/KWVmkUp3pa2FdHK7Cj8pGH6XsICV1kLvuf0
43TVpO0Qo2xZaIlMTNhEEmCgWFjcTyYQ/GZsdvSLstBLgzF0FDnF+Uf8yEWGT751hyj+uQkSLmUU
F0zhMjFeoudbcYWxiIfC6X7/UvLeP/szZOpax7O2BYiW4J8ZGkZYc4FI3LavoExWX2anmwUNRKQ9
H8OhV2kz26Wf0opI4b55QcoJwO9K6Z/t7Qn8VQW/YtIC0Cpllg5SijBt4Q0wMMXmi4y/FuYE7UbV
+BiRsNy5R1NcR6aWMyeAC5bWU6YnDZA5PKxsRnULlie9PbJM9Gd/qZIIq8Vk+5s8NNS80evDx4qV
lOaNFfGrbOplyynoK60hRqpKnsEWJq9H61s8phRDVx0lcCRyygUazMEp50CxFFs0vPBclPk8H+QU
xepg3OOf3G41UT3Zxl59Z7oxk2DaxuMyP14wpXGv4MmFzVmNCLaN2kitAk2U4oULxKd7f3Bl7+nm
k21vFefkrfNn0vLTD0blSkxmA+QO8yisgUpa8rLkfzc1RZnTzzjEHdJxZ1oUp/OC+CuJcsSuV+XT
dJlQVCQ1cyCiErWNPgG7bB/1hWzS5CuxjuaHQ3wAe7V3Q2Hdw1ZxDzvWeIOxjWgC+QMt2EE+1iIN
vVZ17lFMs8l1xEfoAd5R9vPQmb6NMSFGVz3q9bUD15nLFh8UVs0Tfo3smINI3Ho8dMBwIvAO1E7X
dW4l3w72bh9AO62voco+JxZzRcozc0SKOD7ETiEJHRGAZQqmFGr2KBiBSBI7qZrt61dsIo8LDGXE
HLDDw0pr5FUYKAZxwBbdSoyXcO2AhDAzMV+JWENz5hPxVRekCuc6uMiw8SUPEFMJuRVEthbvE6gO
5YHOuxkm4NLaUOANI2nUZf/EtnXaXPBaa6YVWa7swSe2N1a5KPDGIPp+bjPOl72olR2x37l5Fdt9
HMDj8zGL1DaAEyd/GShUwRltWEgp0L6uQk52VmZgEKlQ9DPrkAFmWtwFtl1g5svY63fxAhtHeiTH
42yJsx+8pbiP/bYm7/lhYuWlpiUjGDKhZ1v7rLO5olOOlc3V3eSlIBx9dDxpJIoGidtiX+OrChrD
5AYsuaVaE9zmyn4mIl4bLWQhhnkzbVy9wmBxeppoFLV4Bq31heK9SseVlEqutMAtVZKZMuU6u9Mq
FvbEPMgEleWGLf/29w82h8fG33Fk4WqkP19gwKRwjxwTT8uk6H4fY34/kP8gSuzIdCXigCXN3o6G
KqnLG3ZQoTPIulZvIhxvy4XwWd2CyUPfhbXGGqwUFlakfKuMBF7xzhKrCh8UH1flNByNrbu+vG+4
Mwv+thTomRECsiNvBWmGxWqqj26ErX2i8Sg+/LcyUY7AJQVgGEuFI+IpFwEg/LKoRNlGD2IBzqnx
g5gOFYVTGGIqcZ6BL6dEdFvhUUnkNetiI7Yher7UgCbHWmIo38FyoRw2yoY5yrTmkSMZI5pQf7Yx
fLEkLvNWPMTWZGHdZNxkXNJWJh+XVeN6PfZk4E47GcsIMHbWcInS9cZs9fhDmQNB1nMdd96vFO0m
zcVGrKUv1vE5o/b4CIGO3WHoXsFDLX2bYEMcGifdFUVInFt86Lklz39rkCughydmT44Id14Lsna3
3TlLLaQOyUZ6KzM7RkvrbQq1FO1uDsrwF4FgKEQ20JTnFumGXMjFdXXpkf0p1l6EauzFLiCkz9ZW
6RLv2g6XFI3wyJFFtowi3d+64E9Lf+aNzKhNDlBp+ybfez9QR2Es1jDHhu7ACnl0axljIKa06Tia
FI/CW3OWytA5m3ckV3dHgSIRraB042eYX6bPmYLkMaWBYIa5wvYb2IzMyYTn9lCEmC3Xuhl1tK5M
TLL1sxIQhBmrMBjxq5ntI1JsL4FDUXJGpfiYexQDRTPIY8UsJKvQvY+0gUKTaNDh2QI0AXUG1RcC
8Zszn7L8qc7b8GFWBegONChuo31ICKPe+5PYi9XHPdCl49+uWy7bagjpAOfUuKHsyyERlTvgIjWf
LpjUmcolEAsZxgiTrVn2u0yUKykWG5AZbZJ1lvjdBII+lCJtZhqJ7hztP0He/UdPaJpU7xtqYcKh
Alogw5XgBkrsjE0pYtYYp0KltLyRZjoAd7c3ulzS+qaqo6ZqRreqmqxghMvg1Poxo89spjnpCTBo
6eN+EjBEuj6MG/9+/NVzGu+xA4SU6O0KCg4ejHg7jMassPiJLaaSm4sPel8PT3zAbxlXhJzScLin
CW7vX0GJ2jSdsdW0XkuLN5Z+vZVqSk7Jipo2BMh+9Q3NhtgR0B/n3h1DZsBynkor/7xsz5MsA5u9
kp0T3Iw0lSMZ2nmtEJfC6jt3Hif9PixgSVQ2+zoNYxi4xTGti1DMNaL7Utr5oGqiRx9UA+vq6SRy
8OIZZpSJ13IAR/o+Jg1a7XEyeDjic06fv09uJB2fuUEWvGXyUQSLU6CVGkEgjuZpYC8d8RqNVAPT
HC5uvCgAP9C91PuKRFXiAlXTEehfI9NevFHhtVqPxiYjrgylMvhunyPJXCE0iimAtREHQ1aA+qSh
dvElZgvMq4kidGLHuYHt3YmirJTPXV7G4UdwNWYl4mski5K4nz+PYtGbOctXLkyK3fWh6xDjH9mF
d39VXJg+BHMt75Or0wImoBYsHdjmhVR7tMk38sXVYb4nYQKiQytWnAxpF0cnbfoDepu2SPVEZPgZ
9ox4hz3l4uaCQeQhf0sN/E0v+6j8NqyL+sQ5BMoiz/Ro7cXMf+SfxIsbX9XPgGCU8lQ7rP9iRb3c
BxSG1VyZetVxDUzg7Y3kJhGU4H8on4WdIiwoBs+BnU9T2uSy/GgDquPYLpueVP5h2VjVs+uOJBhH
5Ku4D8T0O5j+KpZeHbzAmzitwqCwAdenvc4OIPCgihAPmKH13llpIO3aHB/uDw6q+bE5S4Zi77Ph
id6ABCrVQ9P6NJtPmuKyj9OFv4+D7bAK4tb78uCG1mtTVSrLohOzuuUiUS1BDdY2p4cTvrTgFZLW
vUQUj1ctgPjwDHOq/YPE4ceVoUVNevCqWspmwLoiWLMMfEDSSmtoeLPdZiP+HaKZG0Rcx7VxxxfC
pkTX8bvoBRm5P5yF8DmGlCPNPJ9ckr81oCuiChMWo3DjmdEHI1RU2g4nEK3uJ2pI5F1gYv4c9g29
LSI3AeWAfnZPIvww43qKhx432sI17wcTudAmG6Jgnl+PntEtw45MAMFv/y9RMF5yfQNDhYcG/x4y
69Vq02TBB1ehfmi+qoHDX37KPoo2U6UZK9fnEHZY+DyOfCXg7REqogRgvIfGouo9O3cxwAzvYHHr
PuWqCKLicXr4Itk5+UV2NER1w9YWez1qb/V4AbMyHx9wSE45LjECDY86Sc9lKosojeR1Ca7f2tlq
kJXhbXiDfiuPu4dB6dWVtkEQT8Xjpe7ksSUFb5LbZA5cUn72Q+1sEWQSroMNEsQ0vUMO0Hexh85w
K3QMtpXX6Zi56SAr5Iwv+VdvysRqLFUEPqtJofNDFKtRmkZamo6MGssu3iycXNasNWNFlvd3S1tp
HoLzona7y2hv+O9+9yqmWKThI3ZhLgYXKoKcxHaWgqiWEPaR5N4Z3SFmXFPpKEickHb1o3jE5F23
5fdJEBp/Lwz4Moc0ujIRc2Ywhlm2SJ4b2lh2CrHm5d8z0s5KOmXUwGIpOJ83k1I88ZJDa24yq5j2
qKvAtbkjPIBD5EkEeyhBGzTNWS2NgIFwgBf2316IsBdVyIWAiaXS1MRFotfBp5K+LmEQtnG1tj0b
JHOEjq2CphCBe80OQcz7buQn+VDqbdR8YfYngsODoyzGHIez6XmbQ0Zo/GFuBpqjFs8Y5DCkNXnE
NQQK67qrR4tpPr6rF7R92CKCyFC0/QEQUy6qj1rL2l3kyhMu/ivyjtBw6M8iFALKbH0HQe88q0Gx
yWM6Dyu4MCkW4g247buKhOsax5Aj0CsJZEHoo5+B3YDier8hD0SczBMhaITVqPOagBV1E9t2Fw7p
xomrDz4J1NT/UQN6Ye1l7EcXTOrLYU4RZW/JJ1zitAXrqg208YkP1V+NleI7nC3v3lEPIG/YPeo+
DyipkJ05ZfX6nTzOvHf4Pim30tPTPQrdvUreC4NU2/xbTt/CcKTieYaAqUv7gGH/lvPwKucS4R73
YrKUznJqlypYhsipdTXsSLMlK43lBV4oEXYEMN3NZLxD+hrK0c2uc+py3rhUxs9V20NdwND6ZyGM
I4UKBAclYOcwjrtl5PLkBxDlGDG3+3SUJh7duqXROB4963f9+EXzkp9WxiL8HviHxck9WG3d0uBl
AlpngeS+MpBNe1ZQwmfwb4CxZrTbVWj/6oIlpqzTs9QaxL6aqkiKOw7GVw4xF8RuokXKAO42lkjC
S7uAl2ODgfIiR9vTzq0J/ZZwacuG85uGqOLPjfTjyydzmORI1RUR/y2KiAZZgCUGBzkVvZU9IYyL
ak+oBMPvyMe2ZjWIohvoI/2aYMr9EGJNBTAssYdRJ+vj3d/C6pGZV0CLSaCEOZZoqkzdo/cC71RI
7WFrKNvONECkJ0MOgm5y7tn303Y49C1GdUZdqKHcwQWZcu8KnPmdhOB2cPIjwCI1BaWLgJkfSL0K
3KOQNR6cKJY8JhDHh5vTWhxxzdxKi9v5+znxy+yY7/w0Z0eWijGml8fuKGglRMqsxbURtLaYszU/
CyaY0TFhjvVnUsxiRjaAUEgGLYs99dvJ+lg77XyuAQ7If3dIccPZmAYib9/tlnyILtryJl9UPMOv
SgDenp82e+8BZ7HImdNQ0/0loLI+UzufBzsJkOPhTbrAX39SzptcLuYf4utr9Ijs8ZvTpzZGFgXA
oWC2yiSgX8dV7XPy90RORsqtmeyvW3UwBeAGDQs6J0dTq1pTtL1VS4yS78webYR4Ih79snkJQ4aC
vp+BYKnXPgDTAQE/qar2ddm0ipKAtqL2PFyvIz/TmFhKVRg7sZKaUM1t8+eErmpb+BhEP3YrDcX0
ZTNhAqP0Y/KSPWX5YGBERWz6P1qSoQ5mm4oZKn2cA8lwQRLAWR5Iq6BawpRKtUqodYX79EJLy1ou
AGmnBYNGR8fT1i4EnvE/Jx9DYYSfqynanuVR5Ipi1IgFSRIIgGGB0Lenwor7Pv9ihqnwG3lyQEqs
7DBWijXdBwb/G/FYlCuNHx3DTNkjUavWoFeifTufIH4yqwb0bShptd5TYyx12c2gsag8Z+V2Ajd5
jU50pfAbSKOfLCIzxwyqLxpoDUiZbfQZESqhQLpZmAl/dMyxAnMzcqOrVImKqU3b1xNCI+QdOUkX
nuj4WYxuHssQq2QFxQJRtlSxzdYRx2o008gqvQFfvQBL305DduZa4wEdNAAN7bZTJKusfiwfw7bM
xdSGrr8eD+XsyrP+x57hdguah7tUbIPcDdpx2H+XRQBAO/yAZN5jqBeXoZwrHGBlyEGHtZVi6znz
U3Ef+mg8X3BuarKnU8Y5TWco7k3krgbzOVzoGGGCMgxPwUAA2JMbiOnYIbWrC/fylP0ATdPwbwoy
exx7qNB18G/FxOTbQatogCjFeEmqpQ0Vw0RWThHmsNMIb/v++854Sr2Y9lSvmddtL3kOKp1WekXP
UXr4Z14CxJudm+iRPZujyW+7jsw9ebu0ddsUAYt4ppsynxMidlMzNSGy+I/GdJE5Wo//zNWmWtan
g0qOJHeze8Nc10Byr7k2mIVvhf3v4jA7vh68oMWHn7pYrl4bBaCzlnwRwkx9wDMApmgJpMLxX2C0
70zWRXFFLwYSUuN4W7mH1eRm6cI+9vx93YsckPPVwnaFNGGRMkJpbsr0wWG/IPqDs5lF7pRwLsAh
M7X3KHDr6+vgXrsBznf3x4527kAdsAtZ4mRyj/zzp5jiDV4mjCK3aj46sdlA5HfzOl2kv7RjzyJn
hmxx57gD41k9MgBdjQrygJc18+rw0BOmfZZalNAJ5GG4fjDSb3MycvJeY+45ZqYqCXFocsfexFz2
DGlH0qNrSVVTqn4fe8Ke728nFzRucvqDYT4/IN50tV5Nf49hEQ0wG0qFD6hEfueUsyA+n6ZxapB2
soofwMZ82H/6aa4AIsK0uz10j0BVhD7WvP9bQVfO+R/qg6MXfxY8E81cZ3z2Zlji0f3OdWv+qmPU
AzBMt6hipCAytHgym6g3wqz2EhAYV46k+9oxHfK+5ZWeyYJo7i8+iI23irMih7s6JeKJJTqrZxSn
XvX6fqSSPBRLA3O5v2UptLaRSdgQfh+CeIGJmTdBcSKQll1J0pLP49EjsLBoguZvi/y1/UvuLaAC
DJlCqyP0d0+Y1tzgmDnktnkpEfDStJGx1HXxAeVfLoD8gXvGzd/671pKhtEmv0OWPj0UnqE6jECe
ft7kaFpYEgpgm2ZZT2dORca8DAqWD80+o9uBBidazjM/ENLFJohLjkcNFl+IuCUQH4FLtQP5Fv/+
G0k6l3ugzW8LMBA4U1vJmXh84V2GLEPvQwSUxFnUoaxsi4A4TGoVReTXHIxTRYQXVI6WJTj3poYD
RcO/Bm/G4MAqBczXAsGLDtmLe3SbMGl3UeUMnswFh5YABFLVQ/+U5Hai8kujA4J2PGPyWP9NhR11
5hqH+pz4weDlPGxVoRiY5hlVpA1t5fYnPFa8muFIsiZGmK1EpD9SSSj0XnDGbm3KJe5dM1fka3Sk
j5Ho9hhaIwzF9qVUM0wJle573effV5QZW7ivuRZFMQROllX8wAOAbTsIzkgcbdfhrHMTiVTgPXdk
OCMWgTMO1gg4BD3ETGJMNT8hodVVXcfK8V38H42ppG2y/5pt4QVyiVcKHuVaPRD9K3jC60om+CYF
GHB8m04OFRqDe3/bZi+W7yjhMtuB+T0JU/5MH7/xnt5FjeaJpCre1LEtZqc+kn8eS7jLlV2RHyi4
yAvntddjxWW4gahx7lLdSmSvaE4m8D4qZpgdYtisFjt/hrAv28hLCdiGi6+JpEgmURZrH8FW5hdD
ifdls8Pf0201pnSBH4w4Q3SlLRjAKSP2WuXg0Y7ywc5mMjoWm5nqB3BPq4o6oHgFxeYIAAY21btL
Sx1RHgKl8qdHMFLe7ZmYgYU6oQ/9ZfkRzUnTaPdhbwAh/OXTfWEes1XnHI+RwJ2bt4wzqozSqDFm
sRzOC0fe+NJSZ3T0uNA/k8H8N1gVH7pCwQG/sYiIY9ZVKZqUWpQhEr+fkm3FSr0YqRqbhYisrPHm
kwS5WulM1hjtHGlcsEU8jcAbaByxshqNWa/QdD8bQmVj6n3VZ9wzUT87ATaYP+sFQPxm2kpABf9U
J1+huLPDXq4jgVbQnx/vs/AxJK2HtUbv4IypvNl7NZK5Q11194znLHkSJt+S2FBIz1/lNAwrALE/
Y781AM/9rYtI/uXEumurFG/crQjusrv8Det0W+J+QhYbjw6b7QQhboMeHY/j8ountbjfBdn7q8cT
dKaCqCv6yYuzuk+hfnW7U0rZRHCVaAGJutp/gCBaNoyFdbQto8J98Y9goSZTsZHOzaCmfYpMnfRj
Ehpit0Apry9Rj1ycQJK95wdNR1o9wwmM3xYMmTmw/7cSvHdMWfBnqvQJj2gd0fyqVnaXu02RQfx4
E7oITlHPg7RYmDzjClhqJfhrXw5aAMQRNSKLBGemhhtjSZ0Ul3nUX/ClCdV8LubZNpUCT/fsNAr0
zRnbH4e9zScLcD7i/WlGSJUkOwwhgPOOHjKjFKhqwAp6sX4VLEgn8Sh1eQG122g+nJOmXu579wVn
lvA9e9FCm1eQ36Ms41dN6Q9e8aLoucmDyMIvjeEbmIytr5IPUtsS9RVc6c+mddHGoTk4NEHJ3RyZ
q2Ey7+w7Uk7VhjMJ9pkBXNatLrLp/3zhvrUCb2bDTeLb5pD1EV7XWoI6QdP6+XRI+Ws/sCbcROQV
KJnc8/5Xd4I1/OiI3Vp/OAKAYn/xaYdia/MLaq3/GF5gb7GeexkdUAoQBtH1xbTprwBBv+l+JpwS
JDMde9diDdp5j6udun0fJrN/ZKOFsMu/H2F5J2l241uInKJcbv4FosoyRP+Q4VYIEByKkPePpVzI
m4Wea64+Wj+JakiAqXdMKPq0b4hHpWXn71u0053RNhXErAeMPs0mb1b5CtB54nCM5OEpqAo5oabH
UTlBR/P6XSKUdL7NZ0lRVvj8HClb9Ry5vvXJCVd1P9Z1XxxYBmpvud1iqEAgSrN1t3hYSAWUfvO+
9/4mW4STaNHTR9SL+I9lBdflG7rv/K+IjMTQIQAFDolFfhVjYTydJDZ3051WuSvtX+l46YIificE
6zCOWEDY4IFGV/JGfzOPq1L2/LLK+243EaVbNBA239YiCJil+5lnXxRKKjcztrosHpqEXHR0md2C
0U2wnMfkm25ytl9mDuSkSy0/MGzrNfeleIxEOLsmXnNUcf9OaS6455yLsG7lF/X0io3JBvJJMDb7
pNqmxZzN9DvMmQftQp7tJssBypF7DO+4J9hW/2wPs+HdWYDRYb1ql5H1il5o/NCOUR9iTyUkunuY
4DfTPXb96WhrP7EmAV2NH/qHM/1wxXHK/c0ZMP9FMCYOyDJPv3q9BjqbyGprSCn95GrhOcqGBKhn
+F9qPBRgQNhIVVdv/5MLQrB1uR+C5zuwcoaMnguPqMbLm1g95rjYBrMkeh/FdhHj1FFpJ5Gk0Evy
FBu+0oHrk6LfWmGoa0V3Oz+yddjVXCfvgkbwDoP8hKVBrPriwxrcfCzZC4psvTEw3hCQyJcDR39H
NiALQIus1SVn+LjdaqqsBHaECQwIvYVsvoAnyDz+HJwWaF/WIKVL53GSwyF40DNLPXKUSh86hTzw
5hLh78d1lspekGLbbfyLTqUu4IUWQloa3VAb/WQSkRsfk0579A62DQZNJxaKgQTbPJlbF66wLlnL
yIk1toVozsjfegrWkDqfurOQHZnKsk52zFNXf6Q8HFsL7XP2UxSTLcyqT5lHfZVVIHfq9tkErctF
vs5aF3ayk1Cf4ag/MD8vgfo4SM1c3vJuQGh4asJIZ1NkeLlk7LxxCP51Osht1IErwwMuIuwOM7hl
9+dGj/ZI0/cKF/zW8XFY7uq+mmHll7Hp5Mc7kQ2YK+eOHTqn1pyT4dCLvV8KqnDOKWeBqjqvKUDS
1KH+ZZOXwd0bcEJZ+eyqkc0/6R64s8h2gk/HgNVwXh8/xSiPkCq0GftBiiEj3R2FTd6xYseNHbRe
H1vKrJxf0JqGV3I/zGXKoV14WmcRiKLzbxHMaGeC+rPDdJkPfX/ZQ4uMB530GW9kjO54V6InjLpF
eRbKzkxLjywJUtpeBsnIO6gJXHuC4jmbFw2ntxEDmajPIR6h4B+aACpJRdzR+EujhgNIY7/6Qgte
1KdE3NtN4hZLJx7r4kGce13tLHe4loMfT/4cv9hkh3omcGniqVJhRCW2/xVbNy5lY3Es57xLixxH
lcLl/0GEYnzFuSi0NOW1uoGWicEpmHdUNB9cx6O2i4QGfDloqNVVXTD+YQpxDHzT9t6M0js9VM19
UxlQV6qaCPWnb2R4Prpzq1l22JIzV6QlbvZrxCS5mU1jlWJFH15GJ0MQ0XlzMaOY7q7Py3w+RMGZ
WkVRrWhFS3GM9uT/RLUXGaVcyPXFKODE1xD1lJCrIfmotQC5N+pXwY4W53onNYDPgNUE1lG4DIQ+
fYXhRpGzTkGGeGW/YEQ9NFey85mrpfTMU+uI1x3TcbqUgV2yYUOlwg1+WZ/VnmIzamjO7zodcyXo
9u2Wb+5LF+QxxDSMN/iisMYtsIjHs1+BiAYxMp0fDzyYufrotgakgfsmcUnrhE8/MPyCxFdyLiLw
yAOFMoKPbju3JTwt1sYvwEmYAENv2ceZjtqqMzeQrFLOp02i5oq9EGkkPLMpQd+f3CCELyGThHWm
GPuc0HhxY+QolfZ37aHJ0JToLWtvSln2wC8d7E2yT8s1E9qqzP3CX+AfGVQbhOee5UA1W7/l+dc4
J19OJwfa1LSizwg1NqNBF2O/j1JLnfzApWLH1owSsp/V10zaXWfrU8KDu7Dt/xPhAFipGVhUDgNg
vOOurjPclSONzb9K92NQiJ5NvLcnONtHuT6LLeq3i8RSPJ5HXwQtyqJlkx7N1Fla1/k4RhuEb+kz
r5yeatPIM5VEBbLEjuZs5/hV9cV9/LlXQiA0KhjoqOEQfpFUdkt0Ch5CbW7PeaN6xAE/zZEcv72w
3QQjGXGPqoVqTnDkagqNG5CuW4wvrweTL8Y6G7m0SsvGD68bU1AAyU1QW8F8MRMUIYc+Q8ZAd317
O7K/8H0z7qel5+I1AIu5V9zdBb9xUeFtui7vcW7KfTWxWg/GZIKovr/6wtiTy4kXxCfwasOeSSmT
jsAmT1voVu6DxzDaTNljPBhNZlUHpF3eOQCq0cCDcaNUdyJBjD5XZnF64jcLMvijOIFwKB8N7SFK
jyN0ftn72x7ipnhd5x3ZGqTBOJmQ2ltbTp9ljriOdwGKvO8JzNxtg0rxdzwBf8lufiF05okZOVkK
qzETSFDNrlAoh6ElOjqY6uNmnOXhkyqp/d8R+7wVUQ9Y+I3TgTKBEhKqOitp02uTpXuWKKK3WKK3
C008OgHGkOB4iC1qqki+WRhI2d5Hhk787fF3LlVd5kMnazATaoqBei4mLZ+FT5fKxXf/mU5wTc0B
0mQYNlp0ArxqZLS+Vd5NXsodkKrm9Quh9Kq84o2PYfbUhlwmbuLTDg1cANwa9Qt7GEFyuJi9ZAon
Vh/t2c64avBJrgrX2ovOFWWvpP+r8BEKWPwyo7JPA7O6Bq0zKzS0SYiHTqQytuSh9IwOqVBGIVg8
ypWG8/B9e3drqXaLjB8ghjQnLF/CmxA0/0hhf2DuJERSJGqqZM+ju8zqnNfl09Qmhrpxh9YoWGqa
FICAC2iY4B2kcYxJ1gWaMcenoUVEcE15rf1ZUDqB1EuI1cjNu43b0hS820uIXhGvsDh4U5uMt58W
YLlN1Azvn/Neqjb9xF0wYES4Ut/KkxRBx3hVW2ejTGaC6qiHOiMRAtAg/+z52gSwyn1l1dInC+W8
60gtgrzQkjqfaSoqhLrCXUGh97cTNdrKR3gZBVGD6zqspwADoSHvTqtqvsDS3ZVJSPTIfxkH/xI+
VVccqHFnfHXCCd2l/h4zOrtXwBo/PrN9Lvib17emjFt6WN/Vr4IECriiqH6pycE7CkySyOfrRS99
Mse71Jz2C7N8b7vLPaZCv2UaZCCq7C0bT/X//ZIfLoTUbq1Wp4dvLno4iYVixQNOR+GERCfnILB9
vMkY5zaPHv9WfUcodwIIVnx+zm7i131O83/c0flN3poox2/U5ZU/ZfRl5/uwKDbKN8HfdRixrpk/
QMsAOTIIiag0yiNHnZLaF35UCgif+50rQTkxWMoRNQWTuwjtU7vcsnzRh8PjB/+j8PUHfo6miseq
Qm2OqmF85ONokX41LutgNz3QqxS6y2HBU9Oflm8i59H1F79LYjrvbyntYHESpDIJUKnT+AxNjdiV
Y52EQEqhHHgyj/fv2Us80sxheu4QUlQUwchKKDNCgHN52L9MUklxO/+0fwTLh3MnUf5b2X6to/E3
54PmOhdI3MH+AUinxZrHjm0cjtPmYAc0xNECCHgPi/2Z6cai6sJyFyQ+KGf1QIRw9i2NxKbRdZuk
+mlnOqwukamB4K1Dfv5JjO6YfnAoWSV1DaOrpuN+1yaBw85Jlrv1AU3yS5EIvQyngsn5Us/t5DtI
AAD2mrWLcGTolbvDRla13z180gj6YedL/q1GLuj8Nj141XBzHsY8AynSVZtZ3mhcbvqGYT4V+rkg
ZyJgSmn5O1Y8FiexfSx2QjLrdltDVGGiCnngY9MnjhgSOrtFoCHVhqdEQklBdcyyMgoQAmFUguHj
YecA38jqQaxEGCfBagMv/idfAWN2v062AMND4AAuuiIc4oCKA55hK+pZZLAPuPwV7xAU08qc+XSj
Bvtj/8Gg4dF4q56PfBVNUdCf4NCtBTuOOvIKlk5WOJ1S2ZAoF0h7iCBtkrPrQ21ooi9m9GB0sdg0
/ltYzqF3UyM0imd2sUUyoVdd8JnxZbgwxwawn6wbf20lYVdbUf3pIUPXUA//QSl3YSrO2yfo2zGE
40neFZ+TjHEeyEAL+8iysWweIcujtFSoWNtAldV6pzQSxq1aYJIDHlWGSl1gDqpmUgh057WOGOvv
SVfBvjidqj9LWSGb7m/FGliZ821iitq0HorTsRGRlUhUl09+mpwiYHjqi7C3YviIDzZaFKnZtR6P
7VPSIboje5KzrTnFDgxeeSVsMdNNBOOEwUU9nh51kt/LX2QvjABJjkwGPFo/Y+hUkQF0MIRIqJFk
QwItJPDAKkzb71kcU6+uOFh2zta/K+01NrXaCZziUeq4nMTdM6Q835ET19iGO7SOFGLDEZNDRxS1
3BSokD6IHgsCGklVPh/50EpJlNMEOu1NbHXdsG5v+qXoZ5ytL/U8OcodsYepvllhOD+J5N+PDNqu
rBktNb6Ajdi8/N3FNomtfYwerczJUSGGytQ1b9Q5AKEv48+LtRjCO/r8WdukcTvvwUw/p7LKj/F5
FttYUCPIQxSVL6V46oekyN3w8Rhoh9Uwv0twDGxPqXajuBBevx1W6gjUzgq+Crvg0Yhp/oPvtEr5
thpe/5D7HY1LxDyk9wGVkTtKIXEfiqEp7SBRMnywvJo5DFiZpVatZF7Lv6qSeGWuQ7VxzRdtvPrh
3jQAUKTzRP2tlSmJUf89SDQ5B64s00Dgh0GnSbUvvyIamRnIPV9jziZX57uNUkmaNunwxG2Oj4C/
TwanE6IhuBU6e55CB+QhSP0G7hK072dlV9cpPWeEJdPgq2JqqBo2nk1mPILgt6Y+77+ZfsZL9yVM
B85gJguSyCYG++CCrzWQ3XwoPsGwjPWECQnEkMXvFV3xKWBjJA3lhyYtDIEKpmirSKBu4+uZhiCC
k6qGkmccorOEr74mHtqlJIgdKwEnOBmjioaOgPugriO0t9Iusyey1dMUgtbIQcIcsCdY7qbrShKG
DFj0Eb/h4dtrPOQzeUJFWJafANEiyr9+vRqggcRHZaEYLIHLbKcteA0eq4SvIT+5yWuPXUKnZSvH
b1VZVqCodjShUNLtuD+8hMRth8mApJrjGLjrm3A9brxZBaMDvHwS4M1G8E+Qc1w6rtIshjF9E+AR
ad59VD/4J9L9FqLbqRoOuzntb5e7N2UVzsX8lxMNeWUiV6TMTlsFBeUtyzyo6U7Z7RmT1Nr8OVgg
Ywhd0VYK/0F1HJz8GYW2x5cu2EwYdtTwEa/LO7Hc2LK1gdrkdpWWTJyGlmmLwA1LzazNTvqK7KM9
25q0XQdBeCEaF945rvKHABGDX8RbOFJRGFk+Re0KpVEEZLjt7WLMcMec5fyFci2TAixu+oC+0eaV
J4MhVJFe6f5MOkH3slw+9zbNnfdOeP177LaPXc0I/UlxhL40lk5ojzADdqQ+j8p+aqlcWL+4MZpA
sDC9wfA8rZgbvJJOWERcwGYKuTGyaAKer5ufV+KfgyYsKoPuSG/raLusJuGeTPoAezz5xR78Gy+v
SpcQBgzizcxkFOUPm5V+QDnttz6/QWgsjxBQIBKr/BAPRX4lQR/YKeJXy3yfxqrAlDu7mgJHY44J
QLC0owk5GYOtwKsggxgHIY7dVT4M8lG/w3VdI6qvRoAt242vC6FJeLJmvZij7gvGtoI0V+2dbhn3
6r8Eu/ZCIy6ofLXFWbNvxH6uwhi/cXnW6CmSSeO/qCzhbKPNAfHdxUGkK+8mKlXVNEYWmTxgj0AG
BtdX7KsSo6IRGEDY7RvYTm0PSOMfW9o12KdX9Chy9skfwCqdTaH/OVLqmyBOB08Mb8G7qguCW0AD
3vqkjm7wIoWHsWGwet6U069nOsgoTjNLPJdjpPD+Hjxjxq8ukwY5XAAw5jJ1oCQ3AzvW2eJtNJPU
EnfQH7+/sSvHq44+CpdCR3h10j5uLrRrIpQcPFd2vbMgCVK/pgkA8DSr7fTJG/BL8/TmL7Jop6cX
r8dUpEND40RjPIQQmCzD3ngcx1fd9PBObeKhEauKVfKQbIwTZPHOR6KV4o2/ORCaTGFJBDacwTuS
9BumEUl7VEOMuOECsmbK+3+EsrwdmzXZpzAehe9D9mb1i+Yk+t6ryAwDPLlv0cY+yUq6U/m23zoA
+WA+6d0hJe8JVyx6Gd2DEM5dwksmw0iYHmXX7y2UupU/pfOfneWvwFgkl7kwn+dF18GKP/U9oMtR
wNjZZ3nz2B5MNCIQMof00/dx8yeWLHoH3o2emPsnlFICcTEeq1BZGeppBVz2IjRDh4rMQBDbag/M
Rb3orV0N+Ny2vU14/MOhzMkxBklOmJRiAk+DxGWlFXLTWXx/U/ALIkXNj/tnuAuZR3Y506JsDOfq
rVAFRdt87Royb3JPt9YruHtNY9UonQwBIPYD9jmRDA8SuhRYu+Jb+2TO9LgZn6obpju4q2YUQfYX
x/TNEhNMuZI+IuMQH4r6ZjzvaeRJapLIDccUgpQ9WGFTqdYuI8zI58tt0gciIJmJjMtfipokDxcO
ZeR8waO9Iw2YsC3FHB5+jOjIXQZNIGpFby3TedwJjoPbpWwdiSqEwPzL9UqDzpZiuBsJS6eTmViK
vpGy2/mfN1KPCYkgXkre5s4vkvrtnWKDykj5hm3P/oH+KaDVS77CGrObs7rdWHsBWiE4cNykdOf2
6U8H+wWP/V6t7MTIhFa3eBw+lh5WyhaRRiuLUc2UgZzSbnqbeebhLsAW2ToYU3BVRoSH3F0qHelI
UF/KJDEc5RP7JWSCNMstLoc7U5ijoUMxarHEyvWT81hmFyzlpiRnHrKdogGOazTkYQpvohtyaO3o
M2DAdyPp+01wQdKBoSkn3hjdSpUhW9ua1sPNA52K7OIKBDBFThZS/nK4H5NE/JjRzaVI8SH486Sl
gPHHBkTkph7cFjM51+723ECAuUib/du3qCn09vDkTii0Ymf5P9uYiUD651CvfVfOO//TQi94w/sw
16pdJRwz2ch8W3jtnXQl9I9usnv0EATKKTO4ALTetbHV4UfOwtXdlXzC7/L2jpSU9/AbZ6LcMWIl
OgyifNaxJIKEEjg1pm8SshSuQX175BMpM77Ly+A/r4GKInpm2gyQaHOKM47IWwqX1dWLokOuhFTN
9d7fOknC/hr3dgTszZhYAfmzbNF9r2HY04bS11vS6LZ1QgrgdkcEcufH9cL8Na3s3mIsRS9VUya0
ZuP3qwYHQ8bX9Ir3mdwZECN8yKHHcOteAOQcNybyg8kAg+i6BjuoraDZeGpswvluDDqdsTrQ3bAJ
rbkiwFWfIDK25IAkJpAQOHhLy8YuFkWhQXDmKjR0WGscGDIO3AxXNUzT9+fE53fqmqitu0EmRBnD
Fyuc9zIeudLRBmZ7IUhMRwv4jKk2dbtbm/x6wZSwJqLOb/U8AmjBJq90Z25pXSCMyJAYF4GTi5do
dC1IovbruSCwOsXWcoiMrOUNRYIc52YarwARmjCL4Iwray6xVdiAwX8OCLUQAbx38ymO+KxHunkz
91LaK+YuHwjV/uIZgkgO/6pThRGhf7xUZ3CBjEQIqpdkV3babevW6hTd+3tJlTIRZSQYxIXturrp
b+D9gZ7htcpmtIecdzrvgrSyIJSNmQGUXjIeknbdPpXR6H+mTXeiCDWKrDa8P4jqETTAv4f8m57t
ot96dkxMWlhMX3HLKQ3bliWs3aOANKH1R1NJqDjisQXj9Rc8aJBjyVIrNqlFJt0xrOJzT9yQnM/+
1/iSDUYCdDPtUUwQ9uSQTnNELA/TATbs1E+vggnNLRWtgmYuDxE2/w3pNno1pp7XEsXpH0ilX/8v
cRqD8nS1FMYmKPp/0cOp0r2dsanLkEff8zEy5AYxfROHU3i/1KYDCicvpJqMhtCjfqGdqAt7NKHO
/UJwlm2abQ1emSOG29FCOCv+G1RjPXj6yb9EMQwf4+pmdpq3gbnQXLFgigXTBEFiEJapJNfjOuKu
ST51KIbhXzwKwWLv8uK+QVBDj9cJOa+3DUo7IH71VG1LBgkT3SayHeHW7eTBZ44H3dYEraS3Df8i
QLUtcVd5WGLX6YKrQ4NTd+i2Up0RdbN/3sWcHsxfReScqZ8RGL4kVU078iu592vwksBlHwAQEiwl
hRN6zw6wFgmKAKNTAKuUhZDwU7G6iLKqQrGC+igZaz2pBl3505zj4aoOJj+lNw8C1GAS0ccr1kot
ZUPlv+ZwL/iYhe3zssbKgWIMkcHiPj60Tg1k7xpwdcXj6O+4jBxMUpzcqahkAD0PM7T8EYHKF/3N
asRhcgUv1Sbdols99Fdm+CVj7h8itAcTi0EHP2uKl01IHhDz7NB1RKWuY8x1qTuZvcJ03Z+150ju
2L7aK4zlcCjALxUPIj5YEkto5gUW49WfwNCFCAFBwr+fZJBe9GcrfUjnZfkPiXTztfVYBPGbIxKR
7hwGBpXuhURbCpDkbUaAdwyBCiyUMVkVT4oKTzUxE1kSOfRWXxiOJiPwe7Qfl+0KzrIGpKIEhMgI
onmTJYPqDYvt1n7B/3OBWqjcfyVsngSDjMjAxID2kkz9K7Oau39BfehSGLEkYyNN8nnP+ttvXVfu
Y3xlzu/Gplaecd3Vl5A+Cogf7rF8aLvFmG/5rK8nW5gTIkxWUkNwtZ+yofrJ4fMi9tHM4EpqPpAD
RPH9KuKFZZzy24vftbmOUmoKQFFmRi0vpAxFxDH9Z62lVQdQ4TdLEhIlbaHUWqVG0g/hRlM71D1e
S/Na2ox8gLkDyKlaiZoH6731LMFrKc2KIKfTOhK4Rvi7Ulz1RluvnTMNEALXUTpgbi6oW8GQkHKT
rD0EZ+yfLbf0GbUfrtAIT2yfaqCREPS0H9FiA84aGxHPQ2JuJbKMF+gEF7yP9ELQYPjqjmZd6ps7
GQoBaC1v3pThhWw55D+rbkXU+DX7yBdBcMTg/RVU3WWdlO/vG6Ughal0WUPR9Rqa0Eil74MwCeyg
/StspsTkhGgEbHkCgHGCaqoCsOOlKDJV3KUMHOsEEr7kBb03nvygWlXVf1Eq9KPvXEP+OZPgnxp5
Rj9iYyka8/lLA58MTpqXKX2NWZUd2ZN15cEFK0Tu1fBdwmy5VMjgnsndGkhhwXFXk0hnJyvNo1GX
WwoscYIxKD38zR935yMNNqI0jED2vdZlb5dR1qjpZq+laTXGtXi2KRzQz07ik27hoqYS2TZ/0tL8
1RGW7lraaxFiiSnvqhnj5fZzrDvxzZIWI0YAkjgCzEKjJg/cezz+ZiCM+yuRObWJYPixTkiw0s1O
q26NMgZu1NxLSwRm5qBHb1fpW7XfledyKj+pB4hdm8yMuUiOWlBRkOsNnKnGomTTGkDyDylFu1Kf
CMywJdCYDW5mRS3v9/glglNaZtbacFp9SX1VqOmEgdZM+OtoR+Co9kP7GW8Pt8jXEEaTNt/puQ97
DZqKW6wJqyfSQ//TOz3pWanbC5XQLx3eYmO5wZf/pp4eXkckVw8zEdIpkD0cWl2UvcFuzTwO6T7/
jN5Gec+3ZDwwioM+whkrG/ey4B7j4HLTw611LsgCikIlCjgXkE3RpbUsu2o+5C49wFYcu87o9Zi/
51J34osovrEQp7KSKGAhpjZLCncB6GUIFbQhYWM0CKn2xAxXI9SWJ2Os91VEWXbO2TjxD/U2ipVn
nBeAlVNr1QhuusPvJz+3NPzAQWgeBH/UzBl4xwyLQbcuC4VU4jNHeI+c3O7RNvAl9PekyHR5FKR+
hDJFlb9MXq2+Bkg4bMZoqCn+9vs4ePqoIQqGnRv/Gber3K4N2piGX/miaEefGxvMtLxpL8euC9Ot
cKEspnMO3jw8aDzNbZjQcKzMxAYd+awkHadVTWdIOKf7T2xpgNnm//zaHjvquA6eoZCHwikB7f/e
RCndC9DCFnJotwb/4GTFv3n0w5oUXjMEiVTsIOiYUJONdWwpkCidxg0DmBCn7JYmbVFCILoOCNDq
m8X9QH20I3d3W6/Wh4vRdPaG5bmpQ7MvfaAbTJyyMU2CN9swuVIvNTZWeRX0cxce8tTi0Igwg/em
IgrkE+o0qbpGiTFyKELE3iww5jGIFdxILfBUKLvNm+3QGxVUQAmBW7zq82mBT+obdLJWYCOjATVW
Fn1seG8ryo1ezOg4yUjlCPxhJLcTQ5znycsF9A4avPzXAmXdlzvSgjTNDCRKQcLTwbP3gLPbGzuO
DiSSS2iZTqaXuN34IMSxNDfEiUnI9mqTPE2mGRyewF1FBpSc4lEupuS66aUBLPN17FaFG4TLbKNw
vG2gFH34wPcCH80dK1Xuc7WDvDwcMHELt5A8Da1xS2V2zhjLNlIRfDl2fzNvZ0daKAXNR0AQULiV
bX+zXZkeihfXbQqmEtCKWgaX/iYB2fpGt+DqOhs2Ub0UsxWQm1Rt1C27vtgX6SKEEaEnkxgJ4//5
beamiAgpE6yAw7e4yWCBw4sErVXQ3Tu+BzIDKgcou0/7IQPwZSa2QSpVDvLBhI+8sBl6ttM4mNGA
oSF652nQ07Q7frePNyEuOWAJyqHBTHdV6+0pTyb2VZYXSyQJhArlQO3xaSyVMBYfHq3WVtSUIv68
uXwDR5iLKh8TXeXHg0d9XDgGn3AZYTmUvcJGqNJcroX79MS+UEj9msjtmc1Q78GmzFhyna+FT4tV
ldHOowgB7Nl3dwq8sTp/jh5a0oTZkPUbScQbXEvr89E20JdEi5IrbUscN6jTyM3YhjtCNOpNgKk1
l9desKUpTPtGDnxvUO5pd7ApBG9WGBfOf4wbQGxvKA3mKdjzTQXTyxeKST75VOyBwYIFnsZbc0Ah
4w1n6geVajkEckoEJfEKXCoOcHs3JYj2W6EDiApwBx/yANEmjQtnC9+oUPvWkQ4+gW3JPV7MIKtK
NUw0yVP2B8NYCcqy6gtYpwCH4AP39L8ypN3R/zWfE6ePuGn3D6rocX/bzNsE+Fg31OoyvKCwvBMc
+2bv3JjOEOW4jYPanlt3yaQrK1s70GAFgKuim5nyDoosQQHj9YihpyWwNO80Hf/k2Lwl/aai2zXy
Hx6x7nlkO0cvzLqClKtrzWgr/uUG41FPXtdbbQpuDywkR3bYC11X0mqoc/BWisK6kIo+Al1gs5H/
iffq+vwd4kz+lCstsH/pl2TfUk22YOQYqsw8YwHu8dqbtAkIgVD5DEuINJ6Hy8Me8o40GpIQdAr4
s7QwFCmn8CYNllNmlpD6iM3L0/AzA0iPSpP/PEPkHqP3sdAJ/mcY5MROv5daSzbLVj+65g+r4EL1
dry5x3Mjus9adM4UXszda6GzxusfvHiFSoJH26lMQTKv69qzHtoT5uY2RdKIJ0egChDNFU0yYsZq
L5RZhWxmwFEj+pQwyEM56fMfCa2I6B4IuyjNbx+PpDBiwgVNwsvQaH+l+86BG5Eg8t/TwsbehdAi
U2AlLvTV5suOOVaZEKOX5A8yEPp2rxnMxJQBYkSPGZuf2K4/+oGwrlcVn/NXPySedaC5EU6LAq4E
aB8BzH5pbat6SL2tGUp56LM/oLnhMoz/Eu+qCt/3kT/dDRbJCovyPbmVVoa/Z9GU2QLf88W7yuA/
aE/mkYhlkAONeF1YLQXcoAN3KWiW29sXFC30OHvjkzZiOlkyO4yECWf5/jsmKoqgzpD+SeF0VvFN
GEEyFhlBPu13LsbE3FzPD3DWgw6IPoLxDT/GYNDHLpfNSPu+RisDsKr1Q7cHosnnlA2h8RFiMwIb
8+FZmTAfHBgDISTvvbOeDVD+7eRFxqio+fvtTIDapiT+3MtRe9gp0CUI6Xxhc6Zs6ZCap+/QpDKX
/lq/Eg4GzPzRcee4y0H3LyBpNrC7+tzRrelqQvNX8lPTAGEQ/xMKfRR6f8V+wD88foAjIvVMFa35
3Xy+zQSjoczPu8N4XIqpGxJ8CLwWhkFIGNBfZpO2ExB0/rB2YEUvcdVAfJ6L4C1GrEhtsndHHqkv
HO3KAv8sbr06N/eUzr4B6aAx6oBBEt7tDhfBHZFnScqUxn3I3GXpaB8auuO7OloXAVQzUn1B6C1T
6B9GH1IJiDa/0mFUfBx+hTKqBn8+MTiAx7e1NYv5kKAHJZ3guugkFeWvoZEsx5zHqGwouH1halwn
/GeJFGdMkd+6hXz/kNfnltANTtvMZVvXQuJYH3GpWjQPF62yx8qHBx/2Rb8DPJYJXt6RNDeX/gMH
2TVmFrhMbrRIY1KrkIWfFjvxdj5N5IsGt1WbDhLq4kMLaCnnHQX5Wxn5xTFE/ETgyP1pJ9Zv+aj/
kL05xlndZGnhzGV+2f9gDT2U8LGPOz/ASISDNzbBt2u7lcNapWCRT54qZL9zkf8b7A8MaPegBo58
y3a8f7mnHE/PGHc8wQG/WyDfuM3OImqQuYwtmx+J2/O80m72p9I8JVKrpy5RdVvEMWANCtwMTOMI
KhGmTVS3BLpmBGZrBnLe3XlGHXE03vWls1SOPxPVF8gEGB061GX88A3pHXRCNgp0kuPpwyu80oHW
rGcNWgi/zDdWv3wzLOrnBW+9kXDbrxgjmLeh/0y38BM71d2n7kRHSbgC5MqyZgBtVe1Tft1/y3n1
gQYq+iSmCelG/OL2A5SBzLfAEoOTSFK3z7eAIMNdUUsMXjWQZmyjo5QxsXQzMpj21EhbejbhjuHc
xL8iNkX+AQyA25+1JAB2c88t9QGD0zsh4SrAgnrmz4S77KRQPi8xF/1hK/d4KXidNWai12yir/fn
1dI5WU/rLbT1vblBLAn9pdwhGId+H5yFDUMuX2vBHKdtE2rLJepSD6z7cj/66vfkH5TprYpukYHA
Ba/1LLHfq9lLJ1mPxurqrczM6sBrrAiWcFQFW344qfea76eIoNBQ2A0K27V0l91rH95PQoTZoYUI
dqohPGpf+1RLo19VJd2Xv3YM/dlgjgX5G+fb3dVyeBEWMzhWkra8pXtXAdn1/Uq2VCYEipLII46K
BNmqoGIsMytIoIbi+IGd8iTjRfyNUp3P4IfdeAIad6Lu1IDGvd/lOPi7knkfr6X6cClqBSj/gKzX
KcyzOQWUP7z03JlmpNXA/Q3gqnEMCZQlN4f56X9h0AHNIutTf5JbcQJ+1MPPii4GBX5Sc2IFB7YT
lkxo3VQup64ycmshXq8Uni2jy2xr88y0tQ2wX4dkCVvc0nyF6tJj58xaHAnrbs8pKoWcfUCEBQNO
AwjW+JCIzfvzEgtQXNI8tB+khleZdnizKRY8gLucEdISwwu441nFZ+roMC0c4Gv1u1+L1XxUjKXs
VA7ljjAT6N7CkyLRiRzgjCBhLmYGCZ9qfpUhld7GCKr/3DE8N9kLQoB2aRQvBKt1riFUdtpspo3U
SLz5rRKPeQSDHGODcLtlbWr/BYjo/lWRe0i8kPiWCXrRvMWJG/j4wx/4WfUZS/xgU4mXMeX0evGP
02Pb0mmfux6GBcplSteE+9DBpLX3V3lZ/jzIq3y3JoDL0OfYf32R6qAtx/3gNJBV1AltHOaiGs/i
tymWXUPe+63K311/YLspGp/ggLIgUCZx//Fc15TuN0k04kusO363eFPdtDqxfc90Cj8b2Db1OsT3
GMgbBKeNL7XAExIk9H7f9oKyHsg1g92Xzn6BRjmdAvX8UdhBDO+yUYKQErUH3X9pH4WZjQvoRiJc
qmc8ozej3UWNlneGpHEgMinih4j+t4uAj6tmcdWs7lrBHU5BhJgGgi7i4ukogskSJfSnvrFM2iDM
jKvT+pJI6IUW3oKAbq91Xp0PyUlJ/jo+XXcdqJ6+x95ITYyvxmcCWEU5bjXeJN0vKcblGtIj0MAr
kbykiN46GAIIiPZebozxlZLavAyXDsTDN3nJ/0pBVx96l+zrG7+cNy4Xfk7tRbrg5T0wK+uCowaD
IDMcGcXgF+b1mltG7EecfNMi/EEJ6WCcdupAVAIfxh41dqkmHDevDWD5EA4o+7pDn13I8FNtLmWV
u87aJrua1lqXN3xedOh3gs/+6g9TfkJqhhw1GunDPBH7qOqFNb80qfbUbgxbT/hNrZOryp4tehOV
uQnmGNrzkhYsakxAHhdBVXbQeQxQfsvqeSqLeucUx0v3cNUiZjhafHNU6HUEZ9ROyNWnFOKoR2Yd
fI7rRCnur4rgASUN6W7U1vdfhUZA0oAOaTtmTwns1B0MaA6nrPfzZp2fDHaO9WOJE7zvyWskSEP2
9m2icfEaBKOXwkyVtz/RM/Zm4t+dr1bp3s5EW312LboMYa69x/3Mad0jyNZTafD5HsYaAhOWKjdY
xURfcWix1oODmzTdzjb3f1cQR4RaZmG7ucBgkLZMw7GfVusU9mvaVcME2y7g1p/Rx/d2ref2FzoK
jDePqmax921qmIyF5Dr0jKm0piW/nBByIuClidNahCQUu4vMT3uc1S6l4oKCVLU3vsYFuf0DrPr3
2HFer+df+Z6RzJd8HdORgLEGMebsA7ZktJLV2s0+vRt2VjIGl1uABG0W5atsj2S+P8ThQOcLOGEe
laBhG9tS1kG4yI+jUbPRCqBwOIcYJGuUuj7tmm5OuciYLxW2n64QtsXxhkNB+kruUOqzwlwriBqs
N7ngtNtv4XWl9i7ANboawSXyIzpUMNMXI83jHWOT6+UtzIG4WoMlpUY9AN0mtc2TLbkC6V4G77az
nxDAFI9IKCTM4nv3U8bih6mLG2jbqHj6oCHX8ANWkF4geN0iBe83q3Np8d2XEVC0N4fjP9/Czr/Y
ARCkeYjO0y/Bv9oMXoI1VnFKsN5wifLLkfBDeW0b05h97a5MdGLpIvRWfQY23Zf6BmY5tzGKpruj
VKm4WtB/BGvXa8lkg89qFTTk6SXu+v22dg/WfSTaBX591wFHpUh9/XApBXXxtZ/BDo325GI3WoPr
B/SMhh6e6dKTf9qR3gZ8oZebkJK6gZQHsQHAVlegCVz46/AAIiji5klrXfIQxZrgrqzUraD+ZAYg
PLHaNZiPU6sJocQHjrn0J0eKycaVfknctQ/2+2SH6mZ46qtRX3Gdctb0frJia1sRvnMx8qGyi3zE
DsCNpbubo4hwnaN5lNhkCHDOWu6QwHufopeKBw48HD9sC197nFSZZrID16XZmVnVFnch8ASM7OQy
POGT7a8lTtA6/OTxdTAhJjS6R7MKgafqo0uMTbczK7t2P7amBGZaZBr+hjiF5GIKWbCLMlmsf1L6
2zj1iFL2fJvLlqXc3SJATWIPuRMezjsyc6aVyGPNK9eTo74HQoWvA0NemE2/K/Xw2uGcZy6VpQ04
VoAqfdQ5/MXdZLYuOJn4eRXspT+Q0kF2EzhmKB5dsqOBLcYd1KUWb/IB1ijfxfdGtxUBHrHeRwV8
CMPMVMpSr48DQL4TTc1210EOupr35UpngqrzGmHBODFFbVL6aOJwrGQc3XE+upyxiBdIwLMS53+o
clQc2GHv1pgzOnWJ7+EhMZ1727E4hf3+eWJQ3SeLCGePfixZ09GFy29rMGhcJ7bauqmBtguthajz
JZDOJaFXYX/PMqXkfQcaiTwJKAZhjwLTp8lYhe0fRNEWOVEARVyUjkDXunyHqNGW2mb64PWHJWOC
AjZnLyUwexhD9EPUPC5JbCk60TGQ7uKgWvqEBcMTV61LFTZcYu/oRw2bMTjdKdxFxtgx6qAbCFbf
RJ0OsbCW4jPtUEGXsp0ap3LuvhLmTFGOR9KDPMAwdZHF60DPbqdBQVJqO1m3+vDJZSNSsPb99nRm
loJRKPZ6k9yx8GQzUQBIhIYOxhwBjIQfiXd+xRmN6ZPdXMeXLwH6lOatqMYrQ3nBSEaa4SKouTAE
Q2G0BKyBKJ0IlbDw6O7/QOg/V5lkLR65nEQxpkhy2lU4z5t5rhvEIgmKAi913W4l7fVK/Aq03kAd
eiBYgEG/Rn45qP5gH+pWMhxqIs9eTH0hWQAxkevp2ZkUxhOsUHbZzVFPdkUBwBx5Rf+jdb4WZR4W
wlREDnanuT3bNn+JVNbUDMQR725Cc5FUYvwtluof2uKj4CvjFv9h58voDp/O2QUvB3JDXkHrLRXT
1yJV1+aiUZsL1WuxRfLOxaaVmLx+S+AFkChFGhDWaCE0Fi6DEj9LcLADm8sErOumFihAFeiIEAuJ
TBu+37tK+sj2kw3y9JNB+S2N+JzoR6CJiJnj3h3zcF7GCe4Tk/Jld7NVAWXP3cw+cqrM3liXUXuS
13lbeeLg5IJQLzAiI+KswjWCEzTtOZPkWEwgE0SRIOOgVjgi3811iYZP3YRvjVNfH5JeciwWQrwF
KsgzFsETzNBNqK+hZDI2mRUW2yUSpDdhQFXrx/it9Wrbck9Bj15vr5TWxHtCAjGP4R47wGML9DY8
wZABTMXQfXAVMyPxAmY2C/MvkNeSKFAfBmNjdP1ihiOJNQEgNCPTOZM9XGespsBptyPHdAB19fPn
SrSiOjHnvTquL1t+weG8uFqZxqQMX6mBhXYic+Mq2p1QdGuNAmEdsbff0nkkGv+sFwNDntOzvZnK
dNIgFs42ykjudB7xElEbDIL2kLaAUDIpAKQdJNfEmINNRzvnfN9L6QrqGZt4S/Ek4YYeKd7lEi5e
4/Gjw+MhH1ecvIcu/wzsfbRbWBdTM4U1Ej/2iyRowTTND1E0emo2bjEgOCeIHNMkBxg7/hbaVT3K
JiF4z2S6oyzI9oIiudTFCj0RGuLxXtGnltnzyeUeeE9C0gnWCePMTA1Rma/AH5tmt+w8KEhERWIz
KVvFE887W1b9wGXFv7t74yZvH2YjsZvCmCEk7SQ+/5du5gh0TNTL9x1f49rLcDN6coQdP15137fF
SItFdecZiUAsxmFHrKolFcuxGKoHDpyc+goEKz4ly3Fs6UPFHWha9NRwd4XtQEG0kjfiCxt/JAFd
VsAWwaBPWUTG4SkvndKhaXY+YX6R7rqfDS/qismNyuuqepAfmyyu/PwJi6zeTR7Ws3QgiARfShzE
3xmclVNB3xjAkq1706UgQIOSuGpawcv/7kq30BY4kD99yaL+mimjZW9x/svEn9lV//OGtTJmjk4j
Ctst9AZGaPYSJwNLfIsPf09xRM5B8tE/z1dtMVikwyd+trEj3HrvSgPt1LBbiJzu4HSQv93UL//J
z+s1O5E3QB9K87ELZhDnCUv+u0iWcXeOe+njmwSM0QzksG1FD+0WzseVlUUfBUdTNcV9fo/dtEsf
Xiu+MNCHzpsUc6ZIz5ZY5rin9ncA8XzoDb1TQd5kEjqSEezv/8RXRBsPLf2Byuic42DngBcMm4RH
B/s3FeJKSbkmsXJRsyjraWfXqdwHKZ/jofcLAHfPphZkk8vpVtcvWghlMqL5FVqs6BeIeag6F8WY
gUZaYDBvKDkeUqYM8RoVsPOyZRSgcv3uTXKh0NhLFygF0cKtmRYztg5eli73XDB688sDc9NTAOyn
O9LwBwUBViocCl6rlTnQ8mx6Nhgl8I1acDz76yN0Xp/coCB4Z1HeMpdzKWMISIp9aHXKmrO8BuI1
oN8jn/VLzUWCy/wrSll7mHlbVsW8r57S2CcUQoYsuMGauKF6p7GcrtdZUq2ZTNyDePXz4dEdqc1f
+waMzKmzkfM+5bEE6DbLthh7cx+hOdkRHfWsO5LjhJGsJyHJpMu0khBgRMBlumMHjURm8AZf0Lic
x0xEGJ4yPs6IwSbzPLO6tuOZT2FR/OKYebOS3fZCQPPsCWsUGZ6bFKkaLZJtR1x6IbTRgKavL/e+
CZyShAEte1kZzoiaSvetrHJ/jaFT+Tz7bIUZg2bhhRusO+F2sPyL48MoL0cS4pci7oMLSRzDxgGN
PJktYVLbYBlqNvDOmCSB8sSOgYE7GbBubqUwhouzXHKIKxc/aGMaRyx43cfaAM/7m9AWnSfMXEXj
Qa+HhNPqiAAft5sL+cZVAhVzFPvDM1XlCq3xuBQU4wU6/hX0UEY046Ha9sFs5fjp85Z6UeWM0RlE
5LI77JokpbaTnqPLqKHfWMAPuE3MCNP4NTdjlUpoNfCa3KFyXI5SIju5/GpdniJGm3UOj9+hdIOH
aNFLbFimwkmJUvCVuFl3jMHdHWAoVm+/hXcXtXYfdevE4C4qoDCVYKZFikXi8SKvDuRE7PsYCGfW
oV31e/QEFA8ILjKFe7lh86zatuRdTgJBHuijgSNnen7qa1ox6OxiYjfFt89kcugx1eIZpHeSt6NH
eku/ZFGmSXImBZ7weTgjHLR+yh87KrcCiPOsj1pHYGCnwbME5kcxsA2iNhM+acoKlxWmv8DaEP2E
PleLuY2r9etcLJN7r23MRTt0oXF+4xrGhhwmvVlSh6i5S33nkAeKRvTkRNAQ+qJ0HBUYTqHK2FAA
bKttjzZRLMXubAQfmyOAp1PeicoARRoCAIAP9tYfdhthO95FHmUOlJit5rJwmr2BNUZ5j4zD9d8U
6m6NcM//Fr2OKn0QwCWvbT5iQAz/D+e0m9dgOL9TBS8JuhIRl10PPAOBYJycPFGdzgpzs+YIklII
D2rBVgZlhvbYDIaL4lDFTZmFrZvzT6y0FZiud7aOhXfk7wVD/u9rM6iYIUPmRoGSfH0sdjuP9VkF
xPKK4NUQNaCuNa3Ps97HM2xjJi9Yn3I/h93wOiXDSYMlZKHnSVnId5Kqu0ZPj8H/2yJgQl6I+fXU
CrENkkCndTMBg95n5SEg6jHTV9S7kV9hKvFFmpyZ3Iu39fPLZllwdsEJsfNj7XpkxHCMzhBEVgr5
bwOVGAhPBopEQYJRCAhaaJT9xLJOvmJzmgr20eeAEaV8Dj2SfAHiUXYwfZnnT/CpUZ/Xp40F2Q0/
QLc8iGRNeMEsiM+rJ6qWhpK2tc5FxrrN/9PtH6+IL7Zp98dZYpBjlwHO1JxNZSi9WMFgAh8CcsQx
BjMbV1pwZYqEmlcGg4jd7ytC0CCxh9LLwqHWK4VLWFx6EMFkn4YdP+HGfu18koqx2MDmyiRwyhl2
a/RI+fE0MFYVbkPXRUHkqymEou/JSj6A3HD+uO6yaK0J8SslZJwpZZWEtul5Cd1gAvBKxwdugmqh
aRMmV91JXcgeRwVVYiidBJVYIGCrAsTmYLcD2amDnnEmyQQoKL01Me0x0ItVhaztOXVvNI7zPtuR
8lbS0wRj44oZhaOvk+05YvN9H5CEX1lYvkaQlLoZKJuklzyBDYWkeOAOmJBiDkZyjxGClVBrOXIe
18kKepUpgXSH6gFF0Fvj7VJmyI3fJv5wEIrly/msMO/pRjxAG3f5J5483upLnWY09xTpbbSXB+Bm
6Mna86RcLVa9luaAQ2lF85+B5uRXpE3LzjTJc09/QOhH2rOezWJoHYuiE/VEUaApu1fsAUnooqJ9
QxV3uCpm5abCz8OSuSXqmzAxdruKygMOYjr+lD/b2D70qVD8dDETHuT7M6lRJFNpP8HNZaDnEy5x
00jJ0rveohskUb3ETK8pBGuYyXbzeZrrq0T/0Z7t3zslf1VKJMTacmfso34CbSNd/7JFKf5RZMWP
e/9Eu40ws3rhwNH+2AABtDGjRzkaEcVCGWJlHPUqkaFg17lV89GJKkpyTUCCaXpA8HROvnGcSPx9
ZkCCJ1USLHHbStpBrqDor2NrOg9/jJURyGswayKr59z7z3OeKaX2/9iNUcs6ZdNa0i0BXyR4f1O6
kN3ReWiHZCRG2j48O2gF74e7DMqWaj+V/oKyyW6u8EwDjOQ2mxVP8brbv3rOQCqlnh31UUWcybI8
ITVb7Uf2dzk0mNx1zLQGFnKGMnhraKN5rZCCM57b/VKoQslOcvY7pS8kbJf6b09S1C7NDO7ipRQl
wnLheTfafkQ4ZN250kK2gYBF9HVoR7P+GToGj0kRkYxcwJBjbeiH2OrMrrNEeDgceouOZeB4uE/+
zHAuWYtm6p+U76xRLpGJ8FSV3byBjred+dWUcYKRHeJMBPHcEtW5SVuFoQd4BqcoOvGTUX44fsrH
QvrF1VEfdeBloC+T2CWXzO+DEpFGTRlkg2b+nYzfdhOsSDRlj0S4keb/Kkjg0K1GRHwOQnkRgd9w
4GFR0ChUrtwkafza3tAZINHX684o2BS9P0l366AQtU5jOMx8R0zSnXsNMX8olXsmHgfFSAd4lpDH
jPhkPr/pu5S/4fPwREQ9SeNmNCNXY7odxex0YhH+SQu2duW4ck3h2Qvo8fA6U7rVLw8G1Ph8wOX8
YxkERByO9TH0mu5phavNOLAg30026kTS54XsTGyr57MtrK4MOaOMVKfCtKIEjuqAi/iRlCrbNSw9
Fp20W6qILQ/5QVJwO4L+xkBGn+JbWb7waSG0G5pToJtTJNupY6w7m8LYs7CnSWznmDZou8D57oo3
nSuxZpiqtYW/pxVTnifrBvphUqK1VL1wseInv75YZViMHOSk1JjcphPCKdolTpLXsmMRemuQJV5V
nA7KtBP+TwSitWyGaScs8EcxLTHKh+ZrspdmEBKrw3S90hPgGf/1BvU2CzmtfIg5YdBoExWp/Qtk
rytz0dqCRoOx3KDQ0LL7sOv245Yc+LhE0ZI60tYbiYDEQsObiUzoZ8NndoCGv7f+bEUVtxMGUT2v
U8JqGgOoYHyBdmyB4zRC63HbOeAUikjLkbPmm54l+P9eNQ7QNtUrT1cVQbdQ95108ZzGzRpKQMA1
K1HmhWOiW0VsrNopocjf9drdhaQg6AmcbTPyaxlHFAKwymX9Gw82zF1Y9AQzCETnKAsO0sUz8BS4
CZFBttvztibDIvdArTk7Dk2IgYkAaliAgON6EcDlZIISGvgyY71JCm1D6J7EqGygemlXYcLK0Cbk
L5dZtL/qNJrmFEren/lqynCi/h7+Sp/yIb1X1XdKjz0b2yUStz2ay81SVNCbLxpNO0ASwu+YJ9N5
E/knpgcHYjXFMDh9jiNUtkKU0DUch+Ls6iBHUHpfXDgJs0pBOjtXoBtF3Vfbl10kv8GmGLmH9M+Y
f8RBEQMoOK9/DH3dSFvyoMLsUUFMiPlujdeF1Tp0P5W5uUsb5p2MIN/abHwlffYWh0ka2NWOhlkY
KAiNEt8zvYbG5WCKHeoPTWWAma2yuz7+ZL6JP+lcDB1zG/44prCi//0rD5xtF4RyXOXDmCwLl20u
oNs9STTTRGeFrCf10eCc+Sg6iNgQUj248YNg/pMOoK7zR3t7uQtgt6ziIfQpI2zMrBg2FmY6aXnf
FWVxDIbCV5GcfG3lxSH8rQZeKAyyxhggGgDre2JdL0zucJjr2R1/uJuso6HzGC/EpK6SNik26UI/
DXtMYd/tBidzrll7BMID2dj5hfvwVMVJYZULqUK2IEMbCakLjvAuG85x2/T3cqg3TOWWE6DIQrrQ
MMxcuC1Oc9YlUZoJDyfRJXQx69z1Yvfs1WsOkkpc4dMnrwq85JEr7rDmUklRG9UdWHPaUqc2dJTV
JEHIaOPbrwd5Hu99EDGfm1XhuByT74EU1nMOYg27NoDbYwUlADwvuLL8NcIWMnxzCTdV1z9pqfEt
PD1wUzVfLiVkFHEoHXlIcNOUpS/CBo8/9WJS7C2VauPjFEYeFri2CyNjQYLnXer8CUJme47HtUFI
t8xvP6m7QWVyEtGOatqZYv41tXx7eoL6Bu5J5clc4WVpLW8ZNaVJPoB3AV2+qe/Nn6IQC3moEq0Y
xHPp+UmY6jzvdoq6opYWLcOrVJED0EnjAODbJIz5Xffan6lVkDkAUmGBlRG3ggtRWNHIU4YDL5vp
+jXmeqlKZvW9ORTigo/KwCYWIvTo7++KSyONOvirYSkwTIRsI1HaO/0Q/WlWvcRA5eYXwePCFsrm
t6aWs/xv7ebbxFRpMICSFAMz7ebOPvpHgvL/Ff8iEan+GsiZzkzyPvosAFnQqNT3wczyevRhQT8t
2FrCOHtrbMnrSnfZHO/NWmT5jbjDlB0KMWEi9ooEvsPNeY3sF4MXBK6Hsm6UbAlqGuRq97eEFOzq
nqTzdJeA/iKR+cFlnF3XKZMXuBNfdNr4v82tvzP50u9aupsbQ0JepA9Zqsqs3supbCPVsWZxWJuI
fn/qDD7i4Nd1L92jQ+btibuojCQgeJGn11N+kyMPmNWjWm4vHtQMtjUnaJni6DjRBv4Sin7LuCDM
8TInzB1FjnqZGkXDmz/rw0TDgmqlCybwg02mGkxepxoPpk0WML7Qn5H1Ydy++lSGlPMlrrVvWr+7
+B6lNHdxnFxEV89QeE5agGuz318s00+hhKaa52sHu4fgMdkUubg7L/D9cexbfyV5KVqbPefQ9rYW
XYm3NPNGFprlx1DUAz4zYHjGzTRQShQJdzZ+VOctTZj4I/fpIbISZBzAIjIkOQ5NMLTnXCA1dBv/
e94FaZHPQz9nsoplA8JqJzgdYwzbRHWH+Y3Fb0Aw9sDrEe74quzJzs7yzbXC/OfCUt7t90aRpUsT
k/4tXEaSNJgSAiFUmbLaLSe8efgv+1FJLyOnB/nnIUW2cx9GvQBF+uNs6sELxPw7TnZGpfsmdzoY
K1NfHuYZZdW1+aoXkLrHl360v1acUAzniyOp0tuSLur9IabOTSTP8aibfjZ7/s9cHoDOifuTBsU9
Sxq5hJroJuRhXTupm5CHrRA2HOjZrwO2/EitPhBC1Qamb9RxMUGsi1FBAhdC0c1h8PkB+NBng7mH
o3oZEsOw3H4c3uxrAfgfSP6y2dURUYBSMgweuFvB1EhBMGVclx4zSSMzeGckZ4FGOS2MkLD6rwfC
2shzAF7AAg6DTEf39/KOXj3lVhAP5VdtCKNjpHMR2HWYxrbh/ENKFadmQuNYPoobSr4EhDjOxUbh
pLlFHQaMUhkaS67+dkDpz/4Mx/jjR6sq9GEr/LpS7q+wR+UgUYHDai/3ljmlDvsvcliGMeKVQ1Nk
R1+B4N+cV+wliQlKeT82VZmza1Tu5ZhD7IghAuEtQIEzJyluXfBgKPBJBkqDTVapeAzokyVFzSRN
7XE5SlkWEUFfkVCtxPiZWT2il0XOLBZ5oPTCApfMMXMsHGjKTsoS7OClZS38jGYeWuhV8bC0hF5s
xz7Q1rmQDyEy5zE4Ayc6g4Jmzw/0MC/DwZ+TKjC0b0S6lLLzGSz33ksJg788GRd2NdgvRScKBs48
8xXGu6XhCn3u9zRAlKf2mNI4lHqhwqpMjewuX5lRyXLjhFSUsLbf3bnQnQEVor83U3bKFIW9kgtj
5uZ+DVteF33ie+bhRQ7A0mJ7ETFnJgQ6+QneD8n4nXqOrKS76Ie3cyAfqyKyXif2FnHZ7TszaGx1
slcDV12XgtDsVOq6eKc8EX+lCWxFNyAagPnQ/ubh88la2/C5k+PU5HRMFV2iTc7cW2YaVJdjAPAp
2X0LgrJSfJICocxKHN+nnXQ1CAYYB9EWN0xY/sKjo0twPInG/uGiWyOdcM7flUl4yYmyqRRxl8Lb
HJQPiXPIm80abShVebYrWlif7PUq0ImjF3IIkLWfH4eK9fsPCuZUsgLPPtovyvsX9Sq5C8u+d9be
+6teZ18yvMXXXEopz0UqpzgSyrdJtbo2MTM7YyxFjXrYQ3tNDiR0wYN+QpsdB/+WkbneURJ/+aDv
FS/H/lgL2NEnO3XSroHJitUHWKxxDaBUuaLAAoKF/PyofvX5tmZ4839PvdtopkAzkT/4mH6efdaK
B1/xlmJjp8V2BucC0NgWiK5ZEyIeZHZMF8XhRg7AkqmxoQY0SQq+3rCFVpqFehmZfcK8e9aH7yzT
Os7k37+rVYjhOw2hqecoazUZU00S8q4IFtsrsNhw8sYEgH+hM/o5haxj/O1HCs9rdcdquC5CJS9J
upsPU1CAcM9VEKN8Mrj0awyrVszdmpnvPn7UmkL+AePuODOOb+PLHMViD4o4MmWh13CJlhfYoiMK
wS1u3Lm7vFCUG/7tGmt+uevI70yGcdkKgm+/CbXO2Gh9pDTfe6DMSsxSLHtZLwTaIeYE90I6sHby
HNVJYueJ6v9HT9xj9hLR1cskCGRyKn6AFkN0O/umLDvVOVOKirLpWAU4V/T6nDyZSGzD6cUTuQp8
jXIfG+hui3DuelsDHMhRn1ht9hz2pF/G6Uco6cKLRqowjxJ1r6IrlaCeV3ZpXfgZDsKoCuYSilZo
Hv8kUPruP4rEqW8frAfhF4ozCyVrdgk5cLI0ooJSuf+KpTY8gQcGn/JJMYvT43KudpxPKggL/Ax0
B3qjE54Gy203j0+KpXTeXbHz60nDJ7g7Ib4OIUj1f8P8BwYSAxk7HyVWzbC/NyfelVGeBbWeJXSD
/fVQRjufFYIiwjNqW8TVl4CslIBEIqAVTV56cuQJ35V/yKaOIfkppkKL8LTXcMSIMVMLbVS94/Kl
A999DYb2CAUHgdvNBiEF/CjS1B+YHzJFmkNbtAMeZVoNZrZ3MdPoLbzi8Qz2iSi4J8zf8QuWn7pn
d92x7R5KTQXn1mwt0EajVbVyqa1EG5s+xRaMAbitmPnV3axrnb/yKh+He6ojPiCD20HzkfKMSFIO
RuOFZsQx8s8bcZ1ca6C9/66NOK1vm0uF3A9j+9wxKZSxYsslF5gsuO7eNG+aA7SuFVZBP4rNMDL/
stLzSaMvC7xS6LQ5NbFqNBQLwLLAdzqmcyzfMNEbuM+gGQCaX5NQPZX/j2suAP3QKoPJG9pGupgi
sP+9sCr651XGkgTYStvvE9ZnsGQMEJJjQPXU0W6zqmzvz5OKS5ySRJV+n3q69mV14aFKtrQH5HUl
/CogVQIqnaMMmgOwbG67oT4P86ihSJrrE2XokpF66JNnhyQc61bCJcS1Z2eCL8VZBZvV26FSJyOq
kiMYJcCWOaDCPX6AVdTzmEXyWvl4aoEXSQgr0ZqWIAHLzNl6NcbFdjmuwwypDcyDZQGaUvzba09P
WbDKggtA9zxS93n0l+IwAyipM7hd0EaPaEvpo7YEAjobEV5zBID3V1HXnvzeUaNrPQogvshMFyvU
+SXX5v7NvCilbuXC4AkPjyQqYB6lj+bimEcY9uqWlbuPRGji+ExE4sSvnYIn29+NPOA1L9T3dGKr
55y3TggEsVPhwpABGu6Ytpv5gtUKw8zWVv85mXLQMgvdR5F0MqGCSOcnO+T19yV1c4V6sVVhOKy7
DTQOsQQK/2vkmuKhtunAq1vqv+2ox6T8fsYRqeMPEN50Vp4bBDxDIx071FUT7PSA4xxCubB5FSQk
99pz82686Vuzu9JvHe/t2+pm9a42FFxBc8fA9m2mM+nBDOe1zYVRrKzNeexUpz6PgYZAGhyhwJv4
M7HTwQvwlozibsmjVCTMjt+3Dq9gEIhM6stDXeTlbMAesdZV4ic0LEox6JxeC4U/1E+cJYROe7lC
2oA/kdGbBNS5QM99++ahjGLCWCgETOv/tY+jX9ccRg1F/k//yXD0Uu6t6yosANqa+1fl3pJD5fvC
mikqfb62811P2LS8QjWzYGMzg+yJLLGRmlM9NfO4B9glu5znBkV2MCNB4P0CU1FtEGCvVBRDIJkj
63p74YzA+IbYE5O0ukG1c0V5/XQuDzmIZ6yC7ppsmvJO7zHQZ83yrXaiDuisU0ngiH6PG/2Rf/IX
bKnUfs9RAm4KXCQByr6RLMht/9uAuzwSWhTs/eRYZad1nDOlIueOfBSJXFtU3+CSKMPBB1s6ShKR
Kvfy6BMxbnKElEONg8lheAoh8h02Ez0YTECmmCUcwblloeafFQ54VGfaRl/jUNf2SUJHQqZw9+qN
gaBfDc8H/HzkYFBA4/IQJOgr7NG9j5ThSX9xTQWc4cWJ2yVdaMJZyX+QhyfdIICxf5bDFI6JP2wm
wt20dscXNqz9VcWK/X/L/4Cw/bmXB3k/WhFBfbOSRSKKYPrAvbYSlGbxrDtU/YlTNy2FdkGxOB9h
oltMZXlROqLrWUQ7jA6VPd8f/oavaj6ucLVZEt3Niaz3YSbakuQwGnGmmDh9YkTCE4LFqGXdwujp
DAPUzjmbdBZBP7/osboyRhxSkXCCTEct6QkIBV89OnzrbCbA31pkYgg980tsGJIcbBDlhE8D4dFH
SLS5q8pfImzw8QZpciKdqxCRqFk1K723VsCMzANwy1UO/yH5KgVftKwj0LkuyUGBIpHdqfwBTB0z
5iRPPbnzD7yADHLgKpj6KbfQDr69TfN81GDOA9Hy/q1+wJtHdRubWiYBxXwibL6jUoWBEhVY7Ipw
d/NuGOGMRZlUTbRRyvfqHPOaQP+SBPmzp6Fa7l/x9n2WTsLNVxWyCjVbOuKeLVqojCdlcjXmXcEp
2eROiWptfIQDXJaw4se8MLFZT0cG7TlLV4cU4oJajXU3XZb5W3tIoGm59iP3nxHkKII7H+w2fi6K
clo1HoZBlGso2dKyje8ruajTZ9pBtORDnvsy/fBThMLdkUoNh77eQE7MorYTrdjT7XTijg7Ba/Nz
VSuHAxAefQiIiYpVNq3vh4Jndb3GLN9jAxJrnrq46IlQo2XZunR4SUbBfQWXSaaUiZOwTmd3gSqg
0oEf4jWWcezPWRQr7nvZSvoAl38T0WUUk/0l6WCLAtP8jO/mnlSotD/SMgWPkelg76W1niRIRU1g
n8djupdjWbinLxMzYNZSY9Ob03G5AKm01bwBk/hILr16WVBqWTd9FzUFYZ6SwXvCB1R41TBKipFP
65wbnfkpyZu8Cf0Nhjr5FHi7EVQE+lvfgPHsr4ZhRjw7hqukWf10eD5RKNy0a4E0y5sYxB62wqgn
ivvcuFHFXWro4UsRU0Fx6Ddip761iG3RwBvegeiE9lcKIh1/8/EngcBFVsQOrxeVM7fua1Tpz18e
VCNZOlXCsX19uqRA6jqjh8UqoGVAl1N4lTA1mojEqxLQyFB9IfTBVMVEpUCJTX6VBrFXkbpe1y0L
PpFWaO3YO5ysVSRiVtI2QF7MsllTyMsh2co8JRBd/109bapx7VM2ncb6WzaiFEGLIP+o1S83qEXX
PdAJu7McSFXyr30peiHCGIo11/KEdvYY6qyqVeKEllhwvml0IY+L40wLe+s/KQZ3o3mtTEHmWWwV
v/ymFdGSGAEuW7xdoslRQyJXn+jNK//DqoV0TgfgwsDEEgMrDUK+ISEofeLznTRb/TLwxK4UXEsc
I0cSrRFx4Q4r/2CNpg+OzVw3FdoMvCP/lMAXNyTv1i0Nyfpj3GIhCpQyDEpquwrH5Q9dPCpp7HbN
b6QwriDFz8BjdzbtEh0IAGM6xJ+H0SK21L82NPwmUpZls1tWm0udIRnYmgM+LK13O7j6xofp/0rF
HWElK6LNH/innV65oAGua4DmmJutQERMw235aI/ZBEd1ulTsg+5cvh+uXLomEywmPgHKr9yhrvdx
uWXUe1AiFGmPWqpAU5MUZmwCcsZ9VbIIGzLdh+OYJQdgrPfJF+D2wGNkX/4rFLhQy9CV4MZfjlxT
OHOvuB0fGR0TbvUWhqq7uRPmpreNmjx962pz7r7eOJWpusd4vRC5gFQ40fT9Z+3n723uZ0/j+qel
sB1grl4muxaPxAaJYPlHqFfpgipxUud+SHnV1i6S/aELC4kLnlgTZrU8ruqI5jdOVCDLufTq6DeL
h8pCdGvdrUtegc5SjM0NJIg62JrtBW/JOd0mZY17Wxz4j5Z8fvSh5PBl53FCQJphVESne7t2nbqr
1I3YnaHxJx5f0gLRevtACkNfOwPDPhDUs0p/j3ezdMOpk+UHBj99FM43RLZiKM+yB0eG06A4YrEl
6s/2O32FQWNBTpQoZm1K9dAcfC3UWxLYScMUqYY8g4Z/puxnACRalsaJ8iaNtdsoirhwrdIV+KHo
5waG0jo0kCSAQUlLUGZpesVamCnrs1z42Dag/wpWEyLa0kYtsW9vC3y8Fn0z2tnCmZmcS7Aqa1Ao
opQuwMnVEQdiwE7ue9GpqBp6L+D5naa0qY8J0bjBjJam+meHtuFw/5mXwvbBZbGH2wLPUOaxkgyQ
aj0haD/1oxeoyFKViGYoWVAlibDgEu7tUMhwc2YcEPYkz3Ir8Qy/EsTKKtQKGr8gbrgAjQXxsmYU
PptAqmfw1AuSD/1OasUU4duSm2sxM52jUGy+JgPlbrf3IY8fsNQKNiudXAi3whfow5vF2wtHbMGk
/eosFxhcEVQ6xWMR1hPWKxlBhJTkXLnTPADfC8IupW8rKPHaHrwvJfcNzjIukj1YlfrIlZtM0TW0
WtqXIntqb5m2N6gItPSBxfKD6BfDiMtDsdv59DvAzuTEVKQ5X/TSbchQMNk0q6iwTLyMclJTWx1F
tKVZ3vCKF8H+qmt35TBY4KcP+3vtizi12npeEm9CmB3501pM+HyVITYt3RsknXGiks9pl6KKnI2z
S2vpx+J5PQg9MN7fnnhD1VuuOsM+i1aMGU+UckiZGA6t6Ar1SKdYE6doRBEy2moXFn8U7wAp/myC
J4wygrbNHfQ4+NfKfcT4i63UAec94xSsE8wCAi8hkyVz2bdADaHd5KsIOcu5u+milvv+o8AYE+YK
DCUoJjw/aluYTDZ1hhIvJINdjrlYLW1MbESkq+DBxT3OyDuKRXcnyQfaYK8pHjQLPcQprLtvv3D5
2/4uC7wxPoX4PSSxRuZzvKClYkibssE6wEjEDKPK/i1xJS+NTAgJVANiEh7n6t4OrG3FmAykL+bD
otkAnNaY0g5mVwL3J4C2UwZlw/Ov2e91r5U4qlqAUJv5p7che3+RxBvBz4tXqJlsVlq7XsFfLC6a
lQrr3ciDWKiazaLVab/ooxEuB4iHip66n/pyJsCq9KE3YXqlJDoO9vvj7rySRnSlbXw7OQEcDlA8
Zi4h/7r1tvNzyZ7BAXy9+kmU7YOR0B8OyodUFgH79dnbVtGoHqHCKGpbTx/MFmqncqFyleSwAfC3
lDq3GqocdrssWOfly7K2+aO88a5Q8i/yP+YTMIojbuOOvy4mfeoA05UahnQUng583dQ3+P+L7pZB
JiAK4+vYq3M4J+mdeF+4/otOX40D/MGWYoJaBq4IE+FtvyxER51/lVxcK+4eRjIOSlSasGTleidz
kf31grYS7L5cJuURF6r3/SDVjS8I8B1iUB+vSK3W8nmt36/XbJJbCK3dV8+W248pZzyejdOefOBq
Qfrda8P72WV1gKyJa+6BmeDE2Rdyvfx/9RLs4i60qXBOaPJzsFN8tdNnnLD2sMpwzmjUll8K0akl
4nqSO4pDItIzug7QWmiv7pOkORbAuYfa4YjY8BS1lQ/227gNqTsZfUX7TUXtCvwSForfgiSIjA41
LlocOA2O+wA93QfKfwgK/5G8UDiwaDwj5uvvWHm4ad+aij3dRkHqBSbwNfqiHbxTTgOSOro3vbUE
TE5eEDIsaWeD624EitB/nqIX62ZRFriY47nf3TgxQyXLUSsxdM0m7/Bm4+Fd6riB/u1y64IF/C8X
u6isS63ECYOgehePLhYYTCBMW2tydg2u+645tQBX/5JKbTt4X7JWI9I1Gn3Dz+NixnZ/+7ui1iwe
9kLf/4HWBv/38NPBsPk8yfKCt9+8275hwlZj2i6eJZk5ZbE8eWuIhDKlTBBOdsNqNWKPBKF6Zv9Y
co3rirRC5SJ4ct0m1jFJmYw4ZiZ6Jl2cFGkBkrPnZyFX0DFI8rfEyCjmnTrNjt35aa5c/AU4UVOR
N2n1+SHgSy0rNuEgj7xK0SyLDWM1Hcq7u/p+zXf9sjZ4KcOB9r+qq/hvS6nlkY5Z81GZW8wdltaF
IQQ0426kvmN1RW86/n+F3UNmTiZBwAIP79A6JnmlZBA/xT/HNkFyIojIA7yq9LBVYHzg7+rHP0vi
lShUGUijDRFxWI14xDdKBy1l6inAma1PMCwjWiZD8ik/b3rxAX9FaGUKg6xHtzQdZnKfQowkG07B
F9cPtB2DEsY0Rj90AGHf6k9wHmwyaw5CA6PmIG35nTImBhjCjp2hUSUwhV7cZbWGcWabIbeVvEME
M+2F9cgzUKKcx1WmuTyVeS2HzhYltwCV5JvmQVmLtaAsAmIiEBz4c4y300w8LTg7XLobskktXISa
BQouCogdmbERpO48cLkaU4rP7i/32Qdde1239uGshrpSboc13rWpMSBdcvbv6pi6hz7Gm+idjOJa
P1eO4S5tvjOiV7fweeh5TpVPJfrVxch93ApiptN1zUnQawvpGzCVa3FdTCmPC+HTtXxK4+p7h+hI
Pebq5wFxItZZIHh4lg7SccewfZrUiAWM88PZqpo8AX3jOJAZAYPVoAYjfqGqo/YR0w+QYHr44zQA
ZHNO7YhWfv1qHLJLV4uvC3yScJzsyrG0x18EnaMFxX6BHvEU+V5tDxwVTmaRNV/kZHn8C1KLVtGG
Lwv52P2QdmuTcYwuSrkQqgNmNDnMgRCLCFOR/vptNczHO7r4LyY0AQGxwXNZY1wUmIrhRuh9ynoN
iKAfbDRQCagUhA4JuJ30t27SF8gbTNxWN9s6DUQzvU6zQKzXBrTIOqFlX0KW75Afb6Y462xQEoft
nzVpbDAMNZV3raNbjIu9B0PIA/fSHEFY7uit+th0qvm+rt3phi36+ovLD3Ot2GjUH/fxt9QhZ9L5
bF9SmkqaEHlBCZx36xJ7h7QiExsNvKEp+7p1L3yISTuEeyrqqL3zyKWbu1/FnwANEOjl8CqVaCxr
1klZI2wxrdHoA1BlG8FRQ+0DUEcd3vQ0usuI3Qqz7lxvH3s3TfgKukjyFdEotz6ObD0NcZi6CoDl
07ALoqS5iCZkS9Ipti14R3mJQqrSkQdvJEzHlL/zlagprwoTewUUpY6EWWQv7FHIVUG8tB/fGqSg
9p5pug4pttYZ862haPIs9ObEA3YPizk4FwuOlpiPTuCuT8afOOLjwXkOvRsMR+oZxDNtUIoziFSn
KN86Un8ahiQwz39MqSUyRgH6bEUVvJPQbjdWvwZYe/C4sWYgwAmzHEG/Kofm0VQ1cQr3gi2Scysg
1IL/Awr1f4tKZm3ezvDyv41eLfpbYlH2ORTnsBGgPnIWAYeJhqXk/eKZ56agRaU/7cypxrjq1wxL
dKg9KezFwoT3ilgCkAogvlK5cz3ZZCr2mJGmCllyxWtNVLefl7XYNjVaEbGGpJXopkfSZA7WxNMx
28wLHfHvKdbUpi0macOwWkykwY+BjevRFomRJsGkvrHFgwuvxPUig2Uw1NMt3suhbCEibSR3W3A8
CTztnNgbh6owQKbDW8P5s7UdnBEmoSwC1j2SsThHeeFJwe4jXXm0L7T81fR4emzKw2XqMxVLmw81
aB1cSU9IHIweV9VhiFTHxdQX8xyrRHWrlazn5GAiDUM7maXG7tQoIZxP68YARex5p5QGF/BY/wfG
AcAzpla1IKpNz8v/Rci2pCxWvK5Hrd8Syga0G+yU4W0lm7hchvAprcWJH7369HQhzcsZEuZAszHs
LNloQTkShiuKKT6GBGSU/DPw4UStaX3UPBda41y50RZnrKwtNWeFKJs7GoMXSkPfvYKyGosyRuh5
zex5vNO9jbQv/3YRMS4tfSObOLf6nBx+d4yjFjuvgmZZRRVixiPSLM/6ofjkusps1XvSYXVirE7X
tjE1yvneYpiNeEhLXUt0drtW+oc43F5XZ7mSc5LL/dd2nwUt+MjK8Fuuu/k6+EJZtgAakBY4mNpS
uu8Q8FlfSQ/3uQgwOhvXayBB9Y6ZOQDg7y6t+QrKx4dn4LL/McbiBp2HnTofwyp2u79riQpCIUOb
aUhEBf2ayjuOLDy1ID4nbipP2jNwGRIGWZ2iB5TobNEIuX5FiHBul5d8/1OxnhOk2VVMKj3XsLtU
JAxPdlJN9L9f6tk2i4nRRPMWQb+STCEMH0oV2vtSc5x7HCTScl7ej2FUV45sTWwkGVS8iaT0d3mM
zzdge2UqEoVxLEY/YQOMMuCLZAi10527+Bh8Y2O6lipiG6kKTXVChguMX21cYx+7Ol2rglvsXdOb
Q5+IyTleT5smWFUaoFguoSJpLMc89gzusnHh1cXHxwIK+9USvG/jYDyIekpEIL5+tuQAkitm67Jp
X3PUAtTRdidW/gLr0gQ7QOcoEy0e7L353tVuc5vkPb9d8bWFm3v2iPdn8WhCaVQKB1iWCLM6kw5H
4JCxcONYXGlQmu5l+Fq2v2vdiSlXCFqz8g1hfpAqNyW06w524HwvrUht9wqH9PtfJ05SpgBH2ApM
LygpaZehStmJn/InhE49RU18vWPy0UxP9xhuCtvuuN+r81tkXdDtQxXXk7wdLizh2qbhh19jNQX1
m02CoT77MWVtAJpxUwp0bP6o/v35TF2ZAqJxpCQxAqIiqJwWuU0/8pkEuZZbbVcJAKpizRdQADw2
dk3blnT64Pq3q+FN3Z+MAEIc9x+GU7cm6biACWEAWRY6fcc3xBHFTX/Bg3hcii76sMf4FbiW63IK
6btKV8Aqg+D/TigIldNvGTDinIfMbMvNEaDkK8ANHE8F0pWJB8oFvRO7O09r90vmueIYttkMf7p/
hDJrjF7m+/dSe88yG8/QF1QaitRBtG90nb0iHt0siMRbWFwZ7ahgEatVnQCmXmLwAV/dnKn9mX8m
1YunkLIeKGBlxqczkMWWqhpbvCX7vkVi9Zbpv+YmzcHQZcnOfNvykcqZQxbPmknrlXdGK4gXcm9w
u5F2YfxUu4Lat+ukC+Ro33kv6b4TNLNhyoUPxBBChv2ENfslZqMPMvrepWYze1OIO/NbuVA2y7Rr
jSnHk42NgQi553XB5lBd4fIgDCswcrNI3AB1nxA87jAeDJQTAbwrIA0wBdVsOSlheljWKzju+pAA
gGp+tLi8vWNg6i+AW7yE0r10y/8pJRKyayBQAXTUf0PDwNSZoRdJjpDCcGkr5fTrw7taxZeaUTCc
16TgHyFJVs67hC4JYoI764wM/7X+xEq91Db4kElhVsmT2KkhGBeziyUlxmUI72IMUxENwp3vN8aC
rkLQRmuss0vpxFo77DY5J5JpLWLg57LFBdO9QVtn42toY62D456LisZAweqw16u0E+vhQBYSI5Am
jGnB/5weKcF6YXlsOyEisqiBbpkSfpG5XTnGnxeDlJISteqggzz5SGQOzGbkarY/nML0EWLZrfjl
sAYdZ+NAsOE/u3bDbz58swyXzJqfauJq2vcQuoiQHtVqhl2VfQaFil7wAZbDS+ZvDumq3A7HUxAN
B+G3+80EwAlLr5SPj+0Byd18HEQwn/HOSIaGA55ZVDQ6UEIyILA5biyS9ey6J4UBRsqGOIyzwGUe
KuZIw0QnhtBqt2JvOftCXeMyBw2TdzclkcpzDB43CK32AQI6GuoFH1tDrNubzeRBRTQN5SR1YL0S
UnC3TEfcv23cqZqDFC7dSqBxN7Ko1T4KCyrE7kTFMl5DEBvoToKOovIqeNj0tAhdpLNZ5CnBDjR4
A7vn8Hxbi1VKV5mDwJPIC9vNQ0EMBm5Jt/r9xObmKN6BkVf0AHAza13W2bE5BLOa2Q+y6xBJiO4j
QYrvD6xSmedSOcyqiJ77c25X4EJ1tAAwL/ACgdpIU/SI6X1Ygi615x+DeLFESfQEIXm/X/bbxChZ
2U+apBn4eTMMtHtt15cWH9p6nYh+AESBwjHpUyRyO8pqDfRNc3MUkzbtWtBwfBvXuE4HIkM/ABSQ
XcLN3kPGJ/LGpCdYC+TKyYmiPuWF2uUXgEeuBUAnCXhOvxnx/qG8EXfbKR47c0tRQIUWeedLfm28
jPObnSLyXXjiRtSyKYu+Nh+8n/LhA5drcZRen8p6YsBivLp+/cNdm3fcVAp97RBnDOexAraiNljU
MYlCLzHE0GSUk61Wkc9DMKiSrQuPZuMS3301Ou2fUQcKTAJRSvKgcE7KXoCfVGUyH3BF4mEnoYAG
kXDyvuD9jBOUWIw96JASlVIWCOJ0wFnV+khUTeqNqr+2cNS4cfjn7ReKdneuqNuih9XcTL6vIMcV
u9DC8a25taAmH2P1bdjMPSPfFYY5JS2Hpz7URAYI6j0lqA4lDx6qExqL329j4eLrQfOj/0w87i1k
pgeuQPfM2kzFJi0fhgoO13bo26GZ4hTHLu3UqUAU2JFn3ctq4DkWBE64m9uyHSf/zdShKrQ6yzmP
a5SkWM8jNOvioYl2RICUkuXagm8Jb4wWPsShaaPo8L9bXvlpH0351F5+gbW2YWYLgff3j2kcj0RM
V/4OCp2yjs8F0LWhYCtybc7L7IORdCTF3P4B7WQn7BGY2s4BLcpia3oNtXsjiFCD652KckuqS2TX
aws2yEARK+CllNfCDVs1EHiJ/aOnc+jWeIOXx+WlhS8Y8QUJQ0fw/5wrUM3fDj4/5daS7fcMV67s
sswxTI+NoKM91khSPrdRqbtC1hccp8VP1jycI77KLRwRAAepV1zLVQ/JbdqVLq4/+28jgzm2OR/u
jZEDEP0QmMyDwoZ7rHjdu/kfaJqQXvkVYcjQ7d3H45aAQ4+Duue2ebVZuK8vW56gDfhju+N+z4+9
ld3RAaw5MlejazmJexkE8g7UVq/ehURrMPXCr5m2hLmPWvX1ef3YEy+bAlIaZ2ZRlbQMFkWM20lk
CxS80Ba5dC0Fhq39neEH/IvojY5um1Z6nKniVzYxhxxH9cN3jb+hcNfNEFRrt6FeXRGkhGLpDXk3
3YpvDZv19Jt6X+DcCQ0JRSRhPxlRGmhbCaKD/JnkMf0yy1rii3w9zkWAj3lPJ6EF0Md/PnhAGYYM
Nkak8lQPjrbCy7WIyP479Z76pBFvbIfefLtTCE/t2Y3+b7KCCpa7obJeFgPuDdpU9J7ATi2oCtUk
OfEl5wuobj71RVdAjn+Npa9Hg5YV+5LD+Ke6ijbkkZ3nLJCQpg1GxL7GPYnHfnLx6mLXyOpSFU4/
4CnufCLlnEJCflDV/xC9MsvvRxy3CUeTqW0uMM1nfYZ4G1PwvlWaT0D1MM9n2PBuRV0VWn0tV1fN
0/JMf5bakMOHiffe4YWEjcNinSbgzG4ReEpi1od+5gOyR577+83w4v3CMF62nLamNx2h88X/zizi
WMbSOjzSMuXhYEZs+ZIpaOR3uRIpCIlLXhd3rG7n3bLlaXLTnd/ovv57OY+Y+P8evfuRKDDaVC0x
t1c7hoyCylRVcE+T14CIqf7vnXoT2MmN3EY/dJXb8d9sfvPyq4qruNtTuAy6Cap4cn2mVudk3D9t
ky57ij7dbp/7pPwBYmblj+JW4FosQqCJgOexDam67NLePnY+wRDn2tlIJh4ELpyUdtdQRR2zdVuI
dObrHiB3eYLXtwHx8JU/ExvV/DnGQaYBj3MnIglPIT8iNiZcvksHha6E/Rm52SWvrstf+q6WE+tm
Mfs97JHJlKMh0hyP/RJI4ymo9vLqPEUZOyn1peI25KicXEzi9m8vSM650HTSaeb3/D/QKL64aBai
DBJb8UJCRtpIUOhWxZqqHYu3rqVTtKhj3iA5JX4pSzV7oyEdGtEtnM+OSBWWNftV7ZkiFM2HmFHv
pnRX+CRsMgN7dR+JU1JTJ1aBvMDN42Jd9js14EpjjPcZMKDEh0ruGVR75SP97XV22EmWEPzYYjcw
3o1XRgt4c5Oz1I2xn0T4g6EPpdgciGIKEx+yzyH2cmS5cB3wBs80k8dZtzbLICMSA96GbtWMD6ic
bPON9udocoeoDeWxZM8ZY93OKoASPLC9HNClqD50133IrAxVnTDTBYi6oB7x7prygwz3Hb41/Kb+
BoIfX+z2ue2HoqK/rEL/kTDMPle+M3+cHheVf2+RS3+Jh738OOB32C2n6RPJthV54E8Dts4RSSqr
lGRLEQYX+794UKx/u+CTKufvDKmgVa5VRWLTDfOuRh6XgmnU6jweihewjKYVVhYHoZL9f7EDD2XE
8zt3E1AhJFscgNiLmhvDMopOr2M2GFJvsTTIP2WyvvcI/YkKA7T1HhQkkoECKa4UNvJ4F+lhHbMT
XlDT2EMAGxqXZlOFuTK1caNIj94GQnCxIdmcqOCnhgPdsMTXgPTtiMYW2rA5E9DYqPyiTjU61IRG
KoFXR3NAfBlOeH9KB5Pl7OBpD/QT7Lt5DyyrrYjMqJApvRbCbWFaVyV5781jH3eZR9xzm0plnPIk
DA6TBw4ZsjlDdXksCb7IfKnefAYyNMOa22MTm4ljwoF8e3kReU52cWomc4F90279p0wn2FtYAqtd
79B7xiBkuyLSn0YI5xKv+KsTEsMkB040uLJ0u9656ClBI2CqGwQtFd6dTKelIOAMk2us1yUp5oU/
szChjNGhw7HovAp/wjxNCuFknc038vxtxFH0394JDe36IQpI6QucdoNVMHdDcGxc3iUV5OSGAgP6
9XZp7zZeOn3E1qiyEUbAh5NQiEIPY5LXOQzWPC4c7FHqHooEmODC5UPep2/yuVrnNe6twhB/aeVI
HQ/xJcyaQlm+IiM3+91aEsVO+BGCK8cKypVj/UadtomNYhTpe9DYEAXrCDvjVgrco8yjZy3NN1sa
ay2HHGdx1Gl0ooowEEgtjllJR4f2SMDYzdPMKbj6qpg6+Q8mx6uDKOBDUBphcx4p4/15aHMInY0G
Mfh8RPYZ/dkqloBHr7bIwDggvw0jC2ivJzoFqGJMPpaYUirRgcqseTi2HiDpyiII1f/8MJPmBbEb
2fmQyUwuNNQQFbmUGNoMIHYvjl/pJEnA7JTczEhwrbwHTe2gAuAuWKbRz1t6CX4cMMGBUe4eBYls
3MRhycHtncRshiLUGFYnaUfdjnMg3/7Eq4VIKqFGlHhNl0OsPw40/phNvlBdAR5yShHzqZcp2JZr
HfhCn2+n/ZoneLxDnGQwZiLD4EUjZK14ufBHM7zxSCAXs4e2cPqFbz/Yds9yEYJB2x1gZdj1Dor7
A11eBw5wwG2rmptW2RTf+kyJlLGWA7FAxpukq8Q3jBD3x8yUmL3jyK8kfEvKjpcafinKvFWz7wPE
I2VUzimY+6pcMv3/nZSHq20Wh2cZqbkVQZDleT+t/0ahsBzKFhKYznWtjBHWJJXCsa5Q8ZKUNuEb
GjYoSli6gUQXPrm5bjz5tcGvmlFJJhWa1NLgg/1iL6Ze13fruN48+ML3kIZVfGFy5At1diEYyjWc
hUG0S3oZJfgyhWPJefA75T4ltE/F2fZdIY7YMQJs76/d2zxQB997jVwUuD6aCIt2YAd0+VyfSImT
vUDz7zwLSnT2Gis2jsnQG5q8I7BXpBhTgKcDS76g41XjZiLW7/zuBVyI3dYtn/4hqeTvUF04vmY0
Br0v3jn2W9lYa4ZfFL5LUcUJ2TkkY7ATtx4XxHe6S/J3VhZA7cHwBhninvU/FOdJ4X6IFxriVXX8
qvM4CqPWy9UETeZ+C2uEa7phVWbgOTMOCiN7YBs9D+rVELFIwqB63ivEnz+V/7xFBOEbwpLWTWuT
txsljckkgrR8F5vgsqaCUaHMMhXSvgjrawEhZaPDrR5o/gxWZ4USsnHRTsCk7yySP1xO3oew1SQm
2iRVFcz/fdNZm9y9pXSOz+wwLJVTfCD9mDEnCI3imGarYnMdw4PVshDNLIUhqWmlJSEesJHGZqWH
ZYkZs5xLa46zdXvuVgGXy4ffrfgQy2TSOi2vdXJg4hJ5dWbhNdBZhCMLxI/dOnfKukeZvHABI7sa
67zS8Iar1ceZyUAKy6woWw4k+GWdiMH+2HzkwbhIMIL7cvDq4HReE4M5qbSATjq11YVt/cCarX9L
pmi73FkhdZePF7snJz5hkAa4ndQdLnIEV+WHtYEIv+vF10tVsuF9lRa0OmMjH6lr/TbND9MTLiyF
mYQ/dk49tQUWSa1RyFa+TQWA93ifJvUMGjd9l7pDN6sswSmNCbrpCeAWxyQQ48me0p1lAR49NNHs
3IYMpmO5LBiNeeuosrliPFANO9E3Y36az2rACP1sqxH1nitqHBDNm5UCzDmukA/31IqqK7OY3NVJ
AEeqlMEwG6VLULWgHRSVPyzomv0pl1jys8yMv16aUMZjSXJxarTa3UxWCrxE95zrtLsChbvjIEh0
XyUm/3Pu6dYp1PgMcUbBn1nSHlwueCb9I9NTDMdqViGqC4I2Hm0agzYGJnp5vVKicdDgNJjuCp0J
TBWa6K7VzUTUsJF6lJpsxOxGygcVq2zGSTxURp975PA4OIvDo9ybghTTtQzfrIc/8zOKKWPvkQbu
/3jfFvcXIAOTFdJkB8nkVE/MbJ6vL9IyloKBp4EmUv+1ssY9Zy1IK3HJGN2tF9QQfdGwKI+VVKtw
q0b9HJgMhyPTdhEEd5FYvRUGJAJosVmGGf1y6Fhyltu8FSIp8/kfq944zNsfVmn8G9anLFQ7YDrx
7CJRtDjuOw2EaGt1QGJOc6sWqdHskCuGLbzyNmqAIalqSJReeCkR4aYR9KckC/X4zv7oDVL4R8qu
mJYtDOa3vkKCUszlp5o0zytF7goiQYdIVw5t23xb1gn3o3Ad8qx/CEhT3cYT7JxIQJKDW2iXiA60
BKY9XpofYkNpUajEtwNTmfuXDySxq7eR5yNDUN7D9b4I8aK8HDgD90RclTnXr3KYKE/AlaFXKs1Q
9aRF2O8SkMXC37qzOsRb0Id8HWwCT2QEj4f1h/5hAcl+KFKhS+bGd3w9Xd2TLL3x+d/lkIUTtsg3
L/aW+9Efu/u2mm1tOBItiZc92qPKLBSWqK51QlflVzP4CVzUZXtdMWYnSRINKt1O/LZfz0PV3XDq
l7mRWiqdX5LLx2C1m0+cwAHTb7EgXhzOe9YtWTa+sMus6UjOhkAJ20iAaJkB9fM5u4jvjoqFCDpR
R9OTNPrOhf+Uv9KcNpgQ01rG3WaEsJLU9ubkLxTyEmfDeydwES+DyS7IwVIZB/BrOKlXSzYhXGHR
fndPmlURCpkWlt5iq68xzLwBtXDL4Xe1/bQe5pFGThlAyhalqn+q7DGWqFFsiaUlpoZ7piYVPSay
fqIMh/hBygKUl96VL/9ntnv1MpoiKhBCWhjVyjb5LtUBQtXhGPYfkyrw58/oCSB/Tq9jQPjkJfv8
pH0ji5Zw8e+6wOLIdYU8KAt92OzErgXv9MMZ+3uCwLQJDA8KdOdeEGSoSVkLCq9y5KgZs506UQ9l
nx2Q3hjC/s/0pn4/M0j7cJYjEXK6KBusisWybv376ICBGfnDsUz1H9bJhj8e5hqpBKw0k76bZP2N
QIOJo0hPsZ8Eu32Cb/l5TzKv8JrgLVcMNsuFmfTjJGWjX0BHGDeYEFKggbYC/0FZ706H72u4/BI+
QpVQfYdzznDkFctYAMbUFWlKWmHg/kVd3jqB9bzLDQjRKljNXWFNk8fSd9B79B28wtFg9OcghRxP
FG+N9Q1xRdn3MKjc9GCVxEOc3rSI7Xd2XbOAWiiDxC3k/J7IuiUapaSplf1tabzFKYDPusDKw7RL
HC7yQTYeksFTdghT6IL9d6sze8PPxE5bS2w9mSzCPQm00s96JCJtz/i1mfVr/vGRhvcJ5w0xh3D9
4iH9VKyuIQ/WXeyR2FPHnbjhIylrNs/QUoqGgPOto+S/YdTEMPyEZx/ZVBTFUhXBoUhKaKh/yuBY
g1jBLV6ra7g1U6+R5ARRXYfd4Rvjnva7qDQ36NbeNrdQmFZGhof5h7bozGZcOy2H3AfqlkKnSEzH
HI7YVkY+8InW99la/JuJgXlDZI/jgMKkAXVmCul+IiaQpRToiEcfbqnXl++hfDNxUqy71l/hM94t
Ae+kLJJ3GhDZX1KQW1e8zN/0XyCs+vzZhQSXVD/XrH+LXtdCBM91zgjbD5/MaTB7fOJs6SGcsMJU
oaAXiNNbhCAZBFvYKuFHKw7a6N/gUSpS3dsSdMRcQcn+6L/ux7/p/O65xEM8nxWDX+oLNaunG6hp
l81J72RNzmQtyY+r79uxmekqS6nmATGv5Pe3ICdp9KPJy0Svp0rrzUxAFEojWj5svgD0Ey5tl5Td
AM5GTPRM/12Rc3Ci+xc+A/kTh0td8IeX28ejP7TmqnWbVGuQqeFtXbk4Paj8Z6VNwvFWu96QIATW
ZyuSlW4+p2Jw8NZXruPCN1kndTe8c++WhEzBIzVGhrGVgkrlhlfQ1iYd4QvC31ChEYC3MPqCezCX
TQShVW3VPpG0Kwpc/JHRWbbwXYqOB0/zxBiHz3jS9OouvZzOk8Wz0nA+XWy1f4sxF75/en6un+jY
lrHjtQxNn/c+ttGxSRza7mk5Hqt6JYZw8r4AOoK39Nx/0q7gcWtjdPvvktAvZhh8okWEjsSYkqrl
gZoAo/GL+9v502vdcT6IcLVgJx/yd8NyrN3W9YgRYc0vUfcZwdOMjS0mzIxPb2H5Ld1SBxlwv/ku
5tRvYAU2GGybGgBgO9AlrsEuC6+Nr7FRept/pszkirDZmXjDkaYVK8NArAt50VxCRJ0Y0mEP5Ymi
rEdDSlyw40yVmvSggJuIMaxA18EQJHtN0ShUY54hgtBp9E/DUZZcBpSJBHaZAcAELbN+lgM8PeJR
JEeb2eJS0M+5cVytYUgX4+yGOqd8eHPjSO/7BPD/PS9fWD9eENmhlbjuHuPhqset4/U01tkuR2ue
rLxUiFPe9HthhQ0FKlkb4wjwyMczb/y6x6adlnQTM4ewJG5l9djHgjI4pEIhmnQyUtKCpRVozk3I
t74MYXDl3lR6mhpyrrWzyZMQYdad+j/d4Uu59+yMOIwRWJsdjMqZXcGDFENv1y21ySFcXsug9x/v
jPd8nfFOQg/86xx0ph9h05B0E05+aBeSvy1+Je4IeMzc1dcbAg8R4vEhmI2kJWcsBkDPa6YiN3vV
dKQ4b2YQv+WRpX3ZnYCW1SUeBqpDBI8e7YKWihYpUiKiU+Aguq5N7sWY+A395rwsftPhk2pPb7KK
PUXHoo5LrTwOuQTRsDVRU+p7d6o5se+Vb8p/Xa2Cmr3haTJwtVfxEU3ucZRDiHUvLi1xQm6PyHUd
dPklRujFXt/3Caq7yQzJ5ii1RCSconbpzDoq+AGbebp2upvq1GLq3PoCO10jlC8ZnEQvmnsQygyP
NcEPje4Yv85/woyikgkPrM/eYZz2b1H4t2lf7MFhGhvkQProwdmylVe9uWuUm9JtpXsdx8hY0Mxt
4i7eg18jzxP2lJ+XAHIniVBv+uXQL85UIxWCAWijpRz/x3PdR2bQLwAOVUMLASirBIVvjxd3I/6h
nWB+YrAIzy0yZvlwbQeM1k1k7IeJfpqHa5ExMUdPbfteBn+lyvXrQJqZvd7G/UVVcbGLqOxdWqBY
ZcPdDWyqGDKq4CudqkA9ON3o/ndC5KJ0JNLr2DWcGHgXFz9FK2LfCNG3gZLfS607wN+MHl9p5ql+
tbzmJJjco3opJ87wYQ10soIB9NGP/DNJsMa09p8OY38MxGxTIzelGcHITHt+4yq0/SpowdgBsNzQ
tOmZSMQkQyJpavyR90uXak1KVU/UXdj5tUEKvZCrHYZIBJ+kGy9kHw4Ajk7+Od393Alg4K2KN1X/
tgtxU3gLAs4LIdqykWGQbBVMlNnlOr/9h5zzbvDj4X/f66vhdPKY/GIWqVAUb2jNvHyVT/SYkn8J
niL1WvED3EcItgatsdQ8+0h8JXSNZnF6n+oxwZg+Yv11XlD9wLLYTUcyjdqZzEqLy+kAwOrqRY1I
yqcz7/+F/qy4AaXaaQU+HxBKAdpH/LiV3As6n8T0FYA3kHDb1qzySco+llRMirm0SodTlBFbwgAI
vOOeSCIDjNj/wqu4dxSSgee7FjJmXcGTKPJjRFKh86CXVUUzGBZRP7yefe1fhsmpPF2/qaT4+ATY
ry81p+CTDKMPaazuiKmPuk8NfqT33uNvPxhSsskyd7IESJaO22WFaZc1SeRdcIYKqHM7nPRO7F+K
n9C4wPlmJD0x+Oo6N4STjlEexC7Al6U6cGnXRQJJXyuAEvjjmpPvMYrI/e0GOFsRZPdwmkxpbpSC
1szYJb6xJZZdIEy8Xe/hvStPLzzVXnqONKB1U31gSxTeZR15WADH/f+PhNhlv0Qjlg2I2BvmeBU5
xNq632uVWU8QVyw2Zw48hobbJJjBa2IWK83QpODu0B3MrMcqECZZDwAfSMYOvbXy/tyxyg5c+Fnf
eFvldrhZapZ4GB3TX8CvxR7ZDggaHtypxJsuVLUgVF/ojx7YQ5FY7XaKh431P3UUviNAVA0zFjtx
YRu6y0+WtwY7nN7jusArWflCWrcmxkddnh1GYkKVW8m3JUCCcbXlZKuVqFDA/nLSL7BZOIwkCQWA
lsbkDfz5RpCPSFLnwOkthF8ppTzbY6aQTX1fEqDTe8p2zBK0wQoBkC9KPMnba6v4JULMKRNfnwxQ
q+haQem3LgO+TphF6IOUWvoHSEzEUr7CJQca1q0tzR81YRBOUXPvZ/6s7iie7KG3xwRuLdQjp2j1
MPl2VlZDwfYXOnwWD1GxluDJP+Fh4ZRD/eof74g8oyX1qwD11U+1CSaxXKKhdhEWnnsgEQ4rVIX+
naI/lY0UUU5wNL37CAEILGgtJVv6pzpxRdMPaVuFfXrfOTDsoSfwWdISJ8RqbT+hFmngvWecn7Sh
XBRLASAk9H4PmC0GMxeIavWJjWd0VwF6RFfNaHzVoXDRafmFFTVSET3MY7AoW/IpHcI7D48HlyN6
ZttNWgXuDeCjkFqumrO6suO9IudqxNi++veKd+Mt2XCF4Iy38kr4WuUXhhrMZCT55kI7q4ZLxZYY
lspU0lPJwQOWZChbpkKxe/djxp2vyerFzj80bElW0O2sqpDhOz9BXykN0YvRq2iarafE3FGx7n4I
TK1GF2CvjgEnL34fQmZvMSAtzPZkr4jtSA994lqVhlRorMeXWVol4NXmYJf3AV1/2QRrpJV0U8re
mOk39irQlUmoOLM3SIjb8IbLYxMd1yOk1qFwu9FhWEbduMC6QLphiGFEdNOz2SdOolzXj7pNCKKj
t2osmT+mpnZ4TqM+kRk4auZrb4CI/9+lj84qFVCSPigFlL5q48yDbeicxTXwiqs6bfU6gtBwmNS+
wzAOQ8zDDtkOUygVJShSej88JqVtW0JwZFFjlDPar0S3aXtxefupEsPADMbnVjwIAzXY5lKrAKJF
N4ylqrQQQQ1BsGo3NlQA+QnGmITUmBqMZ3pT3MVAZc6pNDZ+kFaSzvfEdJqiaJEEBMI8eSAK4Sd7
DAU5UvXDEcdzBB26QxxnwAtVvGRjsj0G9gNqOSEzHLYKoQORcNfndXEgrkd65vfCDugUChG2W5uk
ppRde4Tqcl3GyDMx4xG+BXX8q0d/8PFLMq/bPxacZEI8ngjd5QKn5tbeaA6ynsJXxTQ2e/d77oeW
lUfCCgzVG4X5twV9OEa8pLq0gjK1oaXSvLJrGR3sPNFtXh5dtZSKIbPftpTAfTnfYFw57Og2fmcJ
FIZE4EaODoGWw1aHBYrnXyIEiVU3h3Sgj1l0OBGE+E+D88lccNBCT+VNm3TR2rqwS243+w9+V1wX
QDWEIQvoudE0+QrHREsfZOIzgE7QneTz02rapZHzHlzdMTDUNMDxbGGZZKzTNlY/oun8T3M4thX7
5KReIXSeFk89EOKeyaCee0reavxoGMTLiGXvF6JpeVEbELfV7HaHO0Fdft8+4Wsz9RQSB+yGFZLG
myIo5+0d6sSgWs6+7tdflDBDSW6raYdszv9Fk/aDYDTu9ENI7fKbU2Uwrnpy29H52Xbv4FwU6cSY
HFDz5A6kLYGnCfWq5njBjVNVMOkjy1Wnb4MlXQSlBeqBi+6qEA7R7ceoXPFAz0OM/TGEGH50+FFF
5yE2X+vzE3rRp2/ApBExc3YA+JvtnprOUjvSyGrkqcr5X3p1+jlvQwTpkUATQZqLFYQ2Eq+I4AoG
cedOWmRjxTbCya4rPBg2yYVKUf+pOvmIUQqHGG/Q2G/A+PyF0ZYTZioPlCO6jslE4wC0RhPdxZ9z
lkUMEYFe+ztrtwVlENDhhUJmWqFRI5rjY3aNt7wOnQgeCz07kcwxL69hnKfEdAnmbnkGM+R2mK1V
OG4mDdTEVOUCxzFrz3mD05WXThg4CUrH4/N6K5HqoDf+euQ1YHon13dqa9MPbFK4LDP0Tl8iEiLx
EX9dtLqfqDM5UT3msd1TK0xHgcbP01njpR++yIeSUQfGYsa3JqrrebxwVOzmOpniOLFu26e1rzDR
AurZSHgVYQQwl+2uaZW9jhppyVRA0RYzLJnLzlUHf3CcKYTtKa249YdUKsjIz1C4Mo2tpyiTl763
IGR8QEdkM3TyRYFOxF9lBv4/c4P2cuglaPT+ZhWzRuqLbzj9p4ytelnVkVwjLrotpUSnkYLbOfsB
nQjXHy5Qk8ZNr0TUPuo1dMPsnYkhlQPsuXEZtMobrvuAGaRrITORb5vMGhY95Nob1FEmmDQvCR0o
NIc+opTJ5833xvBhvy0atpQYDlsk0KlQZBQuYIqWrBvbBLYeMuWrSyZxdnFue8HCRRcidfYsvw5l
+M3CBjyEUNdUb4ECEclSiPXh+bWhilMj4NKlM2CSfQk5tculgasEJPwfgv3TTyxlqbqCX1Xfm2j7
+6mwuC4ojJiUbbU6ZoIsnijH9PqqecsnUCUxz74CdULRUUcjbiwDAQbl0mmJtqWpvlwbXMNlohE1
UsUZabLUfhsmT3lLoqw8Qt/4ILFgV2t0nIu6PLAKns1y+BE7Op+ugY4+Gtfp2sZsqddrGLUlkg07
l5uMgDuHiPlOGzLXxxXjdeeMcvH9TUZbtpVl21tQwfL0TMTukxGacXjGFIUmnJYBuc8RBpyrH6wf
CrEAGBNtN/EIHCa2hAQ8W+3Ty4djsSDNJr2ZBBp6u55VugTBDDp6NRXl2vieJmWzrdD2/LzK0DFx
DYv7svWHhiKvY5rkK7yZkR/v7nhaHU3fVoQiOnmafhnlETnj3CnOUeW1cMbMbbQeDIIRtCAIKOr5
qvrn0PFX8In62e5Jpdo5RvisGUgDfAO04jhggIgFzgmf5ZrNbYAgkKNQNyqjilW6rV14DE1sEjj6
I/bTs/QonYut28AWseN4cV8hArXL4x6vA4wtP38s+kXsdnrvz+We6siytsOFtNGw5EFj93wGlAZ5
apkrjJ+eSh94rjbJQ2BCGg4erUJLYhs0mklmEv8hNkMA8GhnnygbpDC8B43/9xCN0tEFJNZakuYQ
c+yJLYiXDJeM18jQeUJNiGriHGfvlSL8LTpich86wZ2WiyulsfgySqgqEYQEh/3mZvN980pXjvYj
QDUt94uNrCTFNBRq7ItL2pPPXkvv3FOvXMYDalXCDSxpIZZOKwstG6/9tyKaOs6B3kEc2oDK+D1+
ONzCDCWvFC9wRu19xqSMn1539wtSzOx0QE+ZEcXZvfFL2GY+qqAUG3A8UdTZk9wU2BLiMSWlr6HK
7r4I8BC7oddCCS4N4fRtt6LWdQFDq1q9l7J4HVOQD+cNxihtKw0MMwCXOgzR4fFMl/AZcAanhSPM
bxDTZKvTbo5rdMY1Ks6wbieOk5kQToYdL6vehi4+2JXLwc5azD5tHzcjvwu6XRhKFcsOKBdPwe0R
ZVyYFDF3Nle0Guy/5pHHFl0BV/I+1A1kycwvusaFCLwZhhCoV/vJsrz5nuTdWPs7pGk8QRYCFMWo
u1K6Cxj31yuIU2hV6nLuC1FLymGOj33v6M6wCkYKTPKPasbtovW5mqH2R3xmOGQGM/6szHCFW1Sh
bmWqletGHQjxiFz1vEo3F5enxzXqE6sUcJe3FamsRF+TWA6LK6GfNEsaRIIzNXfXi1hhSr5RHj3U
pCQZAXhsJFWZ2f/aDXCjA79zHJnFtdewTg21O6+YnRr76+pzQNGhgCJas1XF5k/85qj0iLvRT5hy
ghI1DopU+quDT23h9MEUGOYWiulOJSaEiLLPzLykJ7ciaGuExCEGp5/QJB45xcx5tteFvVWckOfQ
3GAhYtZpjHphJmdRoI1kvNSFw9gR4kc3O8s28YSCXwLbtmBEEe0SZmIyYREdowlKbP30qhuTmD/C
bea7BTeCtsfBW01W+z+paDp+Ao597KhZZ94CivEG5MX/IfrMkDS1dpy+d9FhfwkUw0YadseUrzhl
vByMCDny2X1rQNw4xyAkZtMlP/oQtivGYpGoQDY6ty02OKF8fZImc6PH2uNvbf+fwjDcmtzO0B1i
LA0RVCetsiAm/MNdkRjGvlZdOJnMZQbMGRC5hPUjbQRCIqZWrn9/2OMFAwG/r03M5B7llaDDGp4W
7GR6y8/UZskoDTscRPM9hMmDgltymdm/MsW6+Sjm4DOcKL97q9vcS59oPIwfHpadt67b39WGW/jO
/IhpUVU6tZmQCcj4cfQixyC8qUZ0M2aN2lQgx5RdvmMvMGSnz1YlayheNeiCzaEPL8Rz44hjyzjb
Bwdt8LQxE5rq6jsHyJYQeAZvF68SnSE1jBitRhGrqCfGmwVpb83MZLaqX85/DGAGSAEfRv3wsw27
zqyDCFxgJlgoDdyQfpTqYotuIwc9oY0UPqpYhHrMMj08ILSfGIVa1wKVTzeB8J2XTpyKWmdV/+F+
otOJrx8RDA7gJYG48vAXYKEsdYc0kWiYWDsNW0N6Wtd4qxAxF4xN7DR/y7KhFhXL915BrYBH6bBm
sJRsK+ECVw/iOQnVadht5Sgc2n43//urgVVHcVAHWkorC09w2g04W3qo3elc/1vA0/KWFAdSMLcv
D/v59zL0rtPFdB++QlIm2ger3dl5xC20osdx1e1yIku6h8rRfKI2qaMR4IPb5LX2c6rGkKiJyGn3
C5vp3U9IPU+CPf9dwjle5hVwsDTrh3eVZL8PfhWLAVTjcjS57htejMJPZdJUJBapGnFBI7ef/8k2
QOmMSovvH+jCozieN9S/lPkD1hxJzu0QxJf8lZ+5QLrVhCRMUZLlgyl6Fo8rgCEW1XHpDSSf7X8E
r3oYPGlhaRkqiZWueNGGNLwa6JxofUUcdcWrzJpoDkUK5AwXmw+pvKz40Q0QT10n2+oFq3BjytX7
gYSKpCiidSPZA5B9ygT47jtfH/z6H3jN+xdhDQDkQr65+G7XxT29KcbBqS/i/4C1dPmiZKTC0Aua
dEHjKd+v9rRUtyuX109y4HwmUfsjPw8BMhvZQ8mSsSroS9T4zADZlXZKxXuYpXUGhNgQ//9VMcI/
WKo4guGtThdvsFoiWyEXiqhbBuGHrmA0THwIIMmKgI02W8ZcR6IC2RqYaSVs5yvgrbiXRy+NDHKm
nPZrjrcmJOweTM99VlYjmFB/DiE1iQXpaTXrrUyBTFhIg5O+VZ+xZfPkAXaqnileCBX4t0sQq4nH
7GwauJ6/z0iHH7eNc/OTH+TfWF5Fx9o1Hun/I0cxfIV5dmXSOrfvKR5xZ3QaIMGh7PYL3Wa6qAxG
1fh8iIQt7sjTvH+bmMn1udvKAygPa6YsSMB9fdHCwqNRkin0XJWKUU+lTIQ5z2eAAnTFJ9P9zNQR
9oUBo2hUERXFTKdxk385B4kHD+adPe0nwEAmnwiOQPB5T57be/BkBuMVWARWGuc5ReKdR2x4XjX9
Ml2+EW4S1hJs6QRQTg87EIrbZPu4EouHAjbSFMG9pO1vzNG1W+jBsesv4Vr3QmT4L+mZ8JWHD7+a
hXmmhs1W/ygrJ2jydbTabszBLFFat2kT9dRA8ZgjgDTCcdGZFbs9ggphbEOu1j+noRey0g0CvTtN
7S/WeU5Wf2bp6krGJ/31eZWx4TfO4hmeXSgTLV2ghHH65lynXoTCpzGIkEON133zTUYjJFJKONjz
jiJYX1ugNtyExpUzUNpvemLLY28cwmmz3DdD933m22NNovlPGMfPgr4ytDmFHsby1/14pRTEn4hs
n0sLHm04Sa7qTjDsQj3HmvfMEldRIx2XBA+7+xBiscaQou7E85gHHunIcns5qt4ba6kM64AanlbZ
u9KINeJAee/RfarzNYUo1T3MSHXOX8WeWxghlg6oqI8cvrW4ZE4E3J5UivUxmZCV3QdNfc1ui7Aw
iwrVHkcp01hGM6pBe0u+3TQqbX8Hxgrl3dGQi4djC1INKHNmmJegUGwPHgLhqdoA+Si9OmIEkKJn
iueDVDiFpjMQj+ks7tHCQjouqEJvLFOJoilGxcbSfx71Qld8viqOOeF0DD5p+1yTO8EGyJ7Bxb69
rpGoRaG6uzIcLfRylHhoB7cei6EAPLmlLgViJ9PO5EnoGQpl9VDBNI+O7hjMhvEsfw9Q6yt5lDnQ
sQa2p4fsplTC2cTd242De9g1P7kl48g1s+spBe1XyEnO/1Cty0PXTBZPvJyKysMVZLM2M9pJCnnX
afZj9D5YqZzwq1oets2dsW01OZ/FbFZ325fAj0V4yJjDDsaFF1iveqBOqmQ5uhPr4F1VYsc3tbsd
fI9R1HMCQwPYscE9p47f76hNZQrrMLClOKs9iu8g7jrs3sZcEuBxWZpWoHiQNcm63waozW+8UXam
bxQaskaML/Z2VnMEzjLwGhtTeyaCkQqGIZhKoC598qxPqt0l1Bb6Un5/GBtDF9byZWjhfdihj4Im
zevFZCAWxQtJAZxYDECUXNvwxMq5wM/PeWS+KPW7x+Ytbunkw2qnW9A/HdlgB15fXYkspAQnVtnQ
FBCfCytUXgwULGzGWURoxD+kq2oHoX786dtfFHXcGIgviFYVXr8/DrvH2LFYYU5jI4ofgVCoJNt2
cqPmwtydnz8u0tqIPw76aLso32ouNeSA9zIUTrKWlpvoEJ8IagG7NIVZGnpedRXnBFoYAU/cVMcq
N7z8JNdU6fT3/vTiT9SJ5w5zeuaC0InyZRcpFjMrgH8D5ynmSGLV5VVe0sTnole0wXxGug5YY5lt
pje3CIaCPr7Vg/aEdJWkurgljWkPq9G6rYiosIQTorzJJxqzx2BY7YKd2KL/R9Ht/g7tO6NuT1LB
w51XEy1+2W6R7g1h7TlhjD3hCfiS2YsrJUSEauDByVUnKZT728u3kiBiHdXu7DzXVSFSLrX1Uojl
yUtepekZnrxuC1ltgoGLMhkOefaoFPUqbkjhvvIN5TfxGJyJmeGaHd9XSeQa4vpsgHnEdTBHc20j
GIJuBrAEVepr7ysBr8hM6Esjtr9mqKcsETGoEKx9g1mlcOcw7NInRlhQhzOBpmO/bgrPzZQOM6ho
Pj9pHwEMubgyPXQl0CdJ/MOpvW/vpvSKIoBvfb82qG58nYBpf5T6x5a6f7XDUtHuhwhPXNFXNSnC
luVfCSRPP615U7lgyjhHj0oQxm7dkndZls8PdPNGQZIlZ/Inn4cNSPf8pMOyGL12ddxHAo8BYWA2
D6xDh68Dmr7F7mwp/9b8PKHTnDdMXDGYu6S/FrDTXSGCrYPMOogYxBSRvMGvxp3qbSGm2STQQrMO
SOfk195z1aWPlcd0787FR1jJiO9kkYDU4UV8x35tgOWQ+ifewXIbk5LDvPE5XIuYDE5pp20oL8so
ZWzwgQ+eqAjGKzHpOL9dATlvPwHSyRKhOQ4B3YAVmW2kRRVouEHkS4VpjotpzrSu1XGfCa/FGbC3
CKYUR3wS8UaWSOOKF4hifm3kol5D/HaYyvWSXlwpxANvcrLs6vsxURkOzviSS4Sgnn5QeSdaOjQf
Fa9e86eVioKtcqXzZXI/K08/rD/H845Qm8hrxgFiv6FdxhrBCQUYMZ3vv7ZpIyQCGzHboRakKO8H
d0g+gY11p//ZAhACQYwLeZ2MWfttADC1ZVgtTf41IlGb8koO2voYMLndQgLy+P6TcT6pjC8VwkgS
mkwzOV4tSoUk7S0JkV/J/hQlZ064tEGdjkkuuM0tFjBUbhFYOHXVxH15c0Ee1SqCwzOuqaiTwfIL
A1u0t88MW4ORg1rQ4ZY3IRBS1fW4JsfyJAQD3USRD/yB09rvKeI7faHjop/ERdZDrWWIBEmf6/rW
hw6KSHZ2IHa3uRCfq9s0xU++jyoSt5tCS5OR0kapJXkMCJBqZkWdBkgzYC9OZhy9jkwzfmsTCgah
X/CowazMdLaR8b1nhgg/ir+4Iw5ZHXAkKNRWw7a4ZL++h8m/rbWcbEc3RfGcIbrO2osVlARIEv7D
RUxUdXeNBYo+rm1Xz8VE4DvsqhUyOXoi4VQeGeZLoqSNqoQFrRpWqchPhfmwST6Vbt9tZ3mHCYYZ
vfPIbNHDCbEw4QDiPdepnTiI87BGCOhXA13WbTZ1fEf6hUSYMccCNDnailvszaW7wLL7BSMT0Li/
J7erNlSJ1EhoSGcNQ8yWjqq1XqFPnWUlwPuZqAnllxWh4TpUx9IAzemXnb7hhibWA8hvh35Ok88q
iyrXjZ7LZ/h2rq9e/y6IiLsJ47k3pRNJ4HxPFgoFgPfAGR2Oz7/xPYbCJ5BH+JB0UN37KMVJsEg3
8vQ4154BpaawgfKr3t201irX7yGoGMOV7d4t3h1c+l0nxXKwKi7d8SMs+ocCZtz3VkbNaphKiRmI
4oOyXVUsRwDGjzDghJAMGTIgECJD8/6VzzjdaBR7943BrmgNb7/LbFNvyExH1dfmXxDPzr1SlLwA
ILPJq6CZ1+U5mSBxP57lv2tqa9C3kNXrjDK1pDW/xjlq6z34y2Tf2oqrWX8mcVZnYGMLFD1W5hL9
DvAut04PXPNxIaIZFUNivH1gyTi2acyLcGg4Ww9/8HQ6nUQZhP7+yLzvBCcnI3HrFCHJhDQElU7E
0seMUYd4GSs6/q1V+L3bFK3SThYq8lKIzZ/cczxrNzVSge6kYoYRmdr+OYcC+bq9/aVJFlOSHM3P
vGjnqbV18kbJBjCpnXGjuyls8CSXXToB31BJcnbQ6yZ6Mjt6B4QhFWVMenkGpHa+/DfzORIuZy4v
g/KDjkaOc5hZnFroyrZ1Sm/vwOmohS3LCZ5liBQ53EDixel1jmQ4oL7aS6RWhH2Gm61QxH0sX3x2
kQE9wZoVnF3ndkoWXOMeY7aNImWAclgleX5TLcd6oZREVZHhh/lYi1RpGZihMUkvwjobfNkJhS2t
ZcQ1ntGteS2HInJV4Fjc6DcPNez0vHzOG39BDdVEn4SOdISAKDxCYHy9GnCYuAqpaH2mGiPGquol
ZQ4v+8sJoJMT1+ka6dkuWQvCml5o5Rkb6XWlHmzO1xNIWbYY/zYHmkDDaLdvvl5DR63SCon8l5SE
xkzFT4jRKVek9/hHh+Bh+JRAiqAOwQKADBMoE3AKQmcvK9bvaFEHldyTZGzrNu2+bfbxJixLaA2W
mC5pghcfL8UwdGirqm81wb59wwpV6C43/L9gRfFzDDwix/EprojqGaGZqU4aCy6QsPYEM32XwVUJ
2xWAO+uQN55ZSdnHlqDROlBBSYihlnTDV/rkUy8cS0S1wJeJkm25GZ5voUpD5xM/RFUqr8MzqVGn
RjHfPTcS2z/koDrojPhwYE77Ic1qY91sVb0YW16+nssfslamX4C+Qi0JT8rM7QNNizsEtdlOWVWB
gebM6FajS0y9d5u/jl25J3CZh1rCVmO0Dsvk0xlfiZfDeVXWVevloE4C+czhLyb3mu3pBe0/MBd9
p2j+4WRuUylPfhaRXYL4haWnkyYU8ebJtR/Vk6CCS6EZUJ8BzH0AgEzMczNQ9djVWQk++/TNsBt4
fn20QrlUT+A/7k4gyvhWFxe6s5uhLwaKWSP7xOZ2dcySD1klNhYZpPQvff0jUzABMWSgdDX72C5+
nU9iE+3KHe72w/1c9auOcdSCoQO8FudnHwKzp7r8Ssgosl8cwcX+sGr+4uUoV9MK0ipxcKDO5Fu5
agkWdWajlMMFZZgGSop49m5PqSViHIrjJ7vjqHyktJZ9GQUaF2zUfF+zupRXOYu8IR0FG381I5AE
VahwYQzAorE9Gbv9f86jpj1w32T1KKfNfY6O8EPGe7PPoT3J85mEljP326Lu/fPH141EQPP3WLtQ
I9MW/LLb1/oMn/6+XiLaJ5nvfDHsuaSYL+4Nh0Kf/6ZQ2/mCjcGjZrJ1meLCopo7eBRvfG822edO
j9EyHBEnwrcrI9dQylEQ6a3aEmyfqkGcGA0zucTS4WRdZ9GIGjq2PaYyafCVl5WL8K47XgbtMdO9
WmgQ59CQm3GZYpPZi8xmExXb8/5aGTOFHSMiLphGFPoestN6fKMIdvbCKD8QQzZzeh4MC9GBV1jB
uzZhHqbjxAbMl5X2Bjkq26u4rzybDlweTLpaWcNDZU6piLpBig2AhzSiwlhB1QxWcDS2ylHajkfD
3lX/mXzOM4g58uSJmbF6rm0mLDBPLKcNHuYvC0XWvgAJ7ySD4RByogec0zOvySC9i34x9HPAUyEW
5YdasBF9X98IE4psCvlLGZ2h6CKhxE4twjDzc+f0G2I5wPsZZSVDKongSUUHzFS7yMBs6NfxrjnW
v5GIZP1z7SX+KYMSPCMbTd5CPrFfH9daDV4rm4z80rM+OB7cE+CgJT1xoOfCo0/uZC6SInCmvyo3
qURbLRRRSnRIllc8TiFdqlGQTbAloWuJaXD8i2pGy42YnZlkYoAtcd3R+HAbr0boZpIm52sQ0L7/
pNcU5IKwCbm8DgJMX8PBZEpmM4cK4AopI90z099KV67SJyzsQNoM/9H3TPwqMfDSwI3eosKy78OG
/ARuRkJYvfQ8V08MjcAQaoUxv3sn0S6726Lp+M8j2JU+0kmsO2sGfbungDPm+LaToAGlb+NAYbHV
HNwab8t9M6jYX3QLHKVHx6N1sLkzhZY2OlE8ftxL/EVQVyQTlOqpAmTrYTJEg97R/RsfzD2ua484
T/5HC9BOLYw8glT2FeV10hXAl92TIA8LvUGF4Heg+mpV264/bu4exKIghx6vc80WFwNHaJBqF5h2
7ioBqbMmj8KYL5dsBCtXt4ILe6xdSgQXaTriEMra86dWk8kHDl8K4IVVkNfrCOIKL3CSI1E9jwrh
r+3B4uAZBuo2KqwXSApPdMQ6Kpk/kPrQN69KU4Gnea1Dz9lmqyCr1u4FNFZLxLD1ifcwSUjOvZe2
gU5ec+eyozwQ3AAC1uFv47rW3UZU6cdeW33C6OZ2H5fMBwFTinoxR2XkDrkx5tpwvZJkd3IewvNf
BlK8RbCJ467eMdIbM+jqUvnNQsJFf76+eHjRKcki1qdJQfDQu918H0DJ0wcuPcGlg2Fr6eosbT1w
bWegnoJ1iM2elkkvXRJUZe7HOi3XxoLBsgO2APCAKxTCMFm8NRSr8GtfliUTA9W634iB8DtIl3gk
CuJWUfdZKFTesRSRreRJJsk8EaREnoXDh8mWizqqMnqRZtulO5S6HPzXnddSHeHwsYo3gv4GbG4f
MhcAskfkgBJYvo9x4trCUdZ1Lxpn0gK+18LVNOB6xMucwfeaSaH2p8r8g7HtQYj7AsejHYHCzYcg
IV8oHR64md3mXgsP1MOTzOXb7EdOx3C3Zsi5nTJVpiI05cIXHeEizLSP85pLxlxGnib6dwR4sS5w
Yt71/4/mzeMifwC9vhpRGKZ4NaitGxGZE9jXV8tBwgyTgdQlvn5VLUjKZNuvYODLdjGKM4zjyDcp
bB89495CmDkajUNNE9vh4tDLN39IvOcXeC+OhnHB0PA9UOuceW8rxy4ZJpdVT4Jk/MM3apuEl54+
GmakFkTDi9tdquA9gbjexdiO0xzjptCXEUSVlYrD6nOzyFulGySe/5PK7zJhNKELHhWDo4+bKjs3
SHgR5vOPqTFpyIhtXSUTZv80oXIwKpud+lCxnJSnhZa9vGldozQXUNJr1q/T80J/VJ1aX8E0yY3b
FwfbOn9YW8/x4vzoAK7uYGZR+wp7TEoUKPJLYEnDWOegisUPOzaisCL+RHceJHMkdOsUQ0rO3H68
vYZn34qf3iHBGlqTrFQQtlhR8LxTGyjRvjwGXGx0bnbTrkcfB359MHmQCNLGTEtX8Gk3kxl8aCSl
gmshCaSVDNvU5Ruz4f6wTnGn7xDVvekR+ZdFt3ff0cozNGApu3vMHMduvK73xhZ7EiQ3/2VKSx3z
aXx3VW/LHwVRlkEvaZNI/5uqkInjaHTv7rglLWnvt6k3TvPSCUS99QFDS1SHVXbXUuJ5Tiz3E1aa
F9zTOElEzj6sz01RHFH+o6Kk4FXotWAqSWSKpIZHqVwOoBD89vkdOtmodCjvWH3WpUn2oF+dFKHs
KLv+oppUXurdCCVv895ePAS8r+roXmCnjRh/Ukcg1BAKRFor0gENRfN8/so9xrKdgPdtt4Lhd/FL
AF8pbm8u3y9OtnnU75UW1W5BglfWJyTr1q0qGLmlYEIl+p5Kt3FqvMZCi4AmpBr/5ZtkHBLN+O/e
ZrSyMqbRs/8i4XlZl33bQvsg8rmG6Y9zFYnu6atZXLZktBlAac7/BDV34g/kTouo1esPtPFk1vi3
05L/j6W93CnhoMaZq+8XGzj631Oycw99sj3uJi5HEiB9kHTXwUT+3NZ4aNE0XUwU43Ks2M39hvL+
UR2kfbgsE//5AloKaqAT1RhwRNIBhJ4uungtDWcC4snd3dJy9b5x9rrLESQYCuTK0EaQsxkmmuVz
cwJQqBlTGF65M1EvnWMYiJELgl/jGQHh8IXbYiAWgHkv33juCEt8+gSCLHcUz0bhnJ8RaBSoxmN7
l9sCP1eRXFk1k9eOz0RzWEMPWJ5CA2Lzdgm6TMuwEM7/9TVLmB1T1KWJvmTnBLq72ds7VrWPLGnH
95/z8wfF9BY5VOn9z94EaBtpe4vBb6ZCrjz9ueHOrRjvihySO9X5j+RqoYmH3Fllr1yCRp3U4rxS
LWtWs/pFPKCasdppHEHPFp2oiRr5PrQsteDTOnpaAhx+wkpsoxcVUx3jV00myZYWNDnj57xqWYtp
CqAxhS56wauqaJKB3SArfnpIjWzP1cVyAN+WFE7yezF2/lHgDiy4BREs/8Fz2Q2orEa6ZU99RyZx
oM9RxAkU5X8kKvDbbs/+2FR0skRUHZ+XuEzPHLDaoL8cDuLZS/1ms97IWqvQMgnYLlFiiWz+NB0C
Uqc0677cUAsy8v+CqT4pnJ9W8OVE5nY8/FOMGhK0NULkxq49mqttbDyjtCLShqd9wyJMKi75hYye
2yXOA0o6ttnnWNJTkpMPqrvSm1Ri7LwcRBydOlGCfA+0iGRgnF7ijzGN2dYdSGPhO8rDFmplVv3B
2KterqVnyJOw98494A/tNVAA1QZEAFUHOa+/FUcispsl1EuEDlFZcmbsL/buZ38mRqf9vjX9popb
b+Qd5IERLif57tWOqJkpES+gnKPlx1RWgIvFS0ozGpJYBuHaKK7DU1P4ojp1J65trPM2exHCEKdQ
WyoUAusn5wXcbDJbK56UEpIdOOw+tYy1IXlVf6dq3iuB1Sus9zHrZlIGiC6rHtcBNDSXw+pkV+JC
TRMkmEK10dUoirgm+5EHzamwxO23Frkr1SiOZmKdC2oxvMrHLB60ALySdt9PQ2LJ+ngmdZglCSd4
dbvHdcAjlISN7lfhve8/5BmRtYyZYbR/PL5mkNJXLRHLEBGqZuvYK3jcmRm5zLzwfEjGhh3xX6rL
lLPKCPc48aJB1WmSSGA5ex2X/pVNp5+lwPQ4/BiG2y6nGQ/0akS/lGQrOYACoOxYpx4TBCtfxs97
OStB29CShuwXNb4qO/8uP/pWUOBPE0Edkzp8JaTS/HvqcsdMgEn9oeFAPh4PiXT8zpYrAyxWUVGo
KLpTQUv7iQiGPukg6YcU4I8dDtwouHkskZdxMc/ScMvyMsBvL+6DYMX0NPKWUwyKnQn3OlO4Uz0O
X9KoEiwc3uMsiDWbBjfmRbuzw054dm0gk5RP0tDGpFHinetWz1dfH2NpBjHPoPvPI07TwRWfV37K
ks/+tW1YtddGTOe4HWYOlXmJsJOeJua6euNl9aS2PK0JCYlu6Grs6vzmrpxziTUQ6bgNQN2lvWAW
jtgZ5DNeNSM5I+IH69+06o1LENJgnhhSw4Vvu5Az9isvyezQt3TDiIMYYTg9OT1kTgC5OcwUdy8D
3/BDZBPc1Yy+MdlRkz+QYDBTzZ6Sy5sowzkni0lXrXuln3cTk8rQMeCxhe3CFDJGjEK/X+u07fk9
wS0QVmUVdMt/gOmIYZY5ZjKpAmVbkcjtgkkrYA3+WbhxQQmm3pcL4JwqfTXWxqeKaJfMPmw+wCF5
Ep3U2cP56dJh7Wj+QYml3tOo7kqjis8hI+pSKlsHwRrHx61Z0lTGo6VU7DEjbmL1501Jylbdb68b
G9CvqiNw27oR6AIn/YIyA8n5txMLPPOE7wlE/PIy0PpQUFHOxeNI0b8Lk0CjfcYKJt0BBcrN8q8r
v+7SoKkq17YAN4BQ2dWavkwEy1KGaLIh51rAC3J4CHPEJKZiWyOAbIy7WZCGpjxaR61aGrXIdb6/
TLT8rhZpF6vOLDxD+6OmpBI9glymaN4o1KRzSBHNSnrJxe6SbxKUxGMM9FsvHNwe9UV5R6Qf3PSR
KfcmzmQM9Y9vtniTPR7fJPoqGMlQA08eXEtGandz3dkANHUR5J4CrSJU1kc9UP0R9c3Prq1if3wD
88v6Gxph9v6Iwr2CDQwIsqU7xixU/uDQZKw/xjxz7F15qayMEuWql/qnAGIlmaFF/AYs69S0jrpj
wbHA0PRyLigqfHao351gQDMiMKA0T7Bas4odnDz1qCys+e3KXBYNaUzPaVUCfcENtv7F4UluXZi1
kEFwuRaPQ7zW10hbIbDfc6T3GAKvJhTepkLnRQX+ayT6+0oXCMG/MkrNzs5dqwVlMaBRdgZErAWk
sna/THA4zXk4HRhkai0sQbKcWDidkBbW2SADhkulkU8/2ZSid6UIvp1utTfO8zfMH85laC9Ih+jl
ahv+H7AHlqMc9HjR1lc+2j3ROD50+U1muIlIgKjD2I8nqSaCRdB8cdDHg6TZW1Xd0UuH4IGuvEUZ
p64WmvZXNAC6Rs2xAp/XDppc/PxywuCxjq0OojZUV04bXjepmsoXOnDj6XIMweT/EGqfGeXeinxM
4hMlo4vzhKUg6Vbhsza/TtJeYZBo998MthZbcYBx2XSzjOFcDfaO5ONOOS8K8LYGu0xugXjPx2PE
M8EV0fTydCvNSfsPBBm6cmv0nLsByHgvZQ+ag1vJJEMFgbZLq1a7e/4lN6oCJg/rnXjZO60OC118
Og099N1jzeGmvtBoLhywGaoK4LDXgpV6cNipMiuV/HrBjkT+iJsOuGnGxn0Wh0bu53gV158afXJT
lBDxH/1QhUOY/fneBtt4/1+rcjNJJJZTzAZSYOVGPP1W11KYIhI+ESuIEoDyu+LSEYu/LGJhqlVe
T9yQIWICb1X31BD/qW/xFiAtjxYPEGOdq2eIDsknhWzZ0rFBBBIzQ8JsjUwc9dX/h5TmpX7WPe5o
zhMemwwudkSDjXRNsfYhKNUY/iCYVH4ZXxXFR4hHkdiQp0wRkSkUR0tNm8C6WiKDQ8wKvQp8CKfO
OyPjv4rEVtjHzFpFZAUwW+jp4I3wNfhF47lkKiK6iYUGyw99pf3YgOV4rnQ0h9LvQd5CAFv08dSa
cjmAlL+hw5+3pcV8UhanBT24mDiO7Y1PCo0jKzKpcCBgppKhMNFFvw9VuXB4og2rExFwGvdZWVwo
LE4e38VsnSpFkoS02PH4XEWIhHQrvJ1/vfEqRhEezBZQ40NjbRdwqig7ftqSHLvL0v4G8pnhTrpV
lIu2hdRd/zs8ZlNYmr+GikkRiznW3+eut094aUAy614jTSj/RwnoRghKINui5RhWQ/MZKK3akns2
DyPhLd0+QAI+DlIWEHrJh9qA4tX0wb7Q/oIGqae22Fm9LOVhSInITbCgQwyWsy38eRjXEUi20gPZ
H6ksjWtc+y1AWrI7GvMXJtoatmc7uoB7JPX2z9FgQzdzkfBAfQqHIqJMfGzx25yUkiOD6Y9xyGZ8
1Ix0+XDESKBzPhysjucEik1SMQHyEC3qUs8aFsW1+UX6VbyVjaM/CGQmcgKHO7ybVH1Ky1gEFp3t
1zDkXekerFzJVCiQtrETAUq1RwBddoJUWTUIlltX37Q4cfC4nX8vy3QRh4vQKuZ2onPQq5YHwus3
BSTbloMapWaMipYRw9LjrnzRXMGgF6W0OoHDeUTEtCS0vHiqVvxT0BazaWk29nuBHCxU+2Yl37gJ
1cImyfTCq5FgYRSKntgDQLQFtKEG/jQTpfMUrX8mnNinnmM73OamPgjIHuax5UHN0pSQIjU2blG5
O2hvJU3olMMQ7jXpsKgTvwC4KwvxnH3p1/UbcbFcqNWAn4TP9A9FN9saxaTqI81mVAeVvHGVR25W
2ApBUCJHiOpSie41qmuCr2LWWwLSyDCnwWc6exBGbGcKJ2yC6AYzmxjTQO8EVhw/nykWjZJr2ERg
PgmTHfMkAc7jF9h7NVABqPk8HGSfMbHEPiEkNNIm87uv5UBjtrJSiED7e3UZOb5WEclP3k5HaWDy
xN0paWXGud+mJfStX8zUGOqnrsW+ypUi2frlZEVJOrwJOTCbwTMBNaVjSIISYhLOlyc5aeNvHDlS
s+PinPKwluvTX8S34V8/HhRPr06JLYiUKmPsjFBDYM2jfbKSisIqyoo8KuPKqv7syI4wgXFk27h5
CzkL3qLoj3XsVSl1GhoO+0cQqVPCVBS46p8HRFkDRUjs3RM3PAumZZW0qWQtj3BhEPnn4IhkT7Hx
qARY+/SXaJdxy9lzxIWhxMjnR2iksJFzRllKEsswXWQLTvtl72jEZdXsT64hT7LA+R7UZUJSmsoM
oruzdDph+dGb7WKbftJIUs+j81ocRrDmesCkiVOjPwYvbeBOM+yt7X+Gt5o8kcPwsrl/mNMoBf6m
mLPxwclvZruqVNogVFX+a0timbXzVQpyJDRJPupU9U47BUUQcg8Kp7irFfolY508qvBScY1XC5QD
cFiCtaRQ2YTvbeGuWSHzGr+RvePQxmPLDiCQufm/pr8cWZToWljyVWykLNIsvBp+YG+tMqrrxJd5
TExTLf251+oZaYAcgI20753/zwtQ0zDre/9ZmK0k1ItYECYqX7U69A3ePA7LTF36i0aTOqQpZ0bz
PSD4BVQruh3yuugpWrRu6vxtvvbmeU1I1hQmglbULBvlISEs1hPLldn4692MaceAIE0tIX6HLOQD
fYniFT0DhM9I5QoocSFFBs1MSvzmHag+S5i9FCOsoHxvrfWtmeQZ6rxl6ntdIMBUkjSheQ2EZyS7
q/EiKZf80lbNE1twb77qt3I/Cntn4yj7XkOeePQrsJ821cjVM6YLEy7ltrakNfL1xmL3cTa6Tv3+
DQBZR07n2oHE0i1aNv0A+IA2/06UAYNPGGb+xrnjzTOpxf89PG6jnByshcv5rjFzDX/Y4YBBEFE1
vYvtOHLVn+cOOzwDRPJsCdJcMHOYPQRAUzlh7ded3gWY//cclWEpdXQdpZKCTMp2cUq2oWhIxsvW
gLW744wyFMzQbQqg8tpOuGIqNJL7GzKvqCMXzPjk/+CfbEU98svidRRn3ZkOrTXJ3wMA3qkjoQxh
UhARlREmzxPUSfAYZ9Jpr20eCC6xMNQh4L4wKIun3uilFoG3LAhPIEUSTrGxS13bQX4rEeWvG62Y
0AxQxJSNJjLTSpamQIkWHmD9rQQoZp9joGrnohte+tXbzwlQD+PRz+CNfRJ7g7kz6s54mRawzUho
0Dz6L9ln+xXwNQujYLLmTZ8v3ggSX5lOEDuhwwXfjf2d8ekJxdN2yxRxkJQ645KSsQ8bkkm4KVLQ
Fz8scBQQHXc8hFrEEloNVBDtJQZY2No2kRQSuK2ms1XW9aWEFak7RunlBg0fUBcsclg8lMzbknlB
9cuiz9NuAxF83S2nfhWTgvHWSDDED6vOcW9ASkVSXoggmvRSqqDcdvGPSD19khukjjgxVFSP3Jma
R9CJnwRBcBqDCNvNamcL/3RmVl8/mh8Rj13HsYCE8R5d1mtdn/PqEmCZcMNDk+BaiSjVoghwYgMU
20Pa/jDCkFkzGWfLbV6oQmNES/xnRk91bo7mktxGOypP9v7rD1db/wOTRRX5e+gxywWJmaY2PHel
Q1PIFqLyczFpdv0Q4CVBeRVQ648YU1hN0FSzNACX8XmRvwqSR0Sgb+ei/k7eVmF35Djt3vf/wAET
1M+Si7R9zxGbJqCgCUpCbR09PG9rVNcDIfhp94fyJLkQ4Dh/SGceiQGSme7Ck759T1IPFUySsBhW
LR/8biJ2W9RVNpl3H3bQR4PeWIrSLQ9VUxAQe9aUMnAKEVgnz6EdU7luI5salUlcw6QSyXqP16dx
6Y04FDKW2Em2BEqDTq6IAURCX3OSetyCcW77Et1mJv459FZrKPQeqw/i5zc46mE4JosQfh849pcs
hZRji8OEThwY2yK//jXG2QFmvvBjTTgrT/+kJIgcEtMdo/f9doXENL9+rcfNnijYMDMSuf0cjGbs
HykbBcFkSV26eopz+WsiXKxxUqpl4upnJ09mGTaUDK6bJj2DjdjKdaQD5DCx4cj5g3tft94jo14E
PGQF9O/HVgc7lMM+hE67LXNeQ+GvsCYBv1s76MlXiI48ixK0ymK5VspzlPEy7IxgSR6Dwx4nFvbX
EfaAqFtA0RmIjis46haABEUrRJKiA5koy0AvS9ZIGnNVZHOZv0NkTI/dNUq/3oBF1UUzXlI1t3nX
YakfmFlDO710EpYekXuJ0FBu4i4RTrkECEAI605mHYI3EAqMMP9OaHUb80rEpbLH+7D7eCKtDjSh
09AYkird5kB7OQpf+L6Mi34cl/zse4xQKSTAteRwMwjcWxNR3YZEEzfJKNBQqosj2qV/NjtTDI4M
Uwg8u1fGyRxUgMCiAv7devitEt2KggQmq54lx+GfePa9Izu2j4THKqJjr8v+aUhkENyZx43TkRAx
2FSYojyn8g8HfRRHdUNnGcOrNAQBdTn5Q/cOYWcVxH0H/T4gnoWP4rGEENr0GhFshIGjQKeulrS9
rkaBLB0hWzv6WM+sEJunrZZOO4fxBETY7sgIdFEm5mk5X4XXF4kPNiKy/xA+/3xC6t2P/Ws2s3zI
x0SAZCWdZXXHPED6/JXYwx9piiIU3MhEndueN9P4y/Sz9qAGdPnem3APJHoNJyx8Io0zJa1B0ZOD
jqHzQ0Bgsx+KFhmy+atJNH8U+MVEX2rs8CYHoDjlTCylLxtxU92UAM/y3IDQu8UE7MgYHtw5nsfB
kZB3Y0/QqWGeV4zqlK0tmGyvrNy0blBSeOQCsDNt0omhkHfs1gDVFuzhNZ4liUfWPfvu5Gplb/EE
iSZKpf4w07TE1jJYvvWS1SqyNPaykhm4Ezq0xN6ku/xb74b6B39G67HrmLLP1LmHfqjqhhvPQJpy
SDYhgEuNm7VPAPdOiwH7WIu+EcVf7woy4vmVKs8yV5WcQ0K0ZN/vihpw0N0sgsKoDAfCju5PbHM1
PgtJlZZKs+ndVCuVk/xmy6hjK8NgC0xpcqpXq+9TaSH3npCjFU6SXoSW9jRgIVYctdXtIEp6uTVm
UceQVUyW38bcL9FcMG1ChnRi3Zfh/jHa0X8wweX9Sfz9LDPjmOsNvt7vDGz+GOX9RbWCncqDF9U9
qbYSfWp/cfgmmTYJBzVGJDELoGgdRuFgMBLLtbxESa4UWfTGVgnx1YHH2y5yuIsmElkSXMLzU304
8Ux2rXqbBWaIZ1/iv53H8FoUWNSPohE82Jnmce3wzKoZXX+MYIejpXyZFtblMTglIOM+0DDlmJl8
sIcChOZQtQdpwzLlu2zCPYnN6FtcdWu+sJYY/dLZ/nlSpxL3VEAL7ncoEHhVcPnpv3uKDE8zQFi7
nbappkCwMeZhsdIfaDtuGrWio9BOg0NS9HXI+NQc5lPSuxk878keVUFwm0dWgAQ+0X5Zbw8iKBGy
QSNvRp3A4pBPcp0PCOBij6pBjyoD9x9riSTgMV7eKCnWlb/BXQ2vjbfVmOMZRTLsIwmoFFsC/l/M
mGYMjg/Af/eobJ4KLQOsXFu38hDtRHjQSR4+UGHyefLrz/hWvm3eTlZenEth+EBzUJh2rwJIzPQC
m5ej2RQkgFzPc74iitoQFIaoSao20+Ur+SxmAFU4hYM4nYFIaWiTmmZZ2wKsgQkh4eu6T3jM4TAD
6dWpCw7yJgWOvpHIfFASox5R1qfolWFHF17h1cjLIsH6OjW9sOO+JytAtE7RonfQ2ER1iuJ/C1vJ
zZiqL8/xtdUX6w7HE7YngVGSjK+K/JrUkqHE4ZeFwCGx9V+GMQCBCX3Es85UPt2qASSPEUC014nc
8ZTdrrDYwppiqQBVQ7jSLEulh9Wr+rxH3UKz7hoKjmjG73CTKuyrDoqcNLW87ol3v7LpRXIxU2sQ
8rRBYfgPhGIc4Ue6FdSOMkb6bXzMWnVA712CDAsKNDBEiZCoSBweABMJwpYpWH0N33KmJLF+4WvL
9RaXY70AXuFj3tGckR3MKwIXwTHl9JX3Zptxn1Le596CHPsR9FfIbPf6rVQLbkgzmZKJ//zXEoRL
7x/PPde9LqtVSC33qOt+eXtf24LWerX1Ern2Tz1SQ3ZX5lexqbStMXoOmxob3H565vwrbtCPQX1V
N+3Ik0eG56eKMMkglyenRgehktvdxdRyEhvO4jL0dBHyJDt+vsoOvJOKV7NAO2ZDD8YZW0C2wSZj
+4zcRFbXvvtYUP2dckpoYHWSyLdHbKaX8RsQAgGjRu2ra1k+6PXldZFufKdwoYGNT8xPulcO39KF
iPt8YvnNiTCKmRJPBxl+O2K1QL9MVVkgJfudJUlV535Ky6xbb+rZIxmZm3n8zFkIbupmtLO7idcx
C4js0GmK8S00ng5uL0Ng8eHJeVt3V7V0LBewOHgqTnaMhlhbMuijS634bOk66s5lP6W8WeuJSj7f
vrqQp3X60kqIFwWL/dIw73/tNlpGMKPUrJroGMWSYKvvucDm6BTLg6PmISuV84Xuxysesw1ZESy7
lovofEWMeZUWjsXlpy9f3hR62tYzQxKTTt/vXBNf2vQGl4L9lmTFc23LICU2f0PenXQebcnw39MW
hU0/1tyc0WP8P17NBr7ybpKR6xbWBRx4Gb+Fr014TfLneL3gpze2SmPC/DIo2RSfU231ADLoUDK3
VVZv+pTqEQTxrt+z2coYdH6IktivCeE+m00Cmxqoy/Hzuf0XFxuGufexGXwsXiUMDE777w54UlB2
VU/U1UhxHlmlltT3J5RzX01HCNV6k67iJIKH2mlxTAufpDXoXZxGTWCj+QOsNUPfuWWICLWrKlpM
EUmhHinOhwA+cbHOdVjCzVS1meyykUNY7FHx5QuuY16L6Os6/5PFtBuH0thWQxFgo5X19Euw+Mds
2h4O03v5JHLVIjA9vkf4Sjo9qBKVkyMhyIkwy8w/oufK87e8UlhsC3z3XwggDewU4DgxRjmHb55M
eljYkgev0fyjQ3LzORuqF0j2R6vBeA9ytJhpT939KMTim00acETMRzz7nqHcSXpJfe6Hs6TiF2a0
k5ldin0tPqYrWb9RXP0vZwWw/gF0awu1KW8Ics4QRLPGh3Nj9mnEcDQSuxEDKraWgONW6QC/Fylv
74d1twhJqa/BA98mX8c4YKTQy7fYkny1SwYAs/CriVca9cbtDJ33itu+flaC+Gs1U3PjAmM6KF+y
0qvV2wmVMZtjaJCBIekBNYRnc5pQHrUQV3YL0RhkQOVxvQkYtJdpYbLtIxRoC9Exoy1jran/v6B9
Zw+NMwl6/ZSH7pZzmv7iiaeg2ok6iWpe67nByC2Nba4A6NuPq90LJVpLGU476dQHvDM76nlPUGzG
AfJKyX/L035rFeBidj73qKSsmNYoIn6B0hF4AVhMsoeqQqzCthznC/QL0wZmajhQ6XAOgEc4i/AZ
4YG2LpwSOGpuI2G4RM8RiRCk/Iii6W3NzdmOKtgMImzSi1X1lm89ab3khTiQresVnSujYyZE//Hw
iFib9OnDIa191IqpTQW8Y1Mnb7t5r0mXtTDClgKp3kf/Il9mggbson8xfDg3Frv4mptVxRXX0rLQ
EoXd0ZOvYkk7cJDvWiHWKXeSUkSLhcvWoy2dK6QeU+z1tQHeE02ohKjVPiko+h/0sKX5qRApsuKV
ApDrD8ye2AgfcyEGLNkcDQUub5w7XqO898wkGCT42QCuGCIuh4O9J4yBYHomHtX39m/jHr9MnyHs
l27/LHicFmi1QY3KLkQ2M+Dy22QO/5ZhfczHSVzQL15TRGmoLpjc6nLK1Xowx3L4NPoUTt+x/Us3
lSdqQ90ROPbgeLAIl8Nt08IBQ3r6Pnblh8KQyoBLfpJowJDY4uIDBptRv5nFA0SztJlSfZVLnCt/
+BEBTg7AFXxUsfBsOW2gX7sw2G+45fzwhkf/yGbAxUSuYl832XsTKRCZUBjzYOXFw6mgoxCirgY5
tFJm8mXEjbG1Dxjy44L+FQo/TBBdqegn25cHvViuoNclevtELdGbm5yJALak4ox1d9ToiFYXHfJk
9Drd+JpnMbdatsQvOq/ByXGtvFTQ2T5YJyCLbLY/YJCZPXMbK7UddlRTmbjuvLyDbJM/YFVSxnf1
qzZyvPghdt0Tulx144AdCyZaUY0mlpN0Hsq7QQuHh6+LkWfF3LxQ2w3l9aWXzU5BaOxmzCB4Ici+
zYc2854FitGAJjvJnBLXd4/T1jpfvON180qILBH6bF6MuJkezEb8T0h4jw8uKYk+rtMxStWAgIVj
uADuRm3PAGX7UN1wNbwfp+CYYY1FI0qoSW5qBbqkyq6GFIZwSP7+3dlThcI4AvgSW+FrAFeyntwx
Zr0sLYCfJZp8DJZqC9DbZ5I7Ae+QVwD5w/nfBFdWy/cfs8jS5ivI1XCOY1F4riD2SroefxVuxHOu
ipGQiyQa6mBdO1HNCXXAJxuyEs76AOFIQawHpnzSOiskfri8UhEVWMFRJEW4tr00OoxTR7Ll0UmG
7CRTuq07VxnmwA+60VbnZFkQF+3SUAHsQ9AHCPSY05rOpEcWwVIlwTXAFUS8D/7x9gHYd59c5be4
ERQGnKdYUMIwanAiLqjtGbwtdvs3dBeXlYss5phf1pezLJJt5MAH0rTL0T/ChepWPfWSAOAojvyw
uZvCNV1OMiOWWaWTAsVfoW1CJqY8gBP3qNtQLvn3DxZtWnR4ODMmnNlQYSDuToS6LkS5rWZSolgN
aGunpcFr6nRHrw/uNLDpMnJpgkxIrKM5pZooiMLe0tiT6NXf8+65QUtN/53stRsGqw4X+hNQELOG
J/KMaBF4R0mteL0Ngqnh2kd2lU6JW1267ZfTu06wn3wGPcbI6slTjg+yKzYAvIkWVRlQbryWPuDY
lzb2TbYQqNhK8GAfzm/UZv/5mww1SL8kjkBi9igkdfC7zhFtB5NbD6VHmNI+1/r7FICDM4wxrQH8
8rdhF9tT8GPkT3uHNAkKoMRrZeLyjaMawLnuE9qiZPWgxBlFA5WeAzAQQ7tlWg0/VmXGqV650grG
Pi6cYJ1L4LkYIHLTXF1wLDwkuoXoOU+8+hlPtivw9s9Poui2poWxi3LtOLHwHssHjP7/Iq9d4II1
P4YSXKCJ43eomSZtXouLFxyU/pGi4c5ylH7Dk02+8eGDYkBxM1lo4ZlUE5l/ybxFtcx1hlacn0hn
MJG5oEOUGPhF6gXutEZ4Jaf2okY43Mgh2ytzuftxRD7F/FM1AILiuYTAFbKMxHiKc55rWVUz76ob
UEO9kzVExkTFvyhM/VomEhqN8pbj/7Nr4u5Xl0x5ycItjs/MSigu1oobfz1XrIDGuCei6K+hOibl
xfSWL1X+VIsLNL6F/h3AWwmXep6yt6psATLSDBMW8bQ7emwDxDuXpgEtE+l7eL8p7ix9kY7/Jtam
VY/JJYYNNVP457vFlX/QJ/yOYp+800uCNhf5L/5Ja2/sK7/H4UPwno51ZI5wjy5ZDkuTxLA8ZHd+
1Z//eX7s96s5HMlFKc2Pt8JpMZkasEieuoWRWJ+BDbFfzsMUZhIwHc1KAhzMJaBQi+4jryVLX74V
68DI6vt5Ivv+BtV7/tt7leaUrLuc0b9MOFWFFO2nWB3itp87zzpxJwaj5bkSuDsvhmcNzSLVPsUA
pBhwUL36hjgazCZBal/d/tknVpJFxZG36AfKBZ0t05jtuqTu7xpeyODproslsK9bfbL6VsXzmY8w
Orw+GdCncpx/z4Kgx3lhcqP+OazD88+M46ss+t8D9jlVyzxmzoCaMFwK3eSeP1v0MDBk+DmKWI4+
+RKo8Mlo15lFt8KjOXiA+k0Zm/JWdn2ARcb75Mmo+Yi+D85gBEK7w3EzueNV566W5+XrTnkfFwyn
EgLXPn8kOzmIEAXklqOgmedL3ZDLAp+YxqcOFjDmUXh5oS6qYYrSPulU69kIGuI+hDpH5UDfQ+fg
HOxeSA63/MiPxZwG7ijo7muQZukQE+cflmRYB2omPd8ZLp6hIquC5pp5A+SbYUGcuC03X1XP2kYK
CdDbEZnb0IzRNDanxAA504tqVtvjiaK4TBoCkwZ2RdpDqEoqMWyYVj0T6zssiObmIAbtyCiT7hxS
WTUypuIaRP6kJ9cMEBsq/aLeaN4mZEPWiR9ZKZt5LzLz5/J2w3rlGITAPXIgrBInSVnC4cHTe4Ia
r+uCr2yYed1zYWtmM3H/HwGaerGWKfUp+So9NSkE1pfM+2V1UHN6kAUOlBatTiOzb4CC+QyAlEL/
knTtIOOtCPtRCAFuPk9OdibsURI4FwWP/ZURpcGorVb3fEHz9u/hFpu1Pr/w1mJrPMWPDkt0/QQV
HWlo4mxlJbmralP6aOezM/LZTXT3/KxCtqYiZnuk9znkUHcAdZLnF4CHU1bC+V6tYojAq4d+Dci6
IKWUQ8biBGIWUovwC88vNulQJgoC/uFaGfUe1HGCdwftMPYVnuP0oCju8wMa+qy9ztBf7UVaJAOW
ltAx79naiVQIUcfyBceD5E2BjNpDEIltiBihp5DpU35NIy9F+M8hbjNvuL02PKUQF2tsqmvAbucI
hFLhs+5/r81/935jWWW3xocBtxfz0SvIKy970NsUXQKVBOi2cURN3U1/xP3CtTEpw/1GyTn8rbF+
ptwPAe+9iPho/E3SwPWfAJchB8KTB3wSZJXvNT8RSOZLCnilJKlhuzRNtcAMCKoW3sjEj33/anGU
xIqsTLFzZFJiLp78UBFelMJ2CHfk/rZJ0fo4J1AH7X16MKqwNzJGmoXTRkOfrZw8JrMYQYytdNbm
bupzTf3ZL3POcszEgXXrLLvkXOh6kYFM0LGumWKTx8G8T1BOLnhMCmXNhT14cB6Cs4bXsZnR1D80
Ypu6aQxA61R7Cc38uxlpuWrsM285/uzTlb2SpLycDAq+C8F/RQsxmbt2NiEgqMAPJS3jKU0/onDL
/VUDBiaPgQmToco9peqEeM1F7htKOUuqYiee7F4XnSlARR5RIPWiUmkEzkuLNTKsb/2xbaR37xL4
N5ZVODrH2aK+l01GKqv2XwPK70eRW5MhJBm4f6BJscAryC/cs2Tv0DGCV3dXqF4zEhY0KEw0b0Ua
6NVobJMHiStUEB141fReoyFEbODRcw7eqafKkqtXjkp3BcihJWaWOCYekoIcBiPjrX3Gtsd+WVpI
J41Ei5O20On7cRqvlTMntxSKJ9tV9DswLEaUqiEt1/L90McBWhmgFMGtreR/f4K/iiautW5dJ2ps
9aVjOOC2EdJn7pJnGvgR2oLyMcMP2Zm9cNccnxhmdFLaSHU2oC/c8ubr6/dSFNQK8aRKMclle8Uc
n+2/jYBEYxJkP5Xh33mj3QIzVR/kcxVX59v4NG8dPkVt0Dkoq4odXk8plB9sFUzCawArhRdvvaFy
LGi5nR8VFE1tq60Ly3x+cMr5LS5XeoaHvL8UwsQFiYmPlVrSb8bH545RF9nHknHahfpxILR017rV
P3mAKGmr1zb6xTpwE6yFCcA/e9MzKCRHliDMqUPOGulxHNv/n5t5OSdUkyWnH9+bn+Mtsnwh1SeC
o6R2Z3upAo4bqdqwQv06mewRXITHK4ynTw/uQ6N4mMmFaVZ4CMk9EBlygDENgHFnYGSdsNeTG1Fn
5xClfd9Ban2g0u7gftJbteRDaSHZ5U0FqTTfj1CTp0+xJbGsruaTTIcvh144JwMW5GnszNfCUegE
V4pH00lSq329tlBB13J1F8AT0q+P7lcM5XFtcEBK00wBhyWjtBacn7yGzPm3rXyqXAwZr6PTr1mx
Mij6xi37ksxcAB/Bk1UevEMqNUw8JFqsOhZfJ7/oZYGZQthiEWR1DWbmpbSCGF0/ZSC5Yo4DJ+2V
qbIhHTBYO6mPs7xGqwURlkXnncNHE1NuYKlB8yX0GLSCbKn4+2ORmkXD0gjZ4NjGrqhxA6OEW9Ig
1ieg3sj88Kucc5CpkpgwJHTLPz8J51W7c+rSs2xOxjqZdHYaIbzqfxYUA/wAjE+v0lRcrVfJcnCV
hCoACUJQzCGjr3F3huwtudHr8MKMken31PfXCFjrx2lkUur1JljThr8HnVHWvJ/XGMuAxSEJJbcE
hp33rVmaioDa++5yVcIMqxTCEdAJewzhK4XG3wuSdIkK91PUqKIGqS1miCO8S8pt2x/fMgbMGKmV
84imhyWnDDfp2KX9nCbDTipxkaH1gbbpt0if23eIjATM2xQpK6v+RdOry+7PjEwqNzac9QyH14lS
DJQJDMBcgdKkAxpfcOG5BtILtu9ROSu9S9iCXfJ1exk9UxmKPMTSE+FGvNVSejTxp9esqG7saIBs
dwOZuB1/sWMoH8D6OE7oHIto98fglcWvcg0K4aN59DKsdPOIXvoTyWAOJ0zqt1hJ3GAualpjI1aW
ozTssqRcbTGWgDYWO6V5M4diMCJzFHmf01zKpgzLwZHBokL63f08iXYlWj3a+iaa7/6yEc0+8vk0
CTpCkLxsVAwqsbG3LUtV8RyTy7YCj1qkX6odaX3qlPMxEG2I26xIlxNQRDyOWiEKO+3x5TD747Wh
PFUwwUUz18/dl7DqFS1PwVeZSnLGmU/OJ27nIJTKxykQCXfdAHL9nBDAwKfaBke5IWVAIosXqrsz
GbzjqUhaTtZ7SirdXpQQbtJvpxU2sd82lJxfhueEkmWiWmqMmCkYXgirCtTC/Xp/k3BJdjwfmMZC
0QHFMpcJ6UpF8n/tUcRFIPP2tQ2CLCoDFBI28f/kWqdIxmhOZG812iQ2steO0Cm6NJ9V+MJcg2YG
mN2EMweF9z51N4jQ1WJulXsYJjkQNDZWVmYDGCVNb84+OEFjLceCer05lB29uuvthaGvVzw1Cp9w
5HwnBz5bla5/ZQIB7DUcmacScR/LnKaWhmR4l6HYoBWNiqyUfUHGC7L6GfZE/Q5Fklvklirc2Rgi
U2rcGMRHmjoSgGpgEi1OY5W3E20IoBTC72n8jlwew6gwmmJ1b3LMQoAtS+YTmwlTdnve6g1wsFA0
jUtnqhjhH/KygzzI4QbyN0CZqnXXp6yyXDbIbDAi0zMWC1dQSPQZbjCH5eVeab/pjX2L95pfvlXB
FObX7pTCQHhZUFKTVqY7TcVDHuO7Q9x3sEAySmiVoQqeFzgFS9s7dRb3MF7DheRcNIjvwJwQ5VIy
vKv+CX13oI5aOxhDPthyzqColbkoiTF4SbqnH3SkzCABsHvavXIi5nfoqdvJIC7HY5I0EkfXfv6L
flg0/pV0qRxx1f8HKoDllsBOdSaY7YglIsznLsqtABK+p1D6bRahNDYN2RjzJU86mmM4xeOR+ILR
r3FQtEW9kNLGGc3bzHRMe4aQsJzLFJ/WxsxJ5YIIzWEQE7lnEteK4EGJs1WJM+NciyJwUui1OftP
F9mmf1sBaoJenBE5nPeKEiK0C6XDvS/xAocNXn3oG/OE1e+1IYAkYFwjo7PiWIHQx1iJGPwgoC/K
6HyUU6nqqTHORdXAjv1hyIYCF+KNcLd8Vt8bSSpLADx31nXJnr+7LZlwe3hBqPLluUKGhjCtsAVy
jL8UhGCRJ5khaPbL2d3Ga0otv+2WIV1GVgfVnaFdwGP5lATGIvTlPMQFi6KmmkYpAYJnTn7+CqfT
gCLnp/0xoBsu0htZgR+5AEHrEiB2IFxkyqT5sdCovkXg0HtyoqSMiku9F+x3PSTiVf6S+M5AEqVe
LOxS6OakxGa4k8uZ1nxWO8ToAE25dT8P+41/sk15+Y77ouM36yKsHPyFQ9HaJI4wV/UsXyWXgb8g
v2YVkC4VFq+Ch/9ZIMpMugOJHtz8ZFOVElqUWRiEQXKnh65wjmJCfbuTDDjo0u2VyLqgs9ngWdFS
zKNEllUJ/Ips78NWXwD2mwbxGyrIUR3fW4wZnI/HkivgmJdWPkmMlY+pq6TzzzVu1M8vgJkb0S+f
curOI4aJNyUQj/3ePCZ63B9c9Su6dYIqvf45Ebo+bKiHSaYaSUQzmW2eHGFgziOjJiq4B1NIeuCN
9wrV7khV22Z/otDJOkiFGWGwymK3NHRVPncdz9lL0MJXRcEQC7oghbc3Q6CAAS1cyKVOdLmqT8It
X6JqvIErWyjuJia2k55fP4ANMHlYWTnV0RK8ugn5uvDL55MmGNXhMC0WLvcTVZKWo+2bDLNAJ1a4
C+hawN7iIrDiXK0VtiQOVIqTBeYBrnB4PHOAVZLN74N26B5L9eW7OxCxpuMCQK2phss1k2mkVPoG
xHGuOi+EuQmcu4WJswVCO+NoUbZsQ3nFggtrQxKl4H3wL4FQXPW4CHWwYFp6aTN5rAHg95v7B5ub
JgT/ZxDWlxhJVyN9RWkxsirZww6PjN0yYxgZsWOd9oUT4IeYIc89MTNR/3hhzL5HN1nuOyswbCL4
11dhpSJtXa55nN7VrOxOipdiLzhd8fbf5JUweL6mdK7pVr4xw4RGTMOwavXmta3Ln9L+6alvvtoH
hghVG/IaILsrmE5QP9csNm8rsOL/7gTU2iEAwUTX4H+dGq9M2nlIcg7ieyJzLz7FNaE0m75JmwcE
HoBmrGDGuKhD8kk2HWgE4hLIIVYOHeZqBpRGOB7o4W6iX21qi9oxYbCzTs3nGPifIE2Cj8svCCsI
Zv69TcFlKpk0qonwIpwbspf+nivroU071v+OwAUc8vuWs1VVPAPcNvOgTtO96O6FgqWA0MW+e70X
sE7RMPma2ChEsMP7/UYblHpFJO5pMN1zeTUpNC9sJBMaxhtWCsI0goHTT1ZzHSLk30BVR4bE1QlB
eVP2H67Gmvrs+BkKlMHUVSmxE1nOO9gFt9sNoGgG/jfX5YdpO6dSaGUt6VIOnx1ndhm1jnTYnaB5
w3ExC8YndFvsqi1FURr0BPf3M2lo0rrQG9euGaMgsK5z2L0ukTXjPGWyK4ga83UUEssWjxy4W9hn
Z9nabSUZiMyGbACZity/trp5yPpV2clZtKSHI97CCfMqjDdLbv1/CfN2NRvEYaeMC61y3/PB7D5a
PCDg0772mip/dGAlGr3GtXIr4L8xv+r0DjECpKfECNDHTsyrG7s+y50XsUhg0eLIrYF/m4Chula4
fKn2026+n2gyeZZCqUgxiEzz/IzbpM36kThcaGJRWJZMfXk43MoEaOkMECJTzAHdlvhNsNsFNDvg
r09bqkAXOkF4hiwn2CrlNP56DjzYbY1/sVjZcMDC0olvLswl5jUM+lr19xBoS4ZZd6R6ehoIqNqy
J6wr13cq35joeGQ4w23565PSXw9y7Py5o6rcWzRwlL5apIVAsqzG3YPrIOAaUx7PR50JHJxnGirD
xKrcBDwZ6dUSw8P6DR/PgOwXQHgm5/OjrS88T53Ir1it68uGmicuxQYgPlOq8QjePlD+9zGiBA39
2SRrYHi7uLBJ7nIW/LoJgN9gymTtCWRoBvurbmGWpkhvtyfowxx0jf6tfdC4urK7XIr63bb/dtMt
AOqtAB/iZ4ZN4fp3grqDkyhWvx56c74FUc8DDoSczS1N9mTJtvHdacnhGF+FrCWsrzqr01gyzxcS
jV3DyDYlWRO45AKPTxvrP6LVMj6Iggyg5NVVOa+8bi9HttTTrW1saM1bV7AFJ3seao1ObInvSg9s
e0LdmNZiR/vpS5DAwY8SyjSAkUBBolE3qHNcdRYX2ttA7PvDwTEdpRb7eHwCJBsJDU5ygpnx8+IM
mltA497eqiFl8fMvuAjxBnXKAhgjwSpSp6Q9GwA6ZQU/pXLw1fiEh/BgmuJqAHHwKGRCi1Zs7x4K
5CpxV8NPusZhFUMHHetbzTfYyB6Gjtgf2H32+IhLt+QHO2lk1Fof2jrPVYChnAOPTE3Kc4CtI5Yc
zbr1yMg9JD810SIZdJw+ilfu+lRrXgRwy0rZFusDmElAO/n4JdgW/y/EA033kC8OyRdowYMhsLea
Mgj1YLVZdVWjZuX+op50PooKAAlfk96tP1yMcefJZZDbwtTkiJbELdetHvIM12IHksCZStZP1HQb
e+aCnMED11AF77BSzmcbqowZjrmojHnCUd05pDCSmqKiqYfmsJ0HSW9HKnEFh7ZvSx+f3aCvHa/D
xKEWrtk/Jld9dcfgAMRLq6GfP6go6QycW2YWRyZQzWJaOmmkIg+vXJ3FGbsl/7J2DCotkDNyFEZ6
+Sv9zcvfweewUR5j1iiT9A9XhkNlmM6m5LFikZnjui5KdOQiPcNIlvJIPDon77Lay+t35qOAsSpN
sxDV1e6x9e8LHgyNDMe6X7D3gZO8oOgQfxtZuINyO5WMrFInycjGzSZXKMZJ8tGHBPC1jAw8TMIo
0HIOiUEwPSyQexSXZ/WguSSSAWpfSzdEgvuvh8GIjcNUUvPFLgs07BqcnFsrQFPTvq4pkT+OIEzD
KQYvWRJoFK7Qe3ddFi5ikBUgtr4EF6lmORkBcNjC3nnb5dtYtxJQDF1FiyI2p/OgtaB33RIywV2J
FVwr4NNNBigKJ0PbqFkk5UoTS1BxncHg/ezK61oLscIUDFDp9ZvMfz7gy6kG+eZbLMzCvRB6STY4
KRkk0/GoEbczvdlOLcCFS8t4Q5zAeLfx6MkcJDKn539FQUVke5JWr9t3eRNKUCZW4ZYioO4n0wuc
o+ScZQVtS6hlFvlisAG/Y+t76j96t9EUcsMaLFGn9da8NchxE5ASBFOF2fZ1Fuz9AQIdMDIbPYlP
FO4RHboMmcEQ8ORz2sFShnfNurWB5aq23d9dZaXBua65aAfan2oJGpd+mY4Z/p/SVFcp8fYq7ZgT
BU7cr6ZyVh0V2rgv4ylbWLn9oVmS3wU9TBR6AfGGbGB3iTZFMdLeu5XeMynvdoHs62q2kqrFbdA5
uIrixPQe3q01mkDp995fTEf0kf0DOBmiCpmxkp6L7rwzEoUc4mcmoUINJqU74SGJIjoakkzdeCVC
6oZAs0CwT/tfemyRlcZTj8Yjenc6gGG383ccdxrI1bULshcLFmWCrgZQCE56MARvfTYNH5DuLNJY
3JBpjNmZzY5+FJ8j7q7zT9Lu1hNN0lX/aw/Dpx284BsE6/LS22pHUXYi0KlMaRAAddHfLJBenekW
QT8MQrRWquYGLCbnJR4ScpW5zn+Mu5f/aLgrmOEsDcBk+VHd8VYA74Esbt8SObCcV2F7wipoGb/W
zDHBuVjjjF5/S+xUUmnn683aH7zFf7sfGr0jT6n39NIdy6q/c7zmNKelaNrcfEKedtZm9f0gj8P9
/WplBX6/g6TARy7KjO0uBJWTvOvXcJZoVKzq6a/wUpv4WebrdeiUuTGeVLJLgaceMproa3T+YWRJ
cKchq9Iz+1npNlXJ16PY7xZcy+Zr/Q33Cr4OTc1xEBJiIgvEBs7vSUGXOJDftUaomJxPPv4ffCnn
laBpMgN3J6G5wBHLeHxZaU4cx/Y8K3CrpAigrz4vzUvkKUQLI8hzpn0AwP6/KPBV58LTcTbsvEya
N+M7IYDc2VmbuGFHEb4lrtVOnPfq3NXr9FK9Aw68qRDqoWnWhHGLYxUB0maBvbFobb0uqS/XAAVH
VBjo4eJS/jf30IXzGoNk+4Y5aOxlgWWK7Ie0jwEoizNjcZcFTK/UFc7ECIZAGsBGene1GYW7/BcL
Qb2Ecj016e6T4GjcmJmAk+S0doTlhPO9VH16CRx3PloyQivf14z7NBxs+Hu88o3vYLxCtPljPshT
7x7Xya3rH5RbpIAQSTuhYRFoBZ16XHYvh3kovAo1RSlnpkFLbTGf1WbcxYuuYRComa0B++IpKtqk
qxeow8gWEpNW2/bCVTwZt5y4Ewmk44Y+MmratL//C8fxw5+IfLQOVYVvl1Sx0qKfa2yQfBN707JC
Im56YOanTo2cf1nv0n1q5H+900zuIaHCX+MojM2Qdje4rX4aD8IfJ9cUb6j+zs+P5C8cMSx0hZGs
+rwLaSUk61s6CwADF7zqSwcgIwuCghSuQA/sBbrEvq7/PruhkysF2vC1vdycyLdOF9egekLuSAoQ
p5mYJzNhVsHhOr8+Eup/gF6Wzlte7TZEmrs4qGAAHcX9Uzk4m9/OJnS+LIlV+oEIbz02Ib+FLYKY
XRdiZHtun4vxzCaUOKZxVeCG6Wi5F4FbuoI8dkiepEMtYg6oZXPAhSS5uuDOVgDAVo+Kr9zLXDbI
drGb4NHTNmlceJMKZWbn++bZrDPJQWiq8wd+qHnh57uTtV4JbLQA9Anx4uyGKT62bYXGsfP4rvsD
5gZruoohZcvETcS8yqW4p1afyl2F7a0JS2UqSlNmWc1sn5rKjqxmXogmhiTC4eueHLrtxFirncVA
8bm7+zcXR2YAx6dN8oUc7thmLAy5R773fm28CVzSzLnsmwZePN0N/3LLJFvqmbwiD9OV3rIhqusl
h5m2gLiYUlIBv7Bo1RYJohhGdGRuVtaa07Yt0/ZzOVtE0QsTObkbxeixVCryv4NwPk9kXQwceZOf
GWwK0LvTWKf/9p81x88/q03Nah6YXVHkFygKG2SpVY0ANyD7HpNvTcD17YEg+lC0Rd+cviD56EEb
1FuLLCy3W2vRnFucg3MrsuPLucOVNd2gImmqwLNMDdqRT/tLT0ReNSzFLIszLeW28q2/tugHX51I
xjmsoSTVKhE5jPienyKFprr49ENrYKcAmR9OxNNEQdZRgbyP7qR4nUGxymh+cEcvmNX+baschWjc
vC5OrrE55VBuJxaP6neVF073awsKZemJZTRSOS+LIIy4dNjcOWUiMY/JHfN4LA+tLZKKuO5VCgQi
JjD/9Xub+2Jy2fEPPQ8LRwPWV+hq9MNHlFNjHsEMWgY4n45pOVhDqEig6JCDyYA49HzFC0ztU/Il
UvxZzYXR2EkvozEVqmBDRb8Mly8yWzIrJFwTt2e6Y1d8PgLz9m1nKmk6R1a2U/f7cipeEoLc+fIP
t5IfgjxJ2lV7aPQcKbpj+AO4BxOefXJGSWeIUHWu/ySzLtXNBDuBkGftlXD7R5yv1k5JtskO8Yy+
e4EPrEmRLpeA2N3uxqoScWQEWNjRI49sqKvDCY5jSaYcaoWbbb3RAuS3UUBDTT93zJlVMUBlJJ+X
msZeLpO4uPtKduYuofFAecYGC8ohDz96x3FodOenW4PxcInCBl7RcCYazlLUIgIoygc3JhaeQYw/
5L0D5u39dh+gAiYFCdMxsCsT9Dsl3W5ojWh28r9kgt3mACEVxEQsUOF/CHD4Cv4JHqfC/asGC/4L
IIsGtMZw675HyK13+0zkPnli9JNrc+MATCK5296Gx7Z/CghpWqwKv71NqjBq6GdIcuWOLuLIsG5V
GVsNOfqi6fFRK3GFSSCp3yN4KO/qftkTB+eJt1mdv9E34m3jFWdL4xfK0yEimTkWvWl0H6Iz6k4i
TKAS3azNQjCpM7/wC7QTuULtln8lbgEpJVPtw/WrPesGjC0/913GuuaUA1fl+eAeaTg0ZurV7ZD3
HH0T9vAfxhnQnOms2An/MbnpxWofa1/oVE09IYu8FH6kfIZqjkPr8WxcwNYy7yW6pe+cQm3ch3rW
SK7VL4KAvPJ82sIz4mIUaaLl0nEOQCsXgRx4KQyu680LkbYdm8zUZayJ5i/EPCzsRcCsQrNP055v
/suy3atEIzsrgqIH9q5/sLe6z0Ww8D9+LAN2vLqBcAYp0oEaq9Z+JEtZs5P56Aj25cX9Nt7CnDx9
C/rNqLCIrnbM6JxPnYeiaydfo8Y8lRYfn+jYRU+XpO3CoQuAiq3uN/shAkwkDvVvhW+4mcgw1hY/
1CmTcCjVGJ4RcsVdkj1TxSmOtl0ut0FEBq5hyn3yPHIQtGc2J7Tvr8g19NVYnMwYB1xFqRnisaqy
MUXEVcJER9y/IR8x8v+2gVzwf0AloTg9CsQpfDcMrDmRAs6tVJ3InHQxO7kOyjViants2gN+76Ex
rzkOKWjr99gwEtio9NDWm4VW359TmeyCEtxuM5XgzteiuDd4ftYxwLoQ6GEyhUN7KYvSSeykyYHI
ngmIef+8PwSr9GDU/JKjOViWZJJVgjZaXcIWjTT2v1FqirVI9qz/Q37XUSgGbSpaVdZvrHOZSmDS
QNNSKBea9VLoKJ/vcFjyI1K8cDNJluk5C3yifyD3YQ97654Rzcth+99adOxf8Omg/Dryy9qRh13k
2Bv/xYxXsevuO42VR+WcpUElB1xTzxZbBO5si5sPxNUdcbfYPMa1r573JOO9hzDqeAueusQD8la0
hkN6BbS/nyBnMT4YDUtrtz1aeR910pcR+KKPhQa75rblC+PPvnzuEChkJ1D441e4Qxv09gSWR4EL
5UxBld/3NQQivtE8B8kLOLDdPLv0e+PDBw5MPxdihy1RYgoMXJqgeJYjxMwu9n99iKlrdKXMHrLv
zog6/vxlleidfIBpX2iiHJubwsxrBscISah9rA6B3UKeMJ1W+zKiDf1aAINrgHirXLtmRrSds4rt
b8J6THe/11uerbql1+w4nW9wWmDcMO4PY2/swGmji4Q6DIKMDo3+sfixFYciZaj1tQ1DM+dwjFi8
7Cnp90QxwiD+ffEPw1ciPSN+XroLdWvXwkQBvmtpQnC0IvecEL4DbPkpsRifyaZfXp7DW29sFYnY
tPbfcg06a3xCvQY6WuXsDqzAfhw4v6gR/QATpYAOH1fyZWJmVBTn+y412TGRcTLUVoWjfasmTbK4
f6+19+o2vaI9b1xyGlAoS8yJ8GEZ5JREfpa1JvZNa282D3HAjrXmGnyxJUcl+o5UC38XvK10N0lk
SeBhuQsAefOhuqWRjPJ/xIQ+aU3hDQKgRo6JAYwZJCDrOvJ7cdVFmgkFup+iw4Cn+2pwsVLGfroR
dvMWB0xGuAD1AgfMyLMVwnMbvKsPccI5SmcDit4QPbxR2hDMSmRqcp2rxBtrsSHXsBXM4qM64dkZ
n9yQ1XtD5PbLSJFgSIXiWhXNg02tAyKFQkbOncxr2AprixXvM3IAee0p8+cRtMmjxrwTuYF9sHgd
0Go5KeXIL+mL9z3W0P5MMbfq+3zyEtzqUaEluu1ut+HLrLC3UiFmLyr0WE5OUHYFReAxIxXZOVgv
7u7wwjEPH6bEtbCvKhOeopmYdCTEDspQJqo/fJRngjTfr/8gF+OmtSUGpu1kM1Fj3DS/AoLDY0ZJ
060XhftAFg+jU5f66PmiHpaPDf8Kn0HwVDwTFs5l+rF7OLYpu57i0Vzpn0c8TklgAX2C942AxWUN
gqqATHTC4XAlMhbs6s1OeUMgTaxJKtE43NiQAQxyk+3Yrz53X+Vo1cHtq9TYKdWJufh1Y3jlQ9MM
2ISpfdYUncF9ehQVujKsCECi10UN8tosUZr2zzREvDw7GxiBUtfx10diThi++Rx4s8ewFnTpKxs2
3O+ioKgQ3Pi7SULiwoQM2TPj1rV04aHGsE2DVYoVIwfSOPDPd6PZkCXaA8mfNWqYI5+AIFZ7R2uw
SFiIUFJ3UprmtQrJQBNQp0eaDP1FyG/uDZ5fTsOSKE0WB/WhgaxxCyrFyT1a5ckC2kyXcjVK/JY2
1KZ0JxXMGDvG4gjhyOBofTg/JqoQDk+NYeAw5W3/MWteFTSM13gdhoRL1ri7A1GpmTL33s4au2HT
PKX+l1bP1RYQDdNF5lx8MyfSihbrZkAcCck54QM/mtY3IPIQwB3oRfp1SMxBkoRAnetNIVG0XvUh
m1J6eALx2JFli3pHSw2DI/C79NKNaguRee9jN3TUo0sU50MEAkJzcGBlj5Th1pJyyfPhgbMpnHCH
rE00lM1eWLUccvYuiwA37oGPyDr8pVEBcs99FnMX9aZgIfI5nOdPSFaQEvtuDWc2Q8YRmdqt4V6H
FzIfntMqBY/fSJFZxeuHjwMGLQKFF1vEnKN4NmZ25k7Tjq0cmolIC3X0K51zORNz6xj7Md9Fe6Qq
8Eg5J19PN3Oa1nnAsEmRHKuA9fUO2DzR6KyWp1+DFlIhhI57vaoHdy50lb6/PFSAtrLZL/PiW7k8
rs7H1lGeMXoqx/rKUx7POSQshgbJj0iCWcmV8EpMatbE1Z5kIeBQ8xMi0zdDmOk44tIIjnpEgv6o
n4S0qNesm4tfzkaRySpbuvaIPugmH8RJ4YX9r2lkuc4ZvM3EU74ahULD3OYOhfUsUjOi18v/4U1n
xhfx/AP2fJR4paskfgkRqiOJ8f0+R5biBJ5QN+BInEQDoGZFxh/t4uykhEz2wqyz71ZgJ24ewLZs
ToW8EAZW///1YywBDFYt7oPWgA6hCxOFuWHm+lTQ/X9xLgIurUDnObO19agCemB+dqY6urxnQ2wO
hawf4SgXnzAkv1eMsmDv9rdOhZ6tyAeUgWqpq/q9ALh+JQobmxGoNRKQXT/CMdULUoXS6MnUJ2w4
+Np2au5HfLxIz9zDpEJt30F0F8xAAFKz/gD2il3I1ZkNRY1iy0zxeG7tLqqFe4ZU1hmTM4kGFiGX
4W/agBmLiQhI8PHLDoIOOIyl+SuK/+qw3K0I94QmlibO2fI3k3+cniQUxjjXCOFewU4wvkjDrh4B
Nh1JVf/cGKqDbDC6K2d47erOv55ejKK9gp1MvYnn+vt4EyzZREpA75eQ+oAB6ZD4/ZRAftT2relP
lskMVB8YLhuy8W0i5M7zaw1TJgLo6jzJIuwBnkFPqLqe+vfmgq8sKfioxQ6L0IyKC2eS6/fj86D2
2nxEa1Y7wPyU3n86aNtQCCw8pKTnGB4b7mioNoH6O3+t36yyKLkTFYue6BBKdWIObrsVJuxnUR6t
RtIjQYYRmaDNKFLBqeMPI9EXK5rJZontVvp1Is9qk7ZM1fMyLGdGH6RgRoOmK15WU5uvc+uixS6e
z/uM2qB/adsopil/WB8JFzsqNqdn9WAU2Pw8wpJbcOAkKpeyeK+w83nqpiWRlyfTjNTEb7P3uTxJ
CotK2mGKEgJl3pjZDhBeG3+l66G0lGPI0wYaun3DEph1xma/36urcYr2hdaAY7XPVerFmnSVErFl
kzjUOGjaD3O0Fa0HEeRZCAad/txa2m2n9iU8DodC/SJUuM4byYpDPQpttbCTGGw/JsQSk6ksOaSp
09d+jaekbLIs7WI/d4puoYnxeN3Bb0Arv3CcIs+BZHPqnMuaVDvrJyUe+d0yHuqzxc+kxcIwlvES
cyXas9nFBiptRH7tQ6C/sBZP65S3QYJ6zxcncWyUKGLzFAKRTKYdzla8gAsylhELrR9LFvzGtRzh
b3XNp0dUVr82yUoxlEVBTXxDEVRZZXlfeuAHBgXEngLxTKd2sUrRMOFWTWBmYIjTWoEAPFAx+sbD
IKgPBvFNIuMFCuBK6RKbzfMFnSlt3v00kDlzWWN6bdWEQhOxa/0oFY/1Vzs/f4GnZz4vrt5Xq/72
OKiPQu4eXzaVgDZ1aVu8gY1azquTmjqmdu3iZGRdAnh2iaEg0pvRvcMA72IOoWn6PCBUgYAyTisb
UY7/5DaOZ4b6XzKVyjfwzL4VE1XsqZBJZoOafX5ewvUcyFre11pEYKEeALnrh2C+7g2DVvrOu9R6
LlBx3dnZpxqPsRIgd4GA3GwLjMJwKxz2qglwCd6QXe2PzWCozmGlM1TVfsQ53bZ2oG277yPT/CnM
1yIQqx1YG0++jV/mek4seYkohi29FmVvY4xm283SlS/6YMR4W6FyIYNbhFGXT0wH7O+UQI8SIqeD
Tlp5aR15dZ7xN3ooOF+NzNq74lYvOAs36gLMVN9Ulb13MZaeQp3Te/5ycOrKhBfoqMO51oU2cuE/
sg/9EkFTxzkTwDv+Xa3rmOiM1xPRjo0xlZNnyx4YLGLIPvnBvG567U8qouRpeIurcghomcSrINI5
ZLWkbeJDqddm7sL1qa/ZoIPoMHoAwbwsj/2y8U4J5Quxx6uLkhdam5pSnMsFLy4g1r+gE6bAlx2V
Zt8zWPSB4uWLuW8a4Um7i8fNXtDpt39aUDJDRygkf3HqZY+4sum7DGnA1GgRIz0cp8uklaTiMVgU
qqfptTEWZjvKAG+mSAO7oQH6JLcNq0pqNbJxmeosVZiSwak/SuaeD42XS3VwWlOcTLkCUJPDECda
Xs8hlycXtwLf0hQ5h6zksefNzMJqkAc5aoY2+T4lHUh2hC7qwFgZAXTjFp1uoG2MOGBE55aFqasa
aznqvJQa6iy+cabc5mkEv/dKo1jz9GSMsyUdczvhhpsM8bwCMb6o3mhdPmngkeZfd+ir+ZD07qeI
5NCRkb8NluIkYXzIqkiON24NHdt4V0XfzRw/UCQ0QcyGctaq/bf715mOxSHNGUzY71qzEI2maFG3
HIPhF/4WEwiAw2J0dxqXWlMBL/fDJr7pGVs/iPP2aFEwfQLEkvSGkAO1MZd8vZmIC/cf5Sr3aB2M
A4m0SlFdZD2SIVvECu39u1JVAgv/IU/FGv9lqdUBtSEvWQhD1GLi5inU1onjjxrtVfgreWdVq0TR
5d5DasRDX0n7i/8yZfel41jEpEVf5pV3dGcvaqEs5di4c6OjQnSEBFUaPzzRlWltYhagJ5yIo0Zd
mhDg+cGZ2Aq3QFnI7wPNaj1Ai9yCCYbvdCjo05Iyo60+Q+aYwwsQpGk6D1f1uXtlXONM2nXRgGvo
aYGXMyG4BeyKG5HCL7OWHmCFwZfg1uKpKKsVNEcsxDTmxomvcb3UHgzj7eJbB6vHckJrNLqwJot3
hWU3Phs2D39aUPOWoazai3aTHVa8lGStnRU8vpe2+ixVR8f7F5hqdiHT8b7mM+8gfejdzh8vGztY
y7relUbTwApgoxe1qMdxF/TCgV7PNsqCHSdDXP5Wq6NGb9VQEjSsam/PDcDhilSDTt6FQUIM7ehB
IjKyZQ2k4mTLftJpp6VBC9uiWdg1CrOGVKW1WyBCFWBWc0QDZPRvIULOl7bHFUXlHeU8QM/w+TJ/
orj0TOH9GWlBKYOeeifgWRxy8MuTGwtxBH03zoYuvvqRgTiGczMlxUc+TohPHKFzyzMeKGCIK3Ao
JcMs9UcGLUM2B2hcM+6hWY+SfQfp/sKwpkCkpfqic/b+T3ofwGRB4P9m25UFVdeen7agehn4KpNE
1D3GF/F+mTB3AAvtNjfclfRa+HtPQxanGhZ/nJwzX1mSot1qJfh9NgkmoD2AakaW2lJqHEw5GQjC
5gQaxRj6ZhjUWDTsyIEmkgOZUatxhHU4Mq0qVWDhcLtQLUhI9mJq8JglaM2EtXq0hDuT3yy6/eIs
SyNaQvmvLPzNaJF1MoNEucBOjSmc/Y5Kl6uQjayNKH5VDIFrHlKp6ILFroold5QC2vi1dzAAN0P2
0oVR5FvhzsClmC4ThbJ8rP61FJRGyXq4x0VvmxDRdl0bwTW/4rYnRfTex6RABtcX/vvkbeZU+mm4
3xGvvJls2imGwnH2gBBlu2eRZ5ftJbrg5XE1WRNslMM/R9JbWvIvoQI3dWMcLS+8d2SrG1k2B4Mh
fAmkdB8bdDf5PNflgg4o0QIXf2cekIZcws8Cyn531+rH5cGusbGWI/KYX6fGC7qaTeKbe9GU1iBx
sx7TkVVGjq500ATfLMWIgb0PPIw+qJF+cj2ONfx+Lvy4yVVhnLV/7JOf8uiwkFhQpHojNYuvOWdw
mpvGFuIK72b1d8poRvErz5ftXPP+S8Twoa1wRSetjTKO5DnuxYziUJN/Yn2/wp2wNmtsa1IA76CS
79t9g0hiIJhjW7BcNNeSUm3h5pJbOom2O0oWcNRZ9GGh1E2T1M/N2yAa9PrI4rJOuPEJaoRbusei
MGnJtlkMv6yhJ2hcqqTDGJgtXd9ZUqP/QONVyYOE9UJsHTwx18fVK/8GGvb0ZeLwWbAXgEibpZjn
/c0M9nHloitfeauEm6vyy+OOOF4TpmiifCyaswxoM26/D6xys+K4u8n1LAw5MoIUoDIZjs9cJ0py
4jRouCr1qf2JxFpJ03L7sYH+fqe2G6+6NbrbI5qR4UiJeX7QFLUFJnMH7nMBt/Rz9zNuoztH/+CX
186fmYq+3iJ6TR98LjXZxiYuGzr2QONGJWPEsyC9m1iChjkKGIOC3ZPsRU4fDHpuEl0CySEYpuGf
LALR8xpnPVADnq/JP3GzBhgaRIUwo3DOaH6NQSDVyDKEfxKKV3rN7D2+NQYZjJ1kCK8vIk4VSeNI
GYKWk2q51kZ1eFeRpd8rl66YUmCLkvXM3dPryklUUdNWeLgspMClMsYvIDGHTnxK73PBxNS8Atg+
YSuhPB1WGrUYfNLdFLEFiS9cYQaLuTfT6nF5TBXdkfPmJExHVQdsmngkG0Xw6fNcFWN7fj9Lx6eV
UpziAdyeJJNJa8WHTV5pL1aMBkH5SDIjq84THkj/5+TRWaGFUhsr3WWR/TYMzJ08fEZaqc8yWJr7
pUUGew/T4XPlfYSUCC/g5Lpp92OfPYn/zIZVIg7wyhfnfISYurp6sfzmB2LyG/3S5Mw3eXaq/gJn
W/aFcgz5O+BefQHbuVy+kJod36y5DX534NA7ryHDc0geijYR6xIhqEJ0aSPUfxZFFo/bzCiB0j4H
a8zfMYQZ+1ZG7QjIImIbGuvfurBJatxMzlF7GjWladSOUKlyUtFUfiJcfKWPF+hzFlofVV5wF3Xu
Xs8wAzeP3KE+exPkk9u5bK2aHM5Q43CEgak/hpFMo4cHcfwKMkRPF0bvgnOn5iyHGB6zdyvYanRi
HHmqBrUITOlfXYtjFKz9NWVt3LT6A9db5EGSbGZlrQi1eFUp3s5FRZIiXcw60mQU8zyBJrteljZg
5jWpNnMF8+J/LF47IUAtf3i9Tm8EfGIf4B9GvfWYrRiFzrepZmY+/BYrv7PGC7TWQWlHJrUDYJtO
82gqj2e6XNuKPFBdodG1RMfz+KGy+EVskjeF8nGN2rnBLp+/eKuoBwoqr34KHpBADsFNE03PTf+p
N50bnH8QlRwbWMXstFvivVytv+R79qaRYbA6v8waSdAXo0r3ucQXrRode7j3JlEz2umAhj8f/Jh9
Bu4cHH12PClhQK7VQw0wdIplLh4dCRl7Go1QUNfNFvc6S4cWzESXEQ1+POhkxvKsRjI21Umwdp4b
bfzP+TmF+31a1XkoOt8+jvEGq2y3IhVgAjxlQiQPBCJ+oADbmivT9P7unAD47+FoHBioWM19c1LZ
7CV14fK4FLKbEhaqUiz1p7MJ9iRu0YoYP7WvSZ5exbkth1+B5P99FTWB9YGm7Xr4J4nT/54AZ1mt
5U0j68e3soSYWbq7bt94seO7Vlg+hTVXMabJg3gZXOBJs4OEKmAewc4y4TRysdFD1bbLopVuE0xp
nHl4fSvQphOZ7xWE46Dy+q+WvNT3LRGLhtL3qnpNC4doVgLMqapuwNaTxtHqPZyzU2EsQlJYHNvt
KlWhKK7dZ3OW8vil4wWv0wdHuibJZR7nw/+jMBNdQJfwYHnbhoI2YgyrR34K9QjyZqPDo5Za3q4N
Iiw1y2QJjF8dSMZIJbi0L1aesmMJ6jK6HFkJbAYs03qxS5FBNJBwPooEb6UCpYgFWeyVH6BlBzF1
1L9A6k1ZJondjHDJGVif0oHq34hkVNQfCc+M01+2Erv4xJKT57FrXnYFHruIc5GTcUxRRASXKl/m
dFL4TPRMpa+4RgWFEqrmMnbJQfHskG/Xhv9HpbywSpzmbZoNq1qFsvy9dm4YgWPyNdRLpnusQKGJ
ga9NNuip4/xRkfJ8a0K60RbH9NtOVGk5lIAr6md7cGu+A+GlkGTokkNQMTCY88r8vx4cB+cx/DG/
lvO14LpnuaMJOBUyp/fvOk7PZawUnhmeh+RLUM3qdb5TIEpYExIfIbZ+gzShVj6KsVQ5XEYlDbP6
OTRUbU4CVBaL88/G8NCnvZhw1v49EDlUFRfZmg7CSBdReedwn0XXOZcSSrwYCo0DxMu8roBAMCeQ
EgiFaFwEqD+1QXzhgmYZ7jGf0DbXoRRp4ker4guDBaUHzsmHT5Myoz2InxyzZ++cgNcGt+wJo/MC
GDXTbeQYYNAb5nzJffK13PfxUJalmIDAdK6z2tk9SHsijC57SZRp8OHJtKglC6l71nS1HODDG+dY
jQpNikxaXP4vrBVydBT128XKLY1sjP9X1HAvf5E4H6FOba9FSyJiFJ2X1guW6KomZdJcJwrMrVd2
5o96Oh07x4mjFrHD2GWBWOzkzYUfe+0HIAhFS0OGK85W62hSXIUh7RfN2thCFME398G1IrcOwVTQ
fOR0N2/MgywO3U+bS+L8qLD8bS+Xo4dykahi1Znl7uzcKkwFcotbaMD5XZCFYDK2KpdI8+G3kl5k
DfFDQcUZoKBlwP44MmZ5XO3l0dqm2Wdx/qddsSfytn6dRc3NGoWsoT2WGvPjl+gkoHdV7jxS4+qZ
XUFrvJNGp/gdLnpFxcyisRpXxMhcyjnUN2xqVBBAUAxzPKughGkppB17KKwW6HpYc+2Gfek6W78C
vYOZGyOUxYFfgmp+BlTtkyHMTRjtHC4q6rqJb252qzEL7wRHBTSMDvJIcQCpq1KtU+6uOuARfKKs
z+4Q0p6K9tPalmxFiFvSTeJnVjeeY0kI8CqSDY6Qx/rGi87iPxBTiUzS9X9KStxrzjnuOdMhZ5QI
c8fOryi0iTfVCbZGRfJS237JOqVpfRGb7KXOmCiOQcSCrep8Mw5eHiSB96FVZfpZFT9AX0ExlP7L
7z5b5olOGHeMw91Ij3OEnr1cgXqiQRKkVMSGRcbn03E+Zd8BRa2yD+SnsVOnmz9o7FptoDkglJ2E
JEUuNLPjfQH8KWdjGo72mHjtxgl2y87HO/St88SpmmJm8laQ4ohG2IYXckHrwbflqTTNrkimPyD7
HFkLsTVUCjm40+u9F4+Db2bfEi5iMdzGTEFYgzt12KMRTv0ME4ESqnKhdvzV0GccTxl/doAdbmWK
ze/KhqbCfA6qiH0aC3njjpy76xDXwpGi9yRxPWvqt9UwtCFzoeKx4cft4WJPsp4Vk+L/qIdF5Pvw
vV+P7GHy1uaULBSqW6lVwbd94rSVceirGiQrOI9TzkApUP/FIS68Y1P3jiJarq1VFadQrLx2EQbj
b49x03DbYew+Gut9Qwhm/wRE9eA9c9Gg1M5KsdJ+2BnxaZak2dKX0qCPsWK3rjzAWtNgjFG7D3S1
V7/2bILuU4/OFP+p5fgs9PDfjW+MDTWb3/e3+CILFIm8cPr7fMTHc3kpS2SmFw6Zndm0UM/DQGwE
pdfeBHHchhGEnDQtrQJ7iO2yBmsJ/9vgBvFZXDLQ2H9gY61+Ea9O3VfyGo3KN11+FyLGHboKCH8b
4TwR7UBFScZmczSVl7rvzTbfXpGhZjhTU+T5DPpl2GYN9+2ajq6vkK1w7GCQvEKbSr59DKiHACxy
UaWeGG8AXkdKIhAEmmD4Sidz2OOJnSexRiz5LCkbVOxrxUuXmIsClJH3TUYHvbV+Shoy/Yb9cx0I
5j7g2gJsgaon0mXfOwMfRTCR7q6BV9Un2yZEtgASTI45o95jkhxKiJSMM2x/JwK639GZrgt2sZdv
+t8E5TXRopay1Fu4iwEY+jJnQQp2n+CQdYJ2tVjPT2ITKeYfeUKiyxftQItLCI/CMVNMuVS5cNHs
TXUyPFg0h5oG3MPnJWJeAhWclb1g4Md5Gdf7yo+nz3vBHmtSEARjZXZGjn9hrvneUsTWoqBIBKVx
AlZdvaG/m9byu5et1Pj9wiIdRr1g9TVj3ZlJJPfY2UPQvG89TZslQIZcNrOK+tcXrqEBEt5BnPRx
7+u0eonFxjN+Txiy/eCS94jp/cnn19b4wQYd9OQWRg04coiOI8eSnJkx0idB5KEvte8HEos1c9J2
aHxSC5RL0FJwFqfNhP69N2xrhW46A9DBcKrzkhvyNQuvVH0aQOHViwL7Et6iAsgAWgVlJaHQL9UR
a+nrV7SDk2SLjCnl45fcLgK0NLwSCJbaEraMsE+aGDCdGNrDccSv5SPuK4NO4uv7I8aaNqPNeURU
f3x1Agt8b5BS4GE2P2AlwFwxeArh0hwRfbCKZnj+TDPtaG+B2iFOKD9w9v3e2/WHWI1cgrzlZvcf
+6w20w/vuyN4AqYdq/Foag5+6NLDIFaxMf1dhXW2fzCjvxQTfLd1YuDjz6gYORxQKZKRcuwtqdQe
AH1lYyxvnHH8L4I2zhSbK5EPJaK8Uty743pbOsDAfr+rrJ/ZabSx1eZ/KoSvEEvpEUPLHp2OlvK3
6tTbmdzN/hkR6lR+BbUwRtN/17FhG4MR2VJVT90JyTkG2QmY5eIfjSSzvwST8Cq9YkRWjBaAQTZa
kkaogA7BXjI81Fo8jGAw4Wfih4ARJVfM08LLel91/0q0zlDjnn1hqe9RA6xuBmX5ksMuegC8DCRu
O0yaj8m/0hLLwBcyY/ZTFp3ovuNDwMPADj3acs3qqgmW+ax4cstN8Sl4OWyUGwIS1onT/PhW3c9K
gedLt6q3yIS8g+cMeEtwFEnw9pKCE9FN7YozWbAvDKMG32nrWBBIavL95o9lCrglqWIaSzXInHHk
WGc1ax8MISyxFvMlKWPg9MbXBgQXLuUU+ubVUAdMEL6qWnNlbiuy1/OPwYdiwJZ9xUdcaASM+AaA
5t1Kts7O+ZFCsiBEPE4a0AN2GxDyiBdi3a9GffCAaGeajeFS8w9o/YfzZU+OIZdZCqfBTEX8Zukb
xfMQaGcmg59YGnVvuzwsfBJNDzb86/dpfM32QYHl0cWcToHrGwXs3vvFZo6AxpfVFM2enBRup2Ts
Ct3W81VBG55MGFpYVIeltF5mYHk9QCUDFM9fgK3nJnLsWWbOpiDVkXe1MgQALkMiSRLs8j2yKMdW
kL6ER4GFVAwz8yy7PX2r35V3vYYqMWr+7oUrOlVu1Ga6Mo7Z4nyBfZPAkX/qbn+AO6i/YWv5id4/
jQIb4KauVshsgTIPtOsFC10pR8jp35kqlXkjjQcKfXPdqSiCsPp4MBxd0hQQIHkhgkj6vDRcwbMC
jzwlcD9Oh2K5zBhgi8RMcv9bzhbFh/RrvWccsS0EZDozZx63iBW6+zCmvKbDkA8U7xpCcXBCcoKU
/3Jwz8MtbPvH7nhL/WH2fjJWJTI0eD0/6pBvD7KlWluQHrWxPpWyWwSW2yge//RfPkd1PLxsDR9E
/aw/Smx6sSWdqePcKkmmVp/B+awGkbJxPhUxjsuVNtyHs5cDk/1drLTPoAPtg9K/hLTS0LJxbDtv
9NlBZNnK0cu6SR+BWkDtR3XPzDYTGeYvJ8LtnKF5eolTLJ8QMotoWxpVqAATEn2noynQUkMMqGRJ
GstdTYE5oM0z9/B3qfpCk9PsHWOeIOBCz/Mx56KQW+44Xf/a9RSL47c5O3/WpidGu1eZtMLU+QSu
nXq8Mb6dLpkTZoTpo+KazByqwvll+yVzYii+8vbkP/7UlYxRfpg8aNBcC6+F35ARe78LVoqfgO7/
l8HxvSW4ANEhGa0/X4X0gQoSwTVpWU4nsAYo+HKx4JhGTSUwxouAFkJ7X5TD0u/kifqJhEEiQsuI
9DcmZDsP+7iXpM0oL2kcoV7+wmNphUPbGlmdVvy6GoYt6pogZBFbeNNq3PjUttYM0AhV/DqhIv1Z
b+UKfuXS8hQCVAGPRkv0wfO92NTNVYzNHpo+G9E6bwIUGxhcYkk+meIdCCXRfOEIWqxZuWLjOn1f
tg3oIAQJHAXhUf0Z3M0oV2qxsOB27q4qkwQ6bi47PCA8SS4MsriJzKXII/AOSgg/rSzoNO46M14P
R2onhmCCzvxqAStHMtAVD3/Y+2PfilEQmDxCS04C5KuEej15UA1LM7lkYyv7D8FFWFN1P3kPtwD2
+zBCRmtqVDf1uJznS3rIeIrUv1H32JcyXy1JEZhOKiUP5pN+gZnsXnm4JF+2UNh3zq/KpvGv8Y6V
2scYSCqx0x1axtK8SjsHOx+gXH8Ny0NhsDsZg92QPbNRtRRog2tNJ88TqX4rIIbocYUEVbqBUUMV
NvJhUlF23YMPWpjJAKlIrdupwjDlrsTt8TcmKBH/8PJZJ6Enn5J7n5YEQSBeopbswxG26220zm11
UYED3JTT7Wz+G4zUx6pPbDsDb+AjyOluVevtm/I1S2XhwFMFKUFax9H5BVV7vYZ78hxhWZJWVRB8
j48u3sC78A8LBFU7Y/Rq5kNMDeidq6BvYqILQDcwLMbHV9VmOmu/nxDEGsC+Tgrm7LqSv6lapPk6
UFehzNNA+CYU/gdw7GVtySG3AXgPHkm28uz2wVbVB19hkR4v7a62g6Nhg4/a1VBPa1H0Vfuj68qZ
NN4UJoZc8R1qGGQhMWgnZDrp/ZxTn1+6p9S8CB56xz2MOiuoN0UW7b3BccnnwnsEg4UOYb+Y64O6
TTLs4rShuZqMRXyZz/P0+VN14xbDdExQt4sd6y/DwR9OEXONGGS3xAVTKRc8tufbDqklxqdTtQrW
Ea4LdNjh6KHbN1CmqJmiASW9bmAn6mkh4QbjjuckhvyIpCDPmyc6XaaSVQFnR4QaZXBxE1w/Seug
0oFw9rQm8Ez4Q8mg/ZAOuZo9oU2JS5VNPGAli+5J+BJK+oWKA6n19D7MXHiM1jhxt5PJa+x3s7Td
E/08AETuIegzvGSkMH5L34Gx/6wxAn/P7MoaA+JWtYL8hR+QDlo7ZyT9X/Z33KsMDWry2jWbkTmd
9fdiV3ZHF6Tdzjoile/JdSVuwzDrqf+AMEy5C1QJZqvpkSSAcOoRtMy3XOAHx5xIJI5oY/1sAg8R
IojBJ+MZe7CkS+b9/+cOsDsi9ZburCzcf7b+P1LYfN03wqWTsfiyrCCUkMs8QIt2cH7zPTlSksfy
fn5BKlCKIjiAkMA1h7qHeGdYxMcM/OGPnPuZX8U5avcAUPKYoGLPj4yFR21EOYQvoVlM0HScS9Mf
G/QJeR9FvYcdyzz/aHVFidpFnsfydFW0excEer1CCyW/2H84sb3c2tVjTKC6l/zH24WLYh8tYQFX
NGmaUavMfSWjv/gfm6+8rxZ189XCx9SkQOQqGxiygz/z0aHD0UVm09OJZDtc91Wi2KJZHJiEcD8p
Sq54mRsUVCU+5q5o6ykNa0Qcl2bRF166izzwnxjgCOwCM+4+lU3SqnJcJ16gWJgWvF0+ghFb3pdG
cSBRTmNUDPW0CnrDNenTApoFQwAqo6ybim6z+IJ1uZwFUEUkMHNgFCm3V6wqztujoKRV5y/N0OE5
/Qm5jzPI45l0rg18Bik8FM26qRg/tto1F5XlObNykYkfDfwakLUffVXJxy9lDh0mxoa1cGlwg/nA
7U5MclJ39aYpky3OuC4yqp4L9nh1q/6TSFgNlf9pqpJUon/EHQksGle8yxaEz1uNgFI97zg6vgKB
nVdp2xXOwQnS3LYDEgX5UpEC2a+e5a4wXXuCrXkvVpFy9Lt1YeJ++zkEXrE22Eek8fv4vK/a3o76
8ko9dXOxJnTcyfZ2dvbt1GUkl9ooqzwXk04R/piWKtY3zanb00+PWDKTemhNddCVpr2e2A2wVDyX
15VPjgnVYJ2IS7NJss7yZuMnwdQLJmawx7EMXZbEq4Nk445XzAyQUutHg+wMGH3w6FPWwXPdjTK6
pKiEAHnpbWQlBTM97p5n8lWwNmJAP5xIMRhjJRgW95wVJTeFZc++GwSMtrsdKV8UoDuBdnhR/69p
lq+IOD98dsY+0UZT2Vb7OLY8wcy9c/JGCsYcqVFrbuc5ZJEdBht8b8KNT2B6MkuPdu/xfS+22wgD
t5wM8e8ykIQ6d8WMeB2km+2kAB2dOAyLxLiTfswte2jRddRLYSWzJk0pt+eJp2Dz2n2ag0rt5ND+
tRPuf1XFTIuIyj24sdVFvQc/+BxidKN2pXZoNMn17mJ7hrKAiXb2ABmWGLUKFhPD8dI1GDAdyVIk
Z3JefQ2DKeMX25NUK/TpCUguW33M9GycJIa4Ffw9IpVg70yFg86SeZBT5VkAuq19WGbiaGXYqt4K
fax+uYn5xI6K+zHKd/vkBkatd2mIzbgVKsQVQ12rFJ79ELDBMSYUN/wwVVmEgy3hp4ppjKwJENPZ
iBKpHgRf1BGNGUxgVR892RGd96lmYceE3LtmReF0ZHknl2H9kDw9R8kG91f+NFLbcVyYRxLRTnd+
ylb/j9ARI72JVSFrf+VAh7U+3Xoe3O1hCkoseZdOv4fpiWAg/4uZCUpU0ANhbwn0uI+8Iaw4BMeH
faVBZHd5AJGvl4xyS//nPN9hi3sg/vnDj2lDCDTN67Acerw9PXF32Zl8oJXbb0zXwzuoXRwXe4IT
I5ycK4ZKluUYx5exHkr39Ivvpep6trLHxKnPnRXid7JvVadl2unReubdzyprWliXCeU9IHL1ZmaW
5yZwgwHe9VMVWs/uwicfLd/onbd1ja5ukyiW6des06t8t9la+6CnMG3Gg0Iist8IOhKNAcG8f425
6KbkRvHJfoO4fdSWPqCKyBKTYpN/ZZNxH3OwJyoebjrqyTHewRahQQAGeQlf7qh8/j892mo0Kvqf
RHiGYrL5Xc+9wwmme+Osm/zhZtYuWGRxUL05a5sRvz3/anRt0a3s3ANqFY+Z2o50keb+wkT+T9Hz
CTjfVKitL5XDMOsfynryCgXvnAQmdpfUjqyyaYQ6fDGM+Ru43BJPM2Mh9Ijtoh++UqnEsaWmSB8a
tmVmq7OcJVPD17UihQPSug1QEYHACQU7cNsURq2O84hawy4harnUkHoD1XureXBreMDHPj4dQ/8e
nj8qNepiUlqk/XfyEtm/ePnSfvcTqfWm7r59svhyG6Rv8KcisE4BgwsfaxzbAiwwVRN63qma0sAJ
qLjqwu8IRpSInSaMT9AU2Qsij7ScU2n+EsYQ2kvmA0fv4oOu1rbKKPjFZjZNTBNz4nwcQUVLXEze
skPhjnDpfw1mS1/9tU0SDWagkJiY1V7tEgcSuWjC+580TO3wrcD1EJMz4Xp1SvuoAslYpvAFYZWO
nMWxpJUI38JTZUGfDYLogzy+rQTOpwkFxIgA7t51eBKgvnVVjK0AstYQbNpWcLVh6T9FBBOMe/kD
sGM2Ip8c6lFHYGiUYuhcActhdok0Agh1axIPfHHB4Yz3vCpK839rCeZx2O8c2aQBrd1+o1fHgS5L
JR30IOa8SMqmZZSUIGHTneKBYeUMDPniYMe3opf58SJzHnlXl32G+59ob/cwP9ljdzE+mP2hg0us
0VMwAUHuEULei9LBls2ADglc/Y7cdLBCndMmjY2HvTzCxnyHoJgi1YmhPlM+eZrU5izVegMcGBeS
ws+ZXgk+sXWxUY0Hqe0inL0UJVfTr0erYJEbe1bm+uDqHfHxfra0MEG9/zVMY23UeBqp4yn/eDLn
YCwGqk7HgXAuyuQUMZNXP6szEfHsrPB7Oh+UVphi+j7ofXS+Si4UGDyGyJ0oPM8qo7DhZtgbzqyr
01zYOqBJf7y1s+DGelWHadghPQ0hP+i03X7y3hNTpfc2n64MNKedwU0TDoc2njkmr6VDCIY2DDLW
9Ys5UHSRWTc56GI+rs8J+uYjG7i+IPg6O+QG8YAeNmmIybiIfS9WD2lhx7Ao/8nExiRHcLdP946p
JBu4nUVCRMqok3hRKW8D21xk17uvEiRnErNtFm+xeebNtqvf5SY1Qe/iLuRmYLLP0q461yQOm7YY
M1fffgG8i1LCKzLWadN1g95BC7SsOpVCJSFwgmp15T0ahQLf2S54zuSC1O8dDjMnOP6gExFbYSZ7
Qsjizx+GSwkAkqrXEUxT4g2lxvb4j7MQ5/32uDQG7TCd9eBQCfxVJwsT9+LDsxI3/6vVNIQ12KZy
vMxvVuykoapOj4S4o3niaj0fMWP6eplm2g5igRlaJASEQZ2OKFAoLPChKs70sDCJXgTnAo88zhWU
r0TdPOgwbUhI/KiA8tVcdjzIBacOHKuMeZw+PbIO75mFxh6hbzTaIZt6N8zWvvSgWmo1p2KG9xt8
xGLMDubeKONOXDB8C5s2TSFsVxAl2Czx0ltS2HNsMJ79YMtt6jpGADIh8xDk39Ghx7j/MBGXTSMV
bReGdkh83Bt1NXSIJxJc5Vy3hWXDsfNHoyd6VzRGMPB2okc6gbyv72jP6N1uejO0a9b842I0oDpe
FR/aP8FYdqWWnIxN/G2R+LXydeRA1RcEyFLYsNEMcBOCh3WNHwJFEjsJS2HSUaLP3pZ99bfKrEei
K0AReOC1iPRcjtVKJgO8FJuG7p3hA8Lsho56+2T05psuG1SuHkqikDmT+WJX9TR4rilbyckh3cEU
jEKr/NFsryWCamrYeeeHTh9oEt1JGvvjFN7Cj/LASE4k9DxvWpvBLjoTnh1V8XwKgZdZZXAas0bC
/KJpBwHYBbJH7Dlv8Ize5CkBGvvQZ/X9ExEuuFi42rt1XrvgscJxrqOkJkk6zdbwtyMMPASj8Kw8
5mZ2Hix8Jw6ihzqfqmFmprpoRDZEu5o87pLEeGn+GtRgW7BW9rvv1X8ZH4xclMfY0Zk3m8xVYf5Z
tM5ffBzAz5WpW+qRmGSlcxKeecVhkQfuxlZ67pCHV3yitxXJb8rrj9W9RJKsYm1dmteEgguLOO2H
6UhM5Vh2TELP8+uBaRUywhOwL+AfCu8pd12BAce9bCOa+t+9BXBGFCZJYGcSIbbTyvrQkIqquo0y
br942y53i2T/33tabjoY+UYEXpVC1s/juCchmBNCAGlTWNOZ3O6+kEy2aykFGPWbXA6yW1ZBchzO
GjWiltNYL6uBnLlgARv/kBPUeWYVdB/Lxm8wrxngwCfWbCcAprMk16bTdlaGkD6EasPGtMs29CdF
k2aNDy9sYnbZQRB37htEhRFjpgaa+qZc/GrZ4ldmTMbVE7wDgHOJIqnyLC2yoIjIDrneI7SzR+53
pXejTX2Mn8koCwS3Qo8c2rTTFEdK+SV0Wn6dbDkIimCeW8CsJWVT+YCcPul2bfQir7C2t2eiPxVB
cKfleFS5sTFs26tWx2/UZENVRWVwKBQtCIzZVuE1T33qpmqffWUpjkh8unM6uazWvaTZPYuIecqi
r4F8PY921ixGAGloeirIhoGCYFOLg5hrWuFxa/6/84XuxPRbCtmOG6IbQqKy5FOVTaYEezDMqCZf
gigiLBp/yT3Uq9XTDHDQpMM+ajiFYZIhwSx7hAdGbHGOQBKduqQ0JoF2aZhKORK50sA6N6IxAxC5
6VP+wcjbgcDKhq1y0IMRtVz+5q8k/75CDbgXsrgDh/WwUNu+ZSXR8F+cD+zuNQNVWGYB4u39ED7e
4OO6SQdBYYlxgB1RVpFBK1aNz63SiRSsqvR4jEy3q+iZxOm+aISEkOj+BNF6Jy8U476gQlAN8d2r
bOob2U7nYIJCAI87zP5d/VuzApdZvgd8QEknOzq6oqHJRlIhzQkNdFU4zaMoqyrAD/yqejaAIg9h
K3sdyC6nr9ffTv+ZhGWVOXXzXzZ4s7qaNHHttIiwu0/E3lHGNWcg2tZNbFpluvO4cKILAsZCDCWO
CXhxVU/e53l/7uZ4BZAK8IQXydnRTWk7K0Wy/RKJUdrIsE3wGZpc8zA7TIl/8sle3eGemjfxpOXi
2cO/nluuGSwfVfanzW9Zz0xhvDn5Wo0TcssyFCDS7xqS3L0LTCxyWhHCTPCGhPfx/qQzKpl68A38
zt7w9aj6FkCZ1zSklnRIpzGRkqxF49ZLUS/UTyjeYRSwYw3TSGzDEJtrR6yPgCPUmNEIMg+4A/hu
UotJbbFb0f3xF0HCw5rp1JYJ8aRHW9MdLvKe48/BNTvpNqIWH80Juad3sEbdb973jlvj37Qwedlc
aoYoBV1wMbL6QWXCHMWys1UNAkR9a3Qpuv9XLwVMtgu43SEF7Hb4EOhjzeL/KRqEoewNv5zz4H3b
rjW+rN8FoWFnCr6pl6rRUcDpGY9Lc/yUS6rPoo1N+tiCeQfb9meXGAwZ5IKAVp1UkHUZMnIjGyiS
q6AIgxKZLqCu7z2Lh79XAmrtNia+cH3Yadp23TnpHdTN4/gwInrHQhrhnVpglquOWagffbCv2z92
s72dr92F0pXjJ8YwpOBhHPA+ejXAvvO2ATxKEgTGHTo1gxSCfACl8I+VQBZTmsdmrdfrZV2j5vgg
ZBkWbgRdDFO42u97PFS5kj3/UXX9EWqJ42NbDN3VbBWq4XDiRl2FNH0IQ53CTJ2Q569VNwPNwjjG
o/auYb5xj75nyAi8GlOhF/fRJBG9uA2kwXu5aGuKk7bI0Gx0ut207rDdzC6tKSdNco61JFF3uqI7
rbM7ODmlXebRiyZR6wi5IhxvS9u2qc+AOpn5DjqI4z465EO23rsJnP8mwHToLcxFXKsFtHYLFGzk
PPg4DlAEkUTaf4sb46O7sLzWeuDFSimM7ycCJJeYPHWqx9cm32cMn6ptL6oSPpLFl4Jvvk46dxJE
JEI4k2UirbLT+qz0s1mVMwzwA4HGm6n2caQzaGm8Q8JAeeoxbSk1MfebQJUizAt/YhUJbmW6gusR
bOIQ5jRb5rBoT8IoSEt0tLCD+FpyMySLMMlhE2Y9KD3isi0iE3Sutye8PNuEcLRXX7vXWnstErcF
T3Wre6JO+CoCgRxU91UufnhM4AK1lTkwVgABEInjNSMptPBSAij6DWWVLXH+A/UtQe0LbWP5MDIx
oS4JjobZL3NbGqnV1BOlTxe8lBdnB8qs6U1zwqTQrn0BBE2DEsjq7lg+HVUjNHIPkuzOC9ikUp0P
PNWUMZRdZM2gmLbPNK3BiIhUOZcbGjUWYksgbUHsuxUNfpx6EkFLRJkQGMUZzuQ7JTfWNvDvHQGb
dFTC8HBPxmx4y68LFpoMe6wYDElBrGrOhg07VlMJJ7St1VItsSBdLgk8mmvY/QyNEdIt4LLZ1Mob
NCxqM6LsoxHr0rCqe+9RcyVzwq4ChY65kZ8egIjbKfiV+bH7RrbadmTrCLLUpweUSuSRnQaTUQiX
WLtqLulsjl14gmxHmkNHB87DlRVILwnB3lpjUC2+DlTas4yKSZWxzanVBTItkfo9bHDpBTRR71M/
Qf3a6NNKuUylGOte6dkaZgsWZbQMiKQ46TP2QGG/4tK27ApLW022sBklkSBVc30ICSNE3zBXe2CL
2Ju8ZnWmHCkS6tNJ6eW96QGfIhsPUhogueXE7otPe835SxBEZybbYMVO8BBy/PxcTtCcaBCmOxtk
DZ75h6YXKKXDqJY/degNpIINzQJzghR/ugynW6LOaykW3xJlLkZLTRLNlvYm+cz9kALgHJqweWfS
XdV3hc+QlRHrLLq2aJC79WStYmPmcq2+zToV4OAl47U+sMfmQWm3L+Mf3rlZucoPqKgr6IGLbm5J
OaEHDKe+uKwx6TqCvHHip6kalLRGoAkLjMF1eH6hGoPw8mNMODacaQNWAep4yw72X1iwtyMoCciV
y7+6VGAt4+26Lb3qxfaBKXZExIj/KosUcVRlFMNxLOMdF9hZ5zaQE8JL3DWxzfpiNKI9YLWl9RHJ
s22GjZZDCa/gTjyc9KjLqgGPmwF/3G2I0aNLOO7RM3pBmuwEYn0zwhjXieSX/MwNOW19u/E0HzdP
fhQhHRWwHkOgjUeWJHRoBAKI3MUs/gjpW4tjs9fSFLuJa36A81DGaxIICs+rcfgAf6s0wUJo2ejh
W8rIokqC7vFL0sgdJ727LB4+2UWQPwsRthqPUF1S1/QcR6CI74R+Z9Y+xDmg56qxp0Q3XF7wAvZo
WltfjjGDPIHd0qeQgqx9ZVpKI369wh8gV4pCryhm2j6ebDSsTxrh8y57ZZYlDkFbrBUctvZ7007C
1ddWZoClcuuguAvs4ENvOahU4lR41zSPBhpz1yMIop1f6mroNc640B15V7V5+YiXpi7yPxoti+kY
krlCSQnQrX0X61X/kQTYXl01WTlvopCFTW/yxiLtMNQ7Oow/Ict1QVQl0IzQTvXWKor4JdkewBo6
8tGqug1S5afrKWyo+gl7y9n8fWc0MU3UfrMwpg3vwMXD3ZCThOXEXsAFp2Mp2ka5HVIjhnQ3Go3O
6o5NmHHM/L9YVCq70PXlQ0EpS7YBd8Jvk8SWs6UIJwiIqyXDxofQQ0dMxACJ4F2kun0IAG1q1byM
hnQMc//8OmJ0hd4WaDe8teOkNNs4PgJu0tzyUhd3A7Dcq42VCd32005CeKC8NZN3IJxaJboX8Y2P
09mte5+zQEHp7HjJ9JIUvIpWsQlYjNhOjT8Tz9P/8nrVpGN5AO+D9sic6rgcopuQ7c/ic1e6t3dr
faCn+4tug93auiMkACwavol4i5wlPnCL3FgKcXc3Z8yScdOH2v4fruMcCC1F46x2KZCXOIlc7xdf
mOyeEFv8jlJHJiAQPF6BAC0wPyrNM3UN7foj85jrtTJeXEaIiHRS+bM28jWL+LTFcQHvWeB/9n0H
IY6C74Ty9O0w1YpymjuMLPJRRUoh1eGWJC4Uv1Oc6pwG4X+ao1zgpZ0yiOyoJR8fKu2XiXgQbqVP
KuB74/OYEaYZ0OVKZ65HDr4bpUJ7YNE3TdzKHxZtnceF29K3vzMGoRdsiGV0gpHpLe3yNOgltyqA
rQwUqGX6lgTvg2OUzlbOQi3E/+41T8eL4NNfIsV/ioFc3kTe7wV5Zf2xfNgHo74pghXjfGw4ePVG
H4jeqKJks5N3glYvvvYY+BXCl4mHFqc0DPSgqu4PUGhTauqplkNkxHZ0nEY8b/Js2P0Y6XJJhYml
9m/0jc4tNWotkQkCxwHaCHMGPOib2djNeLV1dCCsNeGRdeGtDvfIZHK9wtr/erWChiBi+p2l6vS3
NcLQNO5sPyZS2aQx+7TU5pIt5YSAjjJck6HwY6O8m8V99W5gJm/JbE8frKKfyl2GoYkVcSzEs6fO
8TBEE51priBRcVUnfEeATUdTtYjz57Jd8835mynth7u+PkY2tXJ70KqrFPjr7UyHv4OqBGqTJjuy
1RJEnXeWzz88OOAhrA7Hq8c+spCjcXv7lEYR19zd8F+dpPYtHrqwNOXqH1xzHIk3dw0xz5P1xwOQ
fgb4A32OqlqOKrCPuAz+4KGFTPdqALQsNCRq/OHPL3HPz6s5zZ8jDc0sDqPbYuNs91D9x3EQLiJZ
VxC+1L5RlOKlh51PG9UpzfPW7PV12uKTqLSqfNIUjEJ1VbbfHu5qVwA23ysUuXe4ZEWuPGVsdMvx
BuDv+FQ6t2hzd4k+G3rPUOyCy+8KbUm8lwNa2473wH/Zhb3bzFtPGzr5ZAEZl40EHkzUkrYp0ISq
7eM7VtKMFsAzZ6BYlAbMBYGlYtYtZJ7PNEyQjiizfD/YBmAEuSJcdB79wyU/cWAT8qVZg1tcwB36
cgo91CydkqMdNzC0TwxamboOj1XwuZbtOiwTr5Fmne8Df1YVizUDEtM3l5P7Nu6j9VryLHL2I+2u
NaTuVTtka5wkBzSJZO4p2M5vg5tGu2/0JFdO9phgbltL0AhWC3QOJLUsAo4+UUc+qbCvDvfUxkko
pQ1dy+TjwwvaianSuBjNQ/fm/8De5gyyDLA47eOUAHtD9hUM6FuOp9N5HrDJ3RFpRed/goo1hM2J
sYBGRCtHTXJ+DyFPWIp683IdsuaBnW2hx5G5xNOZXmI4Q2v4a/kz7AgBjaEeCKDFcPabWzRU88ju
uOCDRCmQfPzBg9R+ih+KheuOUUUUBldv/QRCAP37z0Dm299A/dARk2gbFgKsn/zYuuznescioPGx
issJlayuzT2dkUO1hiyArDkKdEEfgjjprjbDAnTxhpZPF9aIHYsJNlFAsg//qZbaRtCGjPIVjfJk
pgu2X35mKej+SElHrVzHY3mlLYCAYf1LVpeBDswNYX5dvg303r6FhnlLKK5qz9mOrlbMes6rXTI7
lcZvZ5nfe4GfpoX1zi1NA3qpFlKyLMxyawj7fRdHN5Gmw3EDtAZdwgvzt3InG/WP9aHuy5coLfPz
dGmGRNm8mOYL1WrF+5agyULgEi0hGsJgGX1CXDHdIxEoudBbQdIDpTr9e1cKDBCxddwWvGwI9+6+
yjRkGdUakmssDM4HeUZko3N5fJba4a9gB8xLXYUOMRNs5LWQig/Qq9wt3N1r9oqmEtyyWCym6ayc
WRcwP4YNqG/VAFj/25DnuO3vNuD/Dv/vIyCwLk3muiR4rVEDqWyS0QkjfWsBCowRsiycCcz3nPEl
tifkZTh/hHPKg/l/dP6C0SiCHmbfhuMLU+lh+wDZ4TgK3Oc6tGa4bAhmcpKpXum8Se22C0gqKp65
XngemzcHLYSv/wFO0nYMI+IPOGDMy3/fzw82KqqF7CRfCOb20TXjTV3b1xe1SXTU75YRdGXhj4rj
kwkIhg9nOjLDukjPhZ0qrxBUZDRVEZPduuiigeLBxpoYzlmHc0qfkPL1/uio6C2Nqu9RdCdb+619
nY7nXIs5q8frNR2kpUsQPn8frufPQ7yfOBAkUtio98iGqSXE6hmuK3MpM4bfP4eMuLEh9zIFC+El
RDW/xBadZTwUhbWink0vhslId63ATd2qZVwHqqx3Kp+rrV7xEnsBy2/uVH/l1PqUt6nBFNiHl3QL
JdgXpXotKuXT84jrcMRuxRGg572zeaGaNO+2dEQrEAcgtjwNMXDNv9ms7bHQyTe0IbwQXRSA7o0w
7WV6ew5+pIWrEVFZn934egj3BjB0uje+dtodIBd5LHfMZKyfQxCo6bV2VXVQ4DJralhNKrAhrtqc
JRp8IgcXKR1l3rbaSjY9ho2ddybKSg0S7+oNXI65eZm0nfQ7b58W687WktMVuiC42dnZQ6hLz0qG
VrXM1wUWHV09RvXbqvFsyYRuHjb8HASPjsRtw49XCc8ihBsUzokfC30veMrvZD5+ycgC5Hh1ltF0
OZ03xES3ysMK+yeC84hhkk9aXZKQm+IjGPkuBnvZxlXV3O4FEpytZXk/v6W+M1nku0cPPro6ulaY
fnQNwdDhY3qVhrRYs7p3r+eYoCFiZNqIsZWWViNSYGIXpxWcqNpQXlsZKpGVQrGg/maca0tSrU6L
itWEFugWJ8gOBFB9B6d3gYrEGDZs/U/5tt1eMwCYKBlbnZZbEOM1hBj5vbvIFBosYN2KXJK+kftd
3P2KPWpW+3WUxKNvsYijR6WtIy777GwWZimSYjRi7JUuPhq8X10bO5FpITnNaOMH+PJS+hIER2H9
socmcQdRVEqU7pAU0UlUcZfTYZxMnqXTLWHAQOy0KDn3QIkTO4mLLR/N/4I+7I3n7iFeD8XiFw+U
rSgWuP/pd571lU8ZZVzjykGRigdM4FSH0lhM59g0Xj9KUP7yOHviQtxTLtrwJmAtolmVan1kf3Co
OY3jExiQxWjxmTp3t/JhtbthtbXyECUoVmB+ucxUFgTgqtPOhxUR8D3EbNY+fVn+l6Q7FYJ3xo4P
EsmKoCTX+StxYtaICS1XqkfrGinUTl5QLOZAfFmQLzIv/j/RK4YN3b+tO05S4U7HNl1y2LtEzdqo
rLqkpLgbBuUGiyh1UVify96AYpqglWOaeaN+39X1N12cReaV9ucWxKaCPqCAHenKqF3h/qrKLaHj
V0V2ZlTWLhBPOl8rXgkBYPHrWhEUIEPjq28Mbx4oQR8SCV27HAM92BUBa4lr30USAuJ4VXH+EEyR
CLkDVqu18I/ZQ0swKndXrIi3PlD9lG5B2GP99SpzxLN9Q3b7Xao+ZBJyvJ62aveiEvVl85A9UB6N
/mvpMJsnbfTNbi0w4WKgOB6/fCZ4XFyVkdfGe8lu2NsK0KqAX4fJ/oEeEARC26dK3+cJf4HQasYl
Mui3rKKtyg0drfdKk5iBQqdIlTotlBNV38ERcyebp0j/tzOEZzLZ+EBugXqJYPKCA+7Gv88aJDJj
vBMndBjfpfGHvgcrS1FHwWIi4wPgVWfmZxdus5KllT9LZl2A/8ahljYX9prnB9PNxmOcG1N2mcQU
7zptaEjaQ6O8nfdvboPuU3EuojgKpZFPexl6JTTRzFn8y7KeTPaprKIf37TWNg1FwsCq/o73C77U
FOdYdS2qUgJinwERNjC7fD2qwCfNHqQSCMsh5Kh+XHk1ACv+48PvauZTQU0P0SOu9PAfcuVFUyrq
2qH2kUqk8RWTUsZKysxqgR5IgNH5IXfhoEtQfPZ77VbGZYr1pgh0cYcYLHIL/tDxXapwYeM4TdFX
KNfmej+Ii1kcrWTC3qkXrQjRi098OJAOUuTGPKlUqTvFN3qLpX3KDkRHDkyo0zx+AgXuYJyvQc+B
M2BUlqWxXqLlkMC40TYa7iQR0pEB6br3wXYtnQ+/z8TBKQoDUTGigZLB/OSz8TM3xC0oCQDWE4/7
GXObi2N/HoqUgPa4pPRC2Vik8qCfDY9UDsk2UDXYLiVgYcW7wpuqyhQBS6Z4UqxATCBVRYgGNVd0
0EDiBrH+IC7eAkkPz3vNwpfosILWoGqYu5xaWShZFe3Mpkbltz4+Z/BjHSEe6yGwV3INwMnRwU2t
Km7vtkvL+ODIhFiPB4uiltpLlzoqiltTUfpGd9kMHPNgqwQOUC5/BJjsuYPWx4BNFwm4lTV2yV0n
tTefXFOcxw+RPkO2w/XQ0LwAix9Vx91GVpQ5qrpATNIodXGd4txaWtBo7O8PI/23aTnfsUN6DVV3
cv+3PvHt4XEmHRgqyfKP/VNS+oLeMeEPY+ciyIIFlQ2+DEYp+84I0rdiaxZzn+TM7CBrHc0goRRp
2v77WgXEKSz4V9n1sIPT8MROzyJ3z/eOYRrepbXDxm7Q+rFaFanFmYfyDWlU6lVvmzqc3tlMCjfi
t61NA7K5zHdcYdYgvzc6oD+3FuL7q5ersjjagwQYTWD2IGH8rmYrSPfJO5ykR428+rI97ikdC0wr
TQ55iIKBq+4CJCPvhqoGOCFL830L5TGnHh2YN8SHcTfDRczyk8XTZ/GeuK3KZBSjQ1QGzs6paMdD
C7ypfAD6fF8Y081S7YA7GdrQBDgSBwTIXqETnzljqNWIMe7jHRTxKycNHc7JwKrNPUg8BeaDSgAy
RelAe5iecYRGsMvWRqLaIMLlQx8m/yZ5jqaayaH7CHKjiGkUOZ4i9JUgvVLAvEbNnXShFnCzlnI5
xyWb57F1MC0WdxvhX0btDZybWt7LIgsHkzeKXBIAdXzFoeR0Hulw3j5VupbDWRzCczjIG8/1t2OV
z3oZQY6A8ZV908RrPApcqsebFmxbTR7zYYsF6GeMBAJQQrUB6cqFUS3BFtsI35kdQfcfenr4pdaV
h0Mty6CTIquP1HqCAGMWrjrnMCq2WeO/fGJ6nOddX1/S+IwvoUsJmxddI/2ND93CiLRiU5TZYV3T
JL/Zo4ebhGrbEWARBnx6L6zaV7PWkAmj+ZEuYEv/IteqKwF1Nk1vH01fyqkiux2va9vkUClY/nuq
1aiwMReXzNirWAIOiDh6mAJZ24UnAkfXRgfZNSeZ9zIybil6S944RgADJyeD67SnB09xPh3vM+sx
EM9ngtxqDo+sQl5yLj2cuPYKcUz98T8GXkhvJgQC1d0c+VagzOLUOP9uywoVRJ08Wy7Ur9cYyI7q
j30IU6TJOzK2JHYheEeU/MDFXattDhs8zkPp3AKpsGmhFj4qropKhG7C/Vrn1dDnPWeVBThsEhiz
9ccltv4cIf/FjND6/A47cMw5QE58IWKrxdOBleTp/IRvNp6K1s675J8ds7KvqHJ+N2K2WQ5f9zYC
VOQOOqM2oF7pnQIazIUM9KSsWuVRjMaMqy5LPODG5ZNUZz+/nIoERhi3Z4v/9YM4Tm66RMgaeOt/
k85D6mA8JlFGOvwh/acvrE9QdMgfEhHZee9PlYn5gXLCjCRmhu5aFfKb3tjaX9o1NL/R16y2PifN
sqv9/x2xNJmP64b2xwsOSZxKvih4QLTCPpohEja/UqCpULn0BUAd73RtdyBflxDRb8QAg87EazHV
oHtVJCFXhq5k1lLMAsJUh4E8YcKDKR8+fGg6LtJkFwPVUMxMsL+oOKSjcGdqfwGDvDastW3OPQU+
fg6V78DUncv+6I5yDhzgQuuytumrZYd4QF83DeRgGVjMcOYVdcBaUxJnM7PiFs2AoLyvqPzhHiUZ
EeDjUsC3rJX8vLsMdz/GYgcSVm/W6E96Zxy9wY7yyugu+7T6WQGaHw2Xma1HNYsXgtwv1kN5XnKp
20e6Fo4O899CpCwkZ+kWW2WYyoE9deg/fA++fq0YivOAQCCqirOppn4eAdhXVP4tzh5X9mBQ5xIf
/koEXPGCY2gPgH0tLVnBH25QE5Y+XwVmBlqY5Ln92SJ0icC0r1Fwxhm+ggyytnq63zzRkH/3wfbQ
yIXG0iZM3FWcx5NzDMQs4iS0Emli2WXdHgxpg5aZKFyQ/Atqp8kJogxrjNu+yidySjKSsjYkVLaK
NpblxSfO/B32qRekiuSDtg0bpVPrz7vGFMTD6f2N6safGvuqiE1Td83DnhxTJZIjZ5TYhLqZBUm/
7ylY3GsBEGAXgDN6+2m7hG/s6XSUVtiHRCeJzBY9pDJ9pifED+NLP6cseOo92lr6mwKztujip1I5
DDUjIdofs3r7eTHSVSzOC8tXge1bZpxm173xm+ReM0fIi2aVu+V9JPGb8vaRHrqcspP2YTArKvw0
1hJD0pap/UiSTW/B2XLUyD+a3SXfquiH7S7raKkCbtGezzMsbBlsHhJYx2FIv+E3qjH0s9L9uDa+
8XbvgYit/QwLZpJaz9LLlGmfE7zO16gHxuPDgcBZKawVO5HHR3FAFIlIEhx3E0wRAOWTGpAjOosX
2brZpt4yyvOJCX7MjbW/3RoHsZ2cTTdPzXEvDVr3sWYJdnkjKS+UaJUb1c9jgh15GgFAFHCydcwZ
Sj8ieUAA1+nWFI9ATL2bg2dnLe7M1WKaHyJ+MLwocXqJXH1Ucc4FeDw5JF2/qqFzS1lMW45p3WHd
EyPvKtt8GBfGIruxbUeIvdMWKeAqfqH8bHJvDloj1bpHq34hc1o6pD/7xZ8dghOWtCP+fzI9fjuq
96zxp9MFcDP0JTBb1F6xoK6sAuKd/yjait4KZ+q/h4PDv8K0TyfllE+pfd2OB1y0xt/SzpJNeBdC
wQsh1DensJToQk9gf12eoFTX7vAtRdN695+ZhswQ1L2x+5sXgKBeCA+A7OQSamOTMM90iYYFTJhN
LJzawVzwgRiiFDnQxKmfRO2/CkG7kzWElMdhoXyLmLzKPWue04BqEQYJ/cVAtSwj9+pYKphwvmTO
VabhkRGXUtZMTLecRP9CTtZS7L0FrojJ1CoFySKdZ4bzl4UrvZebKI2er6JTagCu44jbaP72sNwX
oYeVzXq0xZdspMZnzw/VtT6ByInNr5QB5T/NjTo1dwIwtGyG4n7umYUctG6zJzq0m+knA1wY0Tbu
NjNWNRzQT7/483J1zsFOjOtbIDLA+VORdn8+m7HTtZ7oALYg62B3qd1aWJCuEO5/HONj2ViRwr1U
jBGOwr6vMnyBh8dl8yjCL9gzPRVfxNcH+GJZCvwOp0dZjU+ZWyxnxlPLINLDVoFNb1xQqjy3QV2U
xubfLHbEJ1B5CAdDKEmia+gcuCeRs8t2ZHkL0zFN3z8m/Xkevr+TWmOQ2BCw24kE0/IA3uWvJpOe
iV8wpYshiwZiopKXcFYRMOWUm4IwuCozypDHl6KF17IWiMvy+C4fULSuHKiFqfBepIhC8qXCfr8W
0r4KmTVBPl3DWmhfe2Pxsuft3YgopidE2ipLtYLctj8RPGPb093ohIuFc8tydTEYPHcSVRbywNad
xF04EwtrJkNr/ZCqDVov7Hr371fSbwYjhNoxixxNrCHXFEK/QS3hKgqTtkzuuDph3GMwR/Ty3j/V
ZDfq1CpGCuCGzgeb/T8hvPm/s+eSeYWHTZk+Ry9Fx3B6aTAH7SB6m5dhNbIEZ3rzZZTE2Atpw7t+
Vhrd2z8SUe0SpFE0KfzwB+qPPWr98dUmUaVHtigNz5VXsmOGTZiszROaKZdDy+HesQp4H7E9f5kQ
+Hvgt5xX/ayps1SPJrWGGBxRlQOhTcx1npgTz5TaM+PhxfT97CXtB6oiunrRQYyVeTYcEPd2vM3I
3TZUM3lCRIjBXZRGYoOp9oAOVWB8K1x4/cA78agljYoCJ/Ta31D+pQ3QmKbRIfmSwznTTasi/Iv3
hz46aFyYSdUCyaAzMf6xtBPw65+HFLgZD6EInOEYFLllQxvauCjUo02pHBJknK6fy8NVhG8zM6hu
jR5gXkn5k8fAelKuMCrPzXnIFbseQ5xjy7u5tH/MvsrGYTHH+zjpsTkqv4ZyfNxOfboQXCcpFbky
Dy/qOB1YbMarmPsnVYB42NF4tQIRttkIUhbjlwgHektoZ/0qosQeILgSxA4kS5sqMFQbuBx4E23w
rdRYs7m4LSl82aZVFDWqXE8sze+kgk714axxf+AeCH1tVZw3c9zWudQ1YnCNGLG4tFVzkza4wz4R
bAnCRb8L3+bZGgMm6cH5MiZSn5woyif+E2qE3c/+hSjxwNB+3SI5+waxpwIACc+HenAJpX+2cKle
ORo19cC31dNSbs+28ptj3SMPzPobB70pC7aCvQk5wTbMdj4uppf4mk6anGim+aDK7hADcgWsNSJ0
xWDILp+g5k/T2amYlU5PTINaBBw8jSXWq4bbqA0qWkiyZg2h96Uq0rODOb5lcnlD87jc2KkYdRCP
kRyUXVSHFSP5B/qZmWeDm2PkfOWRGe5tp3OY0/4U/wx3VlrOAGEBvovwykDpvcftA2lN2dyvHMiX
9QdPe+M1Df4anRlgZyInhzrMJGJdEyFMw80bwv6EDN6zSqhmU9Kzz/AojrQGTMo4VCOAgiXMGg8A
KFOn6TxP6Lk+8GBldMyTRZZ+IDrCEGFnf8OAIlOLq5hSVVPmIrw/O2lE8Vl/g/IgeJ+2v0SW8j9O
A9zHD3isOvxqNX2x1+GSIPK21w04PMlpCpOZK7zSOiBYd7HPGT/+hF5oEmEGSiUrmVeJSQo4wloK
ycnGlub2IAZWBKEwRwvZT2iwrlGWviu6TdiQxORhqDnTlnQ7aw0Cth25umk+X/cfpquh4REFd+p0
01U6/EgN1KE0w4RlPWnoiG5cLHWbuUSPIoJLs8C+CjAMyAp3cNISP9Z4rjwRj1bodjJl+ZT9wYFa
874qAmSsV9I8M0TGhGSas87iWOr7DLriWj9BlcAklFrCQH79vTdPodGkt66MLlc0KnwpAttgQOZF
puycrMQodWIUZLZtlz4N3IkrQIE7GwZHxuR0lSZBHnvD7YGSgSysinvTfCAYAXvlb1GmkBrgbWHU
LwC/tpoKH2nMnA1cojAC5j/klxlxtodKgqA+UvmmGy/yrLy+2OstcUHj+e7akc2PVTELmlfOB5ue
VGxlbsur42uG9JakeMFviqyHtgQeoT02xQVPpi1KRmh8uC5Gf3zTUMB1xW/D1GJvSUg9jJzrMyNU
UTQeX6ttHri0kfThO11EsHg6JV7kMwZ3NN7WpR+jspeTZBsWz1W4cWfrkI7oHbPd6DNhaTeUeV2l
78HRQIBkPTPtsVa+JbzG0DYwjXFRuT/j3iImAy/yIVH+xKcTrLHJMiuPbBo+EcIuMhzW5v6wxUXa
f7H5PKj5P7iLasQdxaXzRj2H/GlCNKajzksDoyhnVQo8f9CWx1SLcnbF6HsKmZAxzpCizS1IvABf
36BZ2M3F7VFcCa2+IXu/0H5u2vdWKM7X1g/62ARoMfAgbPqVAX94swvd+Y1HL7i+VWzjDF7DK9K2
sivfqHYT/+xkoeh8ojv35ZXw5L2TLFQ9wLKGStG3gunDYmTnA2z2qAGK3gmANzFBuhGgIS0vlCYd
qivAdefMgMeYTwh93X4W7eP7unFS8vI+UqhY1RRNv0uXen8x0xhYRNShVFUBznsnjmUKw5NcF+IQ
22MG3EZ8/BZf6uJ0USkSJISUe6KNwRqN7W+iQ18gF3QX+k+nxX+qnIv55bHEoFQF98vbMzmMBAlV
ZljYrEn2jcuiYUyP0VTQxrGG3rPgHiRiTzhgmHBiEbsv04PutERV3wSVCtvIq6ZXq88xBO6Lhhhw
2Npkjs+xxfU4E7yorZETuQ8S+sYQQ2unED6MH3OMCe732kxnuXc9IoKJPrRsQRzxPolq3F63BTYE
0U3Yi9cHZV7LXbhBoaR+d91X7Ob1mwQXPmsK6vggNSRnqJPPFvh/UlGoZ88itVpjuzP2z8Im4oyz
pjcREqrtAFhY8YmU1YMDtZehbxiwr+i5n7Pkvz25bNETk/SqXbcoJXSDXSbRk6T57Tuj+9g6bbxn
sEMtgjxFfzGU2IQVmW5Ak/ddeg7CHQ9F5KD7DazlK/pkAuBXQp6HCZ35iS5VN1vHKSW4XHtY32iU
cPIELRBDqV6HaP4fMvpIxwqa/i/52GQtdhNyvJx60xX/8geFAe0Pq9solykGtabLVufuxgXKqas1
9YA9E7BfU0pG97nIjqaijoBjBdzljFLfV7E6ttI2n0QWCNZC/OfjIubWdQgZo/bXpu+DeoWl8Rq/
Z1ET0dbKxPiVLReisA1yWjr1xowubX0YXhee5eB04bZyPTQuY1AJE9nvwnZQKTwlTvV/8WmatGz+
OKpv57sj1TIgzXTV7rCnmr74V5LfScVnbGXabIfL6CAMG7RxLG0cDgtZATjOBMJ+q8LaOEPvPJJ+
zH4FfEm4Muk1BL6Z9ry4lgeuKmlAnnEj3uI/K1o7Qiumw87U6g6vo+RCCxbiMVUhXRxvA8LWt9PO
wG9T4+6ZfdYz+nIxy5RN4lykD2hL+m9PKSg2y7GXiXHJ9vFb0QGqhWiG7ZQZY1ebEVBwr+v65qgb
TVtL7/VzDkd3iWIL6u29/fVv//z4hs53OwXnM4eRXqIaC9ybK9UZvRssqvui+VQANyfU/cbhG2kL
AksaxHabWCojpBjw9Vz339WBBzO+Hq75pRugK9NUwjLNMEWP5HrMuQTETbEHg3goRuWS4WKzvN+7
t0wuJXDVflkr/nSfQBXmKR0G8vvTf7ttjZALvWxRzWoOTzaOSE2+BWtD9D83RzJyW2KfErVPGFAC
BTyxG9nyMVF/ya4u2U8mHshOECwXdpmO89UgpnrhBmwe8LLh6+CNn5UlI3AVbYiU9+FdSSQTP9sJ
A/XTWvAsgzetbGLAKhaAiddCjOyR545UaHgrT3FBNoR1Mo8Tac69LkxKickvJRl3TGFctx2COGRJ
mSAdTjm4TeKptdbigsCqnodRIbz/NGQXP6qAcU/HyQgkJNcLtpxmMEXPdC/9y6A00oxZ2OIkpBVY
z4kVmYkBjd2yOvjCNEKbCKtjJAjNhWCROgedpJ6uEt0kseljlY6ueSz3koC5LsLuTH9wH9HkM6O1
Xjo1K31e35eKcwwGjjKWl9INOYTwSK5EZQuj8DQQ7mnJ9CKYiojoVRKaxqigRi3Iz3l67Cw9u9zR
AxaOb73tCFhGvlsYrsZBsck/SGE6wMG6oL6oJxHsC7PrgyBj5w9xr2XrDjLPCco85rX2sNGUakIe
8ft1jCMkb9TGbykzap3ZG17aRXu61jJjqufkLrhP3bFqiRwoK1oU1evczA4Ui9GJh062+LjFlBMw
soZtex89cruAtW32vOurL97hvHeYOp/0jgLIfyYm944ac6VLCa9n0Ky6AGxUjYOtsQGM2yBnTEzm
CABqYSZ1D8xZrRNTvnTbmA95FSKAWSlH9JcQRSfxJXDVHZzB4/pdTDvHUep9a2U4nOCu9EQW0NFw
qDlI6L77AMj1inJLNYNNqGvO2JnCm6Ww223H03mV0f8BUFG2+qq2EJ+/+YyKfX648z1xATGdoSCf
77wv8jtfaN8C7ATrk3fU8tyZQXC96C0IqQk0/1uzMuupgNZD9IvANEEaIRzmEuNKnk9WQ3crJT4S
IbPyhI2swg1NtGo6ZRMTww0KEDAwE/sHKlWTad4WReKYm/yJBoIjAy+qDvddasixSBWw6GXgJGfR
Rw+keFJ7vBl68BqU+/FT5UErDNPgvPqEUer9Yk+Q4PlC/OrOp+Aj464hF1WBirxeDod33pWB3d2D
u2KL+OnkmZohhOPbngkZYrZbzvrf5A5rDu5JzQ4jnabRE3HIeaIffkk9zE9dBWKf3Q3ux7L0ITLR
Zsecnj3T/OoM5pq/kk5MI06ALHkuimmVpNImaIuLWUd0w57fqjdAA1DMTyTa32o5KdWNoI2PdTCc
VRGyIQalxUHTmB1GKYBbrBo2apfJC4lNk2tr48XN8em/2qEfm0j/3HkGtWD3kEEAL+JWCm4RYdZb
2WGc/MCJPjep/guntgoCbp0tiS5x2fZET1BcLs2/iMtAL4yL9HunQzWABi1I/fETacpB4ieEtLIy
/aC1Fg3fApgcrg9cNQ6W4CtNpUso9XS5WBzIUghr2JkUCJPDurEmmYMwf5t7rsKmNyC29f2f1z4S
UG1WU2eU4E34sT6fDte9+yw+a0HS2NT4WYjB3VVXN8qonihfPurO2i7z+N18s8NwzWIWfTeHqSX2
h4kPF2PaoVKPmtChXQ4SjBOHoikV9gP//WX59gVTPT7pc9QBfx7ZIo9qad9PB/NUBMTZ34buQ0Rk
FKAVDTbvVBVBSr7gu60S8fUluTNJlPbq6/JvamtsFj83Il1k4qJS1ZvkDNZHePEdl0r6lonzJukT
7ejlzR9QIxyiD4c9KaOZbSDWAOMPBcWeKplxpxplKzQR6TdmMa7f2psBmBhFnzffTNG0qdDDKn0l
yJ75X72/7cUesIb3fiA+YnDkuGFOyTfUpzb21iWGgK4eNGleuX1SnObYEHfjyv2E09Gy4TNNZf1D
Nc1jdgRdOI8SZvRNr6HcDWPW4UPUCEokToaMHmEN320+Gf98vxAa1fuWXK8BMVqDQ/i8hZH3/UTm
bCVNxP10ehRPX0z2viUjjXomzNRgWlVtXeScxeaGWeKIxNGCELsjLSARySfMCetc3Fl9ssiBmjK8
fxQvzkot65upxbHt0rA2Ji/tkDj+T/eHbx9erzMEDvQuIw1XVjvWcvW0Kw0OcHdTsK6iZiGisHho
S4OpqFgwD1JcAOIIUiC61+PFCXhkiqebEolIa3hwoypmj0gFn9jYvP5fKtYUKt4CepzFuWCA2K7/
XxvKSvVm+IgQds9HhYJvqsaWqJLTQP0ymPw09o9JEK3m9QuQbhdCUBmKfwsT3MHkun+8K8/gvXr3
VNsHZlWe+xnH7rkFPI/jAw2gYOckF1+6PwB2Xy3y1WvGlJnbF/xrVoRNU57IgL8dK0HbvTnRN+qB
2oyQu4R5BVAG7cQmZK9VU58dojCOx2ow7JKTCsLL6/nShxDjoDGCUNEa3F3b0IPvPYL41IA5MKw+
Q+xK9GBORzVt78Oq1+tp9LL6CGn4TrmDBWixQoRTlz2koD2sJDofHD3yySu1NK57Ia1xvXrK/Dzi
YnnrF7qSlEVhEgi5xkZd1YJfjVAEjoJZsFXkkBqxkLj6yL3OmCl12fFLGLugmZ0yisCLyIMluZ/e
KFUtRlto2NYHULgn6fx0dROVHZy7vVKQDGqJ9PxBBVZYhCXHhLJC/Y21R/JYyDTq3wXZXX7UxbUL
qapeWOUrBCYr3oXIkkbNobw+N9/nrMzAgUk3RHXfLevyAxRvBBVXOZrYHD28etUChmi5FA7M/MXT
DXHYOvgZ9EQgQ5fl6046dv+XDRygLMHL3kK47OzpXNh6srJaYwYrV2aoQVgIAnuJaoh8vCu/DLe3
s85mBu8PtgsMH2GdbVAbqT3sumR/gYyPY2RllX5HOIrK8tvlYGQuXQK/butGGFJB4SlN3VP7ZpKD
bRy/2ka9COjdKjg3RQAd8tYeZzIma4GyF/tmH6wK32tUJHy9bzhtrczgEjJr1ido8OKSKGNkYiet
zYDOBUqmpLbzCp/zTYLoZk2sKwxgaoHupaw6yGKNim2iTLitL2C95f0UXjpIt+BQItFQr3sPLS8F
PtU+H5TMH9iXkaoSs4jc0Tu7VajUEg8C+0mfR2pP49BSy4UDjLxuFHyKoLqTRicj1PFmxWmD4HZ9
r614O8aeHnH5CYWC/p131QcOjROUcWmN850TP1JO5HLw+C8iXi1rd1fOBDZiydPr4O61xUv/0pFF
4GC1oQJGgeEusuxsk3WwSRCTfJyviK2FPMu2RUKYD2DMesM/ypXh/NOwTUboFrMp9zoJ7RCjUp0x
c0GuExZFC5Triio6q1vcSH7KmOdWJrIhw2qbYLIX8KXaUqCDLUywGUJcldC6IJt/IiZtSeA6KtHU
1rZDz50+nGab8jZScVk1FpQ0Hm4SmkSRA5H6+kbkSy1OdYDbZIYuWhATDOKTIueg0V+EQhzIgPxK
z7di5QFPl0Vv4GlhRuHCSPVbeI4tGJ52mw/yBOJ+QrvjZg68EP081M+AUiaTDBSan9jCSRnPZopn
qAUkYAsl074YO+/9tDz4doDorY++hNnDTmcuyCFv3Is4rt2Yw84WhJGPFIYdGrBWiJy7ktXRj4Ju
b+m9yyd+SB3prQNSH5DHbzmZ1neCR3zzJdsKiSgr3WpRW7VnyW3EldnK/PyxmjwPr04LRkX7iEPD
ogQ1/xavzTuV8v7+PYzTN0va4Mi+Gb6Hwa+WMKKzgbnKU5A5gioEhnhaAGOR6HrX9s1xqysa+Mqk
eW5f38gp8QvcHuTWJ3YsRhJvN/6Mj84uEYyC6J3WfHhZYS2UdlraFdHrghh1FqWlvdUiNH/aObyS
k8fKc1o8juY4xIkvXlP9nwhn8ICh5ZVqZ8cnB1KFTPxKPKaANUQzxCfM2bForeAY3x5BLLRYaU39
lMFGa9MFzQF3mlnY65Y92f3pO2te+72m6K1smhgatJsuYMP6+o6l/b0srogZdubZUvhadO8FkwpR
PSlQaSZIjAJAHxbyNhT3ey00PRDWMLWuYe/hfGqtzuWuZC3XdH5MIZ9560odEpLSgoCwNMyxQz5h
HybO2KfUCfbArbdwlX+QCKd57YOEutzhTe7MdeRcXSPHI61CwHHL+kuQ623UEgNI822MRd0BPDyr
UGLLGD+KqJJv8v08i890iMXvj/M2zeqv5e373GUHsI7DifWJnvf72ijOlgNkvUKizA43+sYPyRn0
o4oqpDTogA4/zP8R4BVzI6Jrlz6SV4kkdcLCLjoTa2ltIl6rK10j54ZZsFvniHiOvNVfe55KJKCZ
gR8MT9NZPTe6K76c/fZcwsp4Lo0yZInqyKXulgVP0GjZ7Pi9NZRvB9nkU/DCPnJ18S19nHh+5EMP
Vpbd385BoStpmivSlZuEO7g/mtKbDmKV5TUIRKiffMALaW7sqXDQ41Uizy80CnYk26n36UQ2lDR/
iPHdrTr44fd3VehNW5iJ3//RpMdSBqD7IwKjrUW4HrWQ/TeeJtJv8jICV7bjAu0aUS3GIpspyZcb
BlOTZbnneeXtip32oMyarrOIBFZGnkwhkgVot/rI114GI+OvnjrWcHFuOsNkcwZF9WFW6eIG4KVa
6LRQ6M7I3zV5biGmSqnDOrV5VSIEdNxcLMjsIPzydwoyi1SbplpPGoy5YIB9E3+qFvhltmYmsz4T
OCeD0dc8eZ/P/nsgDFBm8f9AUb6VVANQuvFjkBWyC70tBkLezdMNIsyAwmdG08Q8nmj2yM3KZE1F
e9G2kb/1rsI/6TjwUd2E6Omnf95slPqClcou/quil+3c0l7MUwigW8Y9YfVoQCXGOW0Sh27sDYR9
unyf/JGVyIvpP3EUxmLZLUvqFuDyNQTyW7ayuGLonJDGlAvIQnjQeHsT6GiQMqATxOJWgc9YjWy+
eHuXteHMj8yYvf3Rs6B/4soq3HCzkgy6x2GVeTe+q/ecFSnwKx1ik2xs/o/v8VgIen/jh32mzmrW
m5j3pMLmcwtNDpsA5c5ynPPSmW/VXfGC3CzeuWvvlUsGGAsnstjtlAGDy8DjvTHQM5Jyb/fUWRZq
DFdNMA2XaTcdTaYf9inSf9Qfctwb2GJXA8LqkNu8ZBDhrd/6XQxOWWPhJXAKiItNN8B3gNXYpM6A
IZ8xN0HE6yR2xizayq+xgqEFyW0swh+IDboeo5mJoSQuhy0PJDQeRD50rvEvUoCLoAVQ/JC+9cEp
6Xtcj2J3P+T0y99R4UNULu+ptqmw+qAjmOX9+kj2IWUn51KEFSdTRW/pGk0o7q51WTZOoX37MaAs
At/+UQwydDlAts7cn2heXrCv8iPESYRc/qORyOhyQ3jhAeVIbIr+LPP/mhs3H7MDaMXSdzOH1Pzt
AvEHsQasYIK1GcKwfaP6WQcVKJa9i/8Yn1ftwo+ArrGsxhyDtGpmNhAP5EU97mQIwmWtiVx/utvB
rBSY3H+ewY9qQLOAamgtwzQRKnkHqskDxGgC3aRitZk2Y0UdhPnIZ3vY+1k+2vx1y8maK2i3l5xF
U5kHV9tsp0yon5+QDeoDl/UY7O4IvOsaYPX5XQeVnXz6FD4J1mQ4jg4BLEmtjlwZRZCwpNxuNwPY
yNuwY+EnN9BvGKImDkReJG8oWiEYRgdn9jWXwMmkJuHQ2h7kXw2Qzo7MC0B5gmtWe7swCsg5a8zQ
b3P6GaBBrWDKY7NYIeM1Bpb3jw8BY1QLbPi/cUv8s93Dp03e4z2nFxeGkgGxBNdX14rg9HiGt6oD
lic2oRyG+x5FobQ5JE9/Fu+vAUS8AP+Iu0VIhHXQ0PJofhia11tW7O+MFqvGxvppG7BJItgsyMa5
e5uTuMYWj7Zk6WrKEQ7PsKEc86d4h411z5soW7ubyzW/4cmBNpLHwOGCnIL9geXqzzGvecNhSJRG
wcsGxDJk4kjjv95hVVKrgoiPNj1QLCuyIWh2xPyuJGsGMOdfHJ0yc/SzY44UdrijVgzgeWltqjL4
SaDTDeIi0/RXVtDcLnKqNPEVyNG0UxnPmOButY6EMdaa+R351hiXnMGNAFBkky7KUWOsJPko4aok
kqpmqaMwuv3dRgsjaZXS3RyqEJ7qoAh2o3fRQIOsdBdmXXIDT7GTCBdYc9j8xiHDIA+37DXof/T5
qbaQC4udVjj48h+nfe4wK+brWUeFNEgI/Q0JLTq7powEt3UmQ34zKXnR4gy338wUvsCrgm3xP78l
g9xxVcyh1AIh/gl8aTsquK/dAPVeJbX/7cSDouV2dJOIL4WUZtAR+4fYMraSAMoVgh2kfz2v/gU8
gctH0l9L5VOLxrInp2MkMyzysgf5vAkhmSAgbHELuhCNoJ2NDph/dXsGpFwNuMKNAsWEyZImj78Y
T5UCip7f+p9/QFQOhOHuIFh5dDGZAykXDdcC0kTwKxrgXxGAqMpgcgFxEj4pE/cjrbZUX5WroQBL
B4M3Qt7RqnjCq6MBHkZgDu2Fub6JcV5soAbe8+3P+0seuGjonhEZ5HlVZu9guoIaoQC4mkPgBkjV
54sgA4YIe6AAr6FQi+QgHu1cuXAYAR5xfnjSw+2owfvWVp8x24wGLPs4e/FjWKThHfBkvfsNi9ly
QChdZ3M0xo/7fwLWD72YB2UrDAsx19kqTLcNgFFpL7uUZ6Nlk78BULzFkrhGa8wUX6b64XPWj8Hx
8pHLQ5VG4fOoFfk0TTkTdATRZUpgAWyG08ZOncJ9c8j8pdVBPY6mIRmCqbtaNacAP8Byd3bHJQH/
O7E15tPJdCH9DlZths1Z/GoNkcbhr1cBdoUjjXwzsflt242Hpo7KjuxVPoHHqlIIyqU09/XVD/Su
0fZS/lC8yoCmn+J8Ld7l17e+AOQHr/uU1TN9a1m1a5yBbE1Pra9gOVWMYiuro0fwCB0U6U90UkoB
w3BxauwwyS3KVUGx5J8XqxhFWh/WXaH1q1Vsighsq0f5jXjkZxR8NKLfVQvDAPVkTNBeKIir+Con
yRW50e6i/nuVVKj7xhUVUZWRfot+cbXPViaQJCUiFIFb4u2GyYtqaU9TxqzQyiAhLs4KhKD1gtHQ
ghTuCF9419qvdVVcb+wIQNrtYm1NkBWdyjVQ2Go/KyXDDrR40e1mMr34IhJJDUtSxXkep6J+Km2b
oDzSa/qoeVQz/lxzXt06am4nAh0SEIWnm8G8ZVkK3SiVVH2iOx7qH2OxDv3x5Jp3JQJR5mdqH3qX
8HGIupFqpX/kj+xyqZ16JiYqdkA17EH5f0UMJWUewXNDbiZQ5PDauOMxvBDfTnXtU3LYDEYMhnDG
L4YtZE1hhO1JkSmgUXhNpPhRrnS4mKhRIBnc+/kWK6MoKS/2sjny3JGHBprnWJbhaqTycxILj72k
oso+0lO7UK6Zh5cPihkA0iohi6DWWssdbP9qQJdjDdGhN0AaORkK+rckX/dWtYTY0TeLyCHcRPUE
LGjO7CzrfN7PnIpNIvUYFqEIZA43PDzOh7C/ArhAGyc08Z/yRWvVTfIYxN3dhiIojiWJkXlE+Rr2
ZkgRZeMcXE1xVhsUwzzjYRfg64K5gOY46KsuESvp614BCHKlmjH0EnJSPga9/v6yezL2MzMHiTwk
4EJnvnPYCVC6CPGa7XCNcqlTtGCRgShJooLnr48Dmex135lbo0qc6HfCEUZDgU8H++ffJeSelOKJ
VrFQZsTTua1J4zMHbfdHIi/FjVkJQngnO0yHeZGEPk6BVeRHJSLL71SwC/R3wurkcfL2QE82REAu
phoDtDjL6guGntKYwKK3PPnfZhS1TU/JWV0utLiO6wKPyTcylJCyY1Nz0n00BdeqxfEQaXX+vgkh
38oW0PZ/icQvplgX53AVnOb5sMGW3Et+jTm+4kS1Go9ssjTq5hpCYm5ei9CLStvB9F7qeKBWrFI+
ymSi4hNE+TFOFEjiuYWsOUH2f/Y82rNo+Bh1abCcGKwWrNJO4LojGjTQ2iEdZH+o7SkRKxHxaFZe
qk61qf86Xz2t05UeVlIxFLSgwu59P+5t46znelGAZkBeIjZdSNJFfxGg02tfyi1szsb/XpOZboY1
k7xfaU9KBuApuLk9jc4eEKL8b7VqvaiAc8II35Dtqz7/IBzhfgXsIkBcbGqZcVUs0rB76FDRtu+5
qnC5fuc1T7Zpp2Fv7/F/HXPlK09bfw5WFgbUoQZBuLeGCj6+GHIiucCYyJiE5MfKipnrE4hkSbtu
LbKlun46RyLrJLWnOQ4fzXJre3bNxWUcLtrU9Ly2bnsek1z/IYlLjLDdpsyAvfLWcNM55Y81P8PJ
nwPdRx1tiNeQX86F6JdgMtO/3P9XkaJkefj1Cx4WLnNuM3W3MG/4OAthN/xgCh1oL8kpJHB4OWND
/kEcmQrNsbhCVPal+xDSvxF7W9msZcnVmY/IwfLUz+HPYJuQh0QJ7ih3riamHewWfQyjgRzpL/kw
ig5vLIIBM472kfn3CSxBbfy4Tbt3e+0l3HS50GQtem/bukM0sMw1/+ZtfxFDWlY1A8gwm9scrMYU
ezxdbAALZJO3E+7pW68yXUoQxbsjUQO+l+jf8ToJu5bpBHBM2AVU0ypDQLjW8cJwgxUEleeG1ZBa
ciBYcKLuTATaYvjqz4uetpy9hpuaLPxnX9qI/MFMNDGVW6K5Wkugq2KUFvbywwFm2bBd7TUfKheb
bENjYVwNaJcdPDgiCgfJQag6t7IzzDd8QzZ3wzcxqZ11Wxa1I1s0Azhl3J3qelrH0u/8biQLvhrF
LIfUYUKREV03UMTrpfv8cdMflGzSUmKrF6TDQwpZsvzhpXFMU1wXQpywTQRLMpFog6qG6xKlRILf
U0EZoHbDu+1fQiqNmUX42uuBUSdf418OnKaP+JKC2qW5r5L0vOfgydSAq9QNJpFaBvbInT4rk100
ARN2wu8BsOFYhC5HJlm4HbF8jwhZbdeQRwh6aAvU6iqSl/TXWYPTF4ufvFzDBi/W3JnYx/mTsAl3
sHSVt92xLwHs9euBWk42edVx+o/tD0uiBIlKZHPGMuKon4xH0kzxroNrNs4mb98goQ5ffm9ickP4
XL3RtM2QjCkcrv1d1ipf4oGO3eohbzwK2/H0L8ZztiHj4+r3BwOCc9LuwiXsFsU/a8ZoMXRshJVx
qeIZvRfw5mEP15PBfyrfLe5AuIVQdE954Xzv4Rx1vRc2Cq/GYA1oeeVpgsWcp0lkGPpktzqYLPpf
gI2jafk2maVQsocUWJGxpJQfGQMCHVVdFAPrhmioqlbw8TGjzrtMrWBa4K/uzApVerEG59q1jE7/
nIKZh0XQvk/iq3SdvraokR79N87JVYCGqHs0R/fxLseMQTYr0plAJiCMpeQUiEwZiHu6WwCfSnib
VAbMx881TS1Cl1DxZhgtYyYYx2f0nRqpPvWPjtYCF3nW3pq6BqWHiGLpD7jtUkDqvmguVNZku8me
7/ukjO9roCMyYmemgn5O9gcb6EMfS7/MluRcJYws4xJEK4e/eaaAtyWFi/HSJHIbzj9F4Ry3Yr7M
aNtj2QLPR4GEgbV0dQlFJ67QKeeAz4Pmo4Y/oBPZssQXqxU/kMCLqAV7NTghZuFOpy25cwn1nnZ+
gwYQZbagFM4Hr3L+nvHBwzqx7m9GJjnxMhMBluZ8U3cIz+AUTe89KcGk0hOzRWSla5yv52DGbrJg
AYqkGt8PpI3z7jh/VYFzly4dlHLzbVOiRIa566SfzRMAnpeE1w8cJjW/FSOyOTgV6Ikz5Q6qr2Tc
fWr6Hb3I8DPCkVXHLNn+iuB54W5NKCVZjMKhEhvaxeMjFFhZ7le0ErK2qHewiuDJ0rCjLX6SbCdp
XzPXHbldmxjdDqbkXCkQ9jobim3UA/MBrCDH1Kgb1TUl5owztcMxJnuEjvUMd3SccKSFr1KKMAFm
bWddEO0Vg/fMr3cNuD3tFZH5Db0n5a/uR54XhfsNLBxwKFAb4ej711/tEm/rHXZ39FEl8vqbVDDo
OA8Ri0pguiPXIRK8IlnBB6ynuBR2TOsVn6qGSjox/W3bxgHyF+kAjOFg9i+K6dlKi1iqPWR6I6z5
ePsnYmyIEHe0TqXC/cSG1imjq3+0T0JkG7eQ+ayU4Dp8uu3E+Qf+i5JoZ1PUae/yZ59TtPhPZqMn
YWKqwBGSfkFdrsSVwVdbBBelbWabEyLt8zYsySGkjNMUEVutXA33akCEzFuqiqCCiVu08oNg9NWZ
dP7ZGTSoysrrWYD2Lc9q6Yh5RQ+CiDsqy5EYujcyjG9QLqdFnyXZWQNIjNzcoQnj0JsBTVt/aSQZ
LbK+jitma6jVLlf6L0SUFGJvXJ0pEakvK3Yz0nbbxqK/hR+ffKUWjxsy2363bEJh6ifYhmDGOVtu
hsfgFoqTdyg1g3M+9tIS11Ge+C1nT5PB3uZiQETe7fC/boIWiO00rqYhEtTqlOCBv1vBMv4gtVVO
kHvPZTaDYH5L+yNK/nYV02kEVuli10dQuTmLryeZEYTiWXPVIpbAhG36uUxefxNbbpjrkRuQ754X
wcNH0zzZSkXiszp88tfjkTixNDwGlqpaTmdPGqbnbdsO7lhKr6I4h0riKeqmA+P6Uv94hZA9Vy1/
ENOcr9cE/JMnr4TWD3Z9fZR72emDHUtqOt2XLqXTgQDJi8b2zMdGScv8sp9RAqholMQ/YOisYWfN
vKrf6Az+0jS1ryEs1Ak8ZB/SukiS1VDqFYdO0xZbMnMDGOfVt8IiWlxoySygRWFBHFe+zjA0qvs4
cN6E7tAEJcUFL5XmlVefCK7+uVEejQTg2rsGIgTQMmHBTcdoqQVG8W5YH9x50y9qvBk0UDu2sw1u
lfynySasWPjdZq2UDElKrfq7sNtLNcVz3OGDKIBrsNRIpayd3I1t4my7h+DJgvZ/V7eh5wG+umST
CxfP66hVjNCt7l+00joenRNOICCfgsBQbadKnbg/E/VgHmFBv6XfYiK0C6oXzZyfccO+EJrNFR0r
RnvDrbrvHSi8AiKVk1HphaTJGx8nH0XDQ7q+mC1rP/YPOY9vAnXJYUrlqLfGCmOqCUUlddh4Ucg7
bbPwvi6Epp/vY4Yp2vFy9sayl3ocoZjL1NdYXfzdacWqN3oGZiTWOatiqJQenGCWFJrZNGW1AlQx
SklNPWuk+OOkiQXM3wbCzitVc07AS3804modU2n0urELgRaleaYEeBpks5X0ccMTreeTCRZ/tNAh
oC6p6UWnwXkuGSRE3gu5otSGeEkIcIL1HjhgP7JEz7pMrrrsx3H0ZViy486gY7IBxgaZkAyzCJhm
akY2LduO2q4yQcfOmMVpEGAXtiEksnDrjkc+n6z3J5fJm51NSwaanFQ8TYwuxg2Y9iSArnOocRu5
zMw01QP6tbBvv3fpyO4j9csv7+mPhaeCL4gRzuGlHeC9satKY+nafng3ot2gd/2m+IkyiY1xqlqB
p7n94HOLoLEOw9m6lhT5YeCe9iBvkGGeHRCIZQGmDS5k1TJFiT6oUUmTC4SY5yK8bw46LzoB84mK
os0+hgI1ICgUH2ai7kOfmJ1MFYW8eNBehjcLkyxt4LQSwDAxlnAsZVpASOJiQczXH9CUcqI6D/EI
DC2SAkaNyTBTokkz+TTyeeYXbeQ5KdYL6hRKnL/9cvSe6s/iqjnowlfe0UKQ9VHlVlnBZhH6OSpm
lCQ+b49UjlsJwyMXmYD4ytX3mL18FaAqMPFJio+a45s9niy1SGq7KfhFEMK3weru49DI0ohABuzk
8XbU+KIqdq32SuyJ30e3LRjGRxS2kBaWeUrHcdmcyILeob72j0OctotFr38aEbdGa3KdGpKfk76r
xeVOxn3lET94ZWtB9Px5ZHSwEOzyuMXbrvS6IRXeQXriM6HPsLc3759YvTUcHR6y0nCgPuJM6+96
9xp43NouPZK9vm0FqW6zTA7vS5QK7XKM+SeWX/rwgGlpJKt3W64hWPOcJ+bvkM/frj8BLfFPa4QB
g7q3hi0BgNI2Uqonu38MhNyaz55A58HzmGZhpZTU2iSDIR18WAwSlZAFO0SVKVBdgz+Tvf8SjIn7
H6IqMuyKzQw7vcMzQ7gtcWSRnlVXq/ALUoLklJ/PJj+gyUGITo22ssTIYzm6fSVnsuSxGA4xMbwS
8CgpeP1KmziEXDIGwcCmiK8XVdTTR+WvC3fiIgRT/c3xoPgjCf7K2XZJVOW0tGP03RWh65AXzyT0
m5LhAiGAGT75x/jV3mW1zHHbH5FmhF2ZmwTtaWkGWHGo4Xu8xZ7nI9pUNP9Znmwq8TnDFAX9T8O7
7xsLmUXqNeYx1urFWWL7G0qGHIkyl1+JZjLyGuHCP4FiqLmWX8hqlNtEG1uBqNShQ0mcUOQ1jpDt
y6UYdkD0VmNNYmeFGGS6H8gZ/e6btCqCPCK7jroq+o+oz/jeFPZU3oOPNdHkop4B/NiVDyLscSLB
5pcYzj7RWqQEGP8HDStEhSgI1JRHWJRWaGO/t2AdJM/2Rc2i2CT5+Noj/NVC4kUZV/5m6UNrLZD+
YMEISp0EQEtKLV7IcMPi4iPZndaMGDa0TPnUheXk6G/YF20fbnkCGJ5nbx59KgBN0gQpJgQfKu/H
aprTHmnmZdR8rQ5VF4Fh1mcMn65v28h9xXNYKY81PVcIAdProxWivRHw81UGuGdZPjpFgIr7uFEA
Oyf5uiTa7KIozlDYOW8FJWG7M/pzCHgkrtyrbHVMqNEK/b1zTtqN9mLTrQAIDu51u3vlx+Oe8P+v
xnn8AP1qFY3GOpaPsYwlMZRSyBZ0JJ/lsgkpo/AiSBIfS9O3ytl+ZPMVHHwKGzSnmIB1pDzWD8jm
6x0X3SAqDnMy3002Yzez7GJn8P8ZNH5QDsq/y88ldEA6GQeV4ofCNa7awI/X+/MfhVUvyT5ac1jo
Qs4OMfQ/X9pG1gFhVKvJiMPzOJlNlev9mI0icyhN6OQe7sg/qL0rXddlFSeh6puYOFPulpE2HDVQ
Oxezfwn0tB4Ykb2BYyhL5hudHXlfWf69qSAI5YO/SyC6Bse/NJ45qlnnGxlg1TgKGBjn38dgG8r5
nfCWvVUBA3jm05TmD5UJJOgaoyVYosI4MkEAKhvmAjwVhnhtTpUPQfkNsc8vq2E+QuKD6srHB3B6
tIRP16K3Sqt0EFB3qcjcjEUNRd1flwDJ/NEXDjsIkjoFhtyfcdDw/e3yYxSvhSBcNBIZRweEjnUA
GAhH4yiiSDUm8LXPTPqT7xaaF9PHcTqxCsNkrNLjlvurE5R0ibdHxJu/g71Thcu1cwQKagXAl9ob
LzExDi5s5Oizlp1ntV7DAvgyrJqGGFF8gAgGnLOh9/sbfPhpb87cl2QZQQMKynPW8Epl7e+d2UUk
lbMa08RyFZoRp7jEdaKUhVE5biyUSuwqXXIfWbwjcnJpDFyK9/3dt7yXZOf+Qj6ddoNJIQZLdrVO
AjBM9S/dixsX5+qYz9oGAAkzZs7wRpYnkZCTnCySmCc2uwXQBM+POMeC0YihH2VJlQI7pQuw06zJ
PAr2hVpv2YtKPtimchHFvKLhryqnDqC56HbLqhXhsNWS6P9No9o3UxY5v+aKWF3lHj2hvWrZWnwl
W41/6Jg8qYj/WKFjzl00QacFliOyYEXXq/GD2HdqhHFRf9LJy7odrQkEFK2WIfgQhVjKCNXegetW
HgQ+YNC8ep1c56pWe0PVp+AHii6vIWFiCi982ZaN6Q+rcqUv+gcKVQWDB8rbSqVm12fx0gsIoXme
gs4wehWaKUMlTJVrzghsNi26/mJ+o8r0Pb489JqusvDhwAtZmGzu58clD1znwOX9dHvbPC96uXm3
5OxnXLGOU5ImfPnE5aeD/IiL7L6RlG0VOPjfZt/nXP7Dpil593NTJo1yLl/3N1R1eIZs2Z09tZHD
7cWPJxggYcyzVG4C3YIE2RmVqnlLNUQMDvsiF4A1RIt2a1wWGGL9nGlFplj8esXwuW3EuivoBR4d
RMWSqPsqXNRmXR/+I7NYu4CTdFM0XQXs9OVblfjvRHapM8WoH3fPMz1qvXbzHKx8kgoqfyrBePsI
QTsGL0AEotJjPalm64UKUpZ60bgn3dFPp+cAzSnuhv5Mrfunl378fwTXCG4mniIPN118ri7VcIj9
hGhEiFgTiHVP9QJwKktTA8yQ367umrnU7xkju+NFq4heFUZ9ArZz0I0vjA+eTSg6djSnt1KytXgO
mTBioh7B+WTnW/lK89wtTllA+fXKZzZGe5Z8Qc8Wqv+QlTA5jU8J2nnm4cmRqKwUhlOfJ3oGkcei
+UgWPIcysWOR1CC4om6l1Slc5PEzqAFZYM1EAq7eY2Uh1c+PyMJ2uiXaf6CtpfcTGgIPEGiUFoLe
On7JrvLNUC/zco4E/3nXQN2Yc92BTuzLS/oSTo5N7V2BftEpWTxC5Wxuj96MQoLeIP/cfZw4vrro
aLb989wuBT6EEXn0C6XaBRe0ke+RJEK0Ukq3jLBAbPvTQ1/bJIo/oCbogDvC74Dev6R4B6/+7XLl
kOU/FaeYg2ERHmKHFMF4URazK3uxFrO+BFd1NzEzuE7sIoWLraTYnfjqpc9TRoBSz3GO2BbxBLab
/LhQE+32mjXZ1JEB3X+obkbIAea7e8M5SwQXJI+sVSOVuqKotnANS2bTMICrHKK4O2+KVSIMB17C
wIc0nOPPftzmYh4UmbvgjlJXlLRi6jqQWxUcSQ+FYKFb3XOuy/N5bvWbRSp7rJT1qemTMh/MvzfQ
4PPDAN210vK2iE/AfaHkPx4MbtSfVVHUfuKODHgxYfhr07U9oUkjAIELh13I+P4SucJK5HUXctDn
6aijxycTADKMAzpN9ehsV8Wrvh3I6lh3A6P4UzPO0S7zulvAINgj+l7mxUY1calBmtGbXIAZEv0j
TcWToZ1qxjSmZMoD8LWFxETx+qt0q0iy+TcpnRBDGxWU6pYPqWn5SWwUOmpeKvVK0S6ZkMcXxmP0
y+6M8u5kDP3YIe8CLbSOwYCz8Zm9Cx5PlVQJzuZ1RCey7b2qOLEgf9Iaj5ywo/keBlDyNTy8fc2w
vYU2xLS+d7ULHPydDuUgewUZVJRKhlt+T5wqy7hhUlVJzYA83RedC3MTF8UAfCIFyM8Z/yggeeus
uJKggy6w/DgAIGgvUrTCwYKU1ZJdza4ah1PwW8+/udd0iklc6syRE0qFwqlUmK/81R8TBLkvC46O
5SgPdKW+dfLvQcuZnFWiurDDjcD7Y/ZdHYxMeMPi8g6Gjsu+s1jAVZ35J4UQxnQUfq0nT5y0OxoR
K1w3x+xnQ1QFUQMVjI81nYHptbeUjU0XfPocszkuTQ15p2+78Zl+8SEeGeCXaADUfbODKO3UcuWz
8gpY+m7SU0D5Rau2bzDO3ZqjAg35EB2j4a9ctv8YUQmHZVQvTk90sBr24SnVa+9wnYgOyffjXaps
7hWrSk3dXFaW2KHzc1AhskEaj3wMlv6XlKACXRzPQXTlGFo+1uE8yPuC1aNUCSsEr55x8PgRhsKH
sJ50jqWuchUlMJUqsHEnRYg/naI9+qPMrzW5zfVclE5Ufjf7AiIggy4JCgoaR/J+cu1+/tBTBei0
6IWQtOwscv8kShu/weSzLkwgn3yTckfjNbB1JBoebotbxqmf9F2gK09sExXbLcoEPaPqEUmZunIL
Q4x/T88DcXcWVwXlKq45oAlg8nhXJO4tm9Nebf3k7jelHq1sGh9bdh6NHq0tzsyeJWFQnPyXSA2l
2RTN+oJH0NF0zWZdBQXsgV1o2Zj2hteQQD/AH5FObdFueUNxRCvBbpC3zzsbRzJbpN5h0/2KJP/P
8z+zt5x+bbaocYBSfBe/PBRFhqUkCkV6AjfmBivPG/FAFxusfily7/VVWv0rc1ErvDHoB18RaPc1
UYrsa+fSffNJLIjbYl2jZ9JR6xiRFG0AAKU0LQAgYenD9ASUfzpq3nbYTyB4cqUOTpnm7ADcnUQa
r5FQMveLBqeO7t3wbnblqF27cL7rVugf7I4QhS4REsm5EFHlcBFVMuB+uMngnckfHdWM4tnN7eyE
yfJ5KE0IXCd/hd3+IA7jvckY57d+vPh92wyFsM6L0Lr8yeD70+PudVf572Vg9PYYyEZ14vvJLb51
VpdloBanMnCMMyZ5oFYfne/2NreUfq33IUsxTqpMUdx0ayB+mk/d3RZ5lQB+/FzKMFGdc/1ZG9rm
bM1KQ/2DqOCUpUKze00RojJv5IWOI50/UvsSgCdvCVr3ECFQ4es+ZQ9GpMynI24ZKiYKNpl8ZG4B
4AnQRuGnDTfGWODheLsBux/ahBl+1DqnQDNHOUWYFlj6HL23TwyIwViSn3wTtftBR4eqSrlNAHQ8
PSW834foqjVbgVvNj/wpGV3n4Te4GbzPs0KecuCgoPObWmyWsr8n1ceMxB4KTGzBBtT0xwhJzFHo
+2gswybgCGZ71dEop6ywdqcqbueFytXolx32mTFheCWPEIPTJ+FC76Lj9bcrgnPkMpJ4a8/stvMA
GlCgmFTGiHsdrz0HEFSwRTw9+OoJpRZpIIkDW444kKZxeP5LG4GiUfCgeUykZOst7tSXdAnYcvbx
b1GOolnFjk7XWGnYTRAfARcviaV8xgZgWPiv150HzE55NI2pAV40dmIw/K2WF7nZe71+HaaPXZ6y
gecuoQsQtzvBkUiOuhUPgvs6B1uAICOS6FD58sRoJZT+PTGQtgKwIqADAclMlBzCSCBFeQjfqUue
LZaUTfzjMmiRo15lMRnzZVQRJPAeIevtYZ8JQq7fXp4r+nbPx2oN+tXGcuff+ORVKSc0XxM2c+L5
ZlXMnk5tLeWrabURDB4qAZRq9jQrIFv3v/sGFMAGB0je/oNRJS3waz/jvIzzbr4EaRejDg7Ql8cn
X/PjRLr01cOP5vKOkrfix2hgJ8zR6LpBXWQyd1aWhy2farkMrbMRM49OACjwKh01dMSl2MGG6qba
llh1mK4g3S5cA+FQW3vvHes+17/3kAMZRZf6MeN5WxpmFaxUesjy/Iw9pgGtD3pz02IzjiQR2uSj
wkXx7NGMch66R0ynrPkmzCmxemRmVBiaQ1UYqCZXjQvP1xuUf6zX5V4n6qJ3LsFsrYnrXh3ir784
QtoEYOON7FCZVOPfwDeIE4U1fQDNZs6CzZe0gF8V7T+rXqayXl+JnnnsZOAnbm1pi1fk1yAn+ZXx
p7+1aB0NPVbA5UQkJs730yl0VQbXwpRy2kzV1l94gWBCE3RJ1KjLD5aLZdak/k+K/c+R1BYUaGvy
XKIxK/D08vMPz5/01zbxMtvec3i9fVQgkdwya2Bt/r4wUJbnj1+3hIpWmiLVwf03kVlFFqHPuQ0T
aBp8BwArCSMyjwr/eGeywg5rFemgBp1CXAqQJE3fIo2iXjNaIOGxJ6Mf2c4Zpf4JdH5WKqZvFIjN
LuYMxBXrbIGh7tV0AHWKmKKym8j6ElSdmhpO7VFRXcE5YXK3QqCidpcwwZMAJK94rpdBI6FvsexE
HSe3tRNuiXxy/Ci32PBy7UFXQCo/HZo0Y0rbuwGgEcm/WfvN/ishDXmN7Wp7IStyrJuRrR7OPSIX
RB7M0C6NKx1pmfv4fzu/ZJhRN1YLgnE/HXvzQpy4I5yysGg3P3PVlPluIpDMlH/hngJ05TdkkSm0
9IYTaj4WAHJJ+qWlX5lc/yTjr0uBGENwelz0W9dqlPS5h3QeX30z0k/zoGEDlXbBWkFRRw1LG9zH
kj1OzaQ0rJ3kkIimYOdDzvKT8U+IH0EgHHpNRl4B/UQvoYuBEaXni4aCWPRmSSROTaA6mQWWVREK
dFyJutN/uuZS5bM2U1q65j1YZtFNK/XKIelE2+HtR2EgkkGVloX3uUqpCw8X0lQLJZq/gx5fe5sW
s+09lH7GQOGjbJMZEp70LR27E/tFNs3tLnifblHQ0GNQ3LyikCFFhnEBbW/wNjOBjBa+2g4OSfat
wBTnfR1OmEQEj7eNi2TKEGRl3ukSnTBNxXhqB82PTKItC84a/F5KfdBqDS4877q6ynD5+wvzeKXM
/CREZK+glmhCRbguXXN5889okn665FWdX0asSRl9BQQtVTsqxPr7wEzDT7191j8133DGXldmdCAh
0R+nuQDCqI21jNCLYAJ2h6q0Mb725G475HNlLyrdxf9vzx3WjhAc7806MgnBsHGpK35IoAngbo6i
caaSZWiGgpKVa6emPjwzYQCycRCPc9wclJ0Ove8Uzf/aYQoWN8xuSZmsPcj6OhHCP/zizRm9nIWj
fAlU2rrGqENSbHsve2aWANvbqUBC0HXyk/htDphx4MEyz79UF9PDkanAE0+/0s1wXju6ZpYTR9hq
QtjXcMB93dOb7i222eo4vLox6q/YyW8AoP8Pc13HqhAnf0Ardj1CVDtaATdsycLiEygtsNAue2Vl
AlW+KPyNqka42GHc9pSPdskF+1nXiyjIo8ZfUE3czDv4TpfeHZuwJVZlaY/MHrWuVm+jwukABm8+
7NDbg8P1WsKt+WRfp0Wj28gfy18ZFCpVBVxn+tKhS3l3Ab+n9MFpLBwIbxPR00rdTMyiqvLt4VFo
JdTGnASzZyJFgAoIMD8en7UaPsIKGi8hH52bXcFWalM2XEAsmYxQp82HpDKkx+Ip08yBlHGrUmjd
VCz9Y7IOvR3Oag8lIxt57Y9ovISAUc2cdhvNd8s1QAzf+/B9K5Tlbuzz4s5IBYCvji0x+tYRjh3Y
y3FBMBJqS9YjWB1AvXxasy0NcssfSbnNjujfk/lq/+QCdRNpnA0bLiWfLiFSnKpbpXDDjtA/Q7A9
eaq0xj6PsDdepYSFuzXDY1QPzrn38nRzhmJNSu9AnXizVzakqB65Yx4FkzzTbgOd5hO3hFGpn7Bd
NB71QqIKWTho/iZcA71s+HzZZhOs3cBAGYT3GCzhLa9+CmmJzI6unVl8wPM12e/7GaYVv5uGBz/n
TvnzIRFQVYNze7XE98A7UFqtmNR4Rxvb2B1vKEktJqfxyJ2f7gtZL4Z2ObVkPMbKF3PymlyM7hdq
0pQNHXXaFkApDuXm/OoEHLLssQqRsX+v209WrXJ6WOYdyywiD68CapnB/nu/RZM3ZPGdBAUF3B0p
69/zYu9jU/JO9zPwIiBWkyT+lGS0Mmt6JpHjtsS9ML5vWR0KZoFQqlKUqnTDKaJ/yqzTrTVf59bH
g5D3M8NbJqvmJP9erq6Oxaaz9EHwdzhh4eZLF9V8OdL1F6zoYOY+U5O5grV8WrC2MLxSlyf9puaA
uwy6SgtBf67LvVR0ntAwtE6Z4RigfyU+VQydJZ0aiYKBOTi77qN3AgnKrCWwUq0BSsCgFi3Y4BGK
3ivFjRV4e2uQXp9tZmFgphBxPsy7OQh3/LAK23cvCwrsXDvNAS4TFHO6NNAq0+KPenjQa39BUneN
5DmIAdQLlLfywfWrBSGIHI0Ij+mkmbqm48wXpSNAbDWhqz27X+kBuCNspzmA8IVhHskIZ2A5jrXx
n8PchLLyNsU9NIhg9XhKim+QV3wgJ5d07diSjXNayfC78Qk5icAnw4rYh3i9VqFTSPBxtSPiaop4
b0ttKqLjUHWW7+K0heGWHJ0r4kK0M8hcyQ6s3kfPxNzQuoroY8p3RnMut1WqW+oEIV3+ZuJou1bL
DVuDUzeRl/7ybS4jSD+xds91dH5zBnjJ4xWYQ4vR1hTkPuwVkmJa2xWCyil2HKXML3fdhPnrNljn
Jp+jYxlvOesYOcO+jNYSK1rC1bU+UhMAi4a4wTZUAS/eJo8ke47Zlv0fepK6NShU6ii2MKwTY5VT
XGJ6EicVIE3Xij73d+RpU11tSoSu36YDT6YjXeMBlVbi2SMpzDAZSnU/kXq1mlSUZsqF8WeiPiB3
igLbHcZlZHKuY4n3ihds3zIi7VFzqg9PYt362M/X94x6Jfot8eo5dO93oHfzkY/iw4fxHV0Qsd8R
16+iOVLdKJgEPY4gGnqmI1Ufl9nyIU6mNcDuoc5mgYQPa3vpvFlveXZDbvPAEBlvjr0UiGSgxv0H
jeJ5HK5YSKv4/gzPEeGmUbPiH1qJxiDrLOQAl39IHmo4BZ3+KMxMV7s96GmW3XB6GJAGmovZpJYT
BuDQbqWGpazk/RSCqjTpMv9T9kquUeCFjgGXWWqwT4L9ONFy98iKNqIXE0wbLrlWVFbCXfTAykrX
4rUXcUdMdaYHU2Oy6WGp7sze9qOGNymbc4h1vK08KErJLtcxiCGvzcvGkoTuIUatlmYTW3SNv9/v
chLVev+KlutKSs0QO91BBfR/ICYdQO5z+i93Y0EyP/U7bA3PWCHkBNShaKyzPR8a6MaZGcvAYvdH
Qaz3fO3JyvgiOoN9+Z41oMIaq61xJsUN7eQjiESfsaCdqWCQF8z2awbdPWwlF2aj9O/8/T9MY9DG
uoNah9h20tgsvBZrL1ygbiUEHwX4DfKiMexGKFjlFXVGSgHblin3n40NJwakVY8H/5YKixYXfngr
lcXLVyXeYr09ZuLjVs1t3Vm6QnJcviwKDCPsnWqougIWvK+RtYaJ+61ZiDAfSd7/VCS71rtTRrHZ
/fxxyyToMwd1ZT92S3pbb/GNZX9qk7frm+MBH1wbmCC4Ya6EJS1iIdfqYn0ZVCCB+OU9/V3efDXa
ND0ac79N5g/NjgsZL8lSe7P1di6Ei+pJmnQNepYTt0OSSg/d2HLwm+kn96XwD/ReCoSlvFzpVaf6
BJnFiFQOF0eqV4Avz7pQlHv12U058M/Hyj2TqSw45z6oTFBBEazo5EsK/N9EJ10JPeXk5b7dyeyY
lbMDDA/rHKsOkAWRh9KH49CkOiSCtprTQSW0kYW3sTx7kLzIYFXgoSlq3Kf4WIwXEzuhFvOacdBJ
Q4Is0963wZVnWtebzJ3SxV52qlS+miY26IgmC02KdI83hXnbDGq20Ed+MQVsa/bu2j9O0doqAXUF
MDiQmqYEXdZ5RvgDbElSDTeB1rwdB4qwfzw2GbvuWw6m1zvVVH0nehcp6rBC8YamAMcJOdzWmSue
anZHSZAVEk4dGHN1J1k1fXqJhDa0nYFanRiNH2gNauzXuSmBRXadSu+Y666j+v9rFrvkkh7kMmq1
BARRSblRBvTs5q6iEaRjgg0wLE6yPtM0OfJmyJazbr11O19KWYxwszmXH90Lsg850krpyPHcjfE1
nF551fEYkWgt1ETqZ/hl8czOrjLLSyEDK+e6jeB1FMFiL1miq1SyeNZ8bynzf4CglfgRr/Cq4xB4
nsc50f9mvDzaB0zcl8puviw17z1hxu4kiYoYEmOCJhcgl52MEWM1UveSbk+rLluzIT61uQ+irtEj
sR4hZ7I34OFKRPgcmQxJ8LznGq3DjkLlE/shmFRNiIudnRll9qTk8VsJNVg0PiyDN+Uj6BBWSIel
mw80099MzpWsnJJA4WavDQ8t0CKKHqRBAClF6/H2JgBac99v4b8PfCwZf7HsE46dDlV9hiwnHJx8
18/rmJLpKH/W9fnC/HBBbyqcmzt3LnizKc+WT8qaZxzSo+rZ9HXSOugf2DsmMQlw4h+H1S5Bd3Rt
4m6ctKlFiBd19aYs4MUa9tDXOG/OWeRTJ4USXSzjbiZHt6TGhnQc/tAtznjNWANPdAxDIIGH+T/x
Q+eq9B0QsIoGfIhocllvOElC2jbYG2QADRxYVdbGvnoW8Tyzx+abjwXyQEu3raQjuhfMOBA2Zl5u
8bPIH+Wd/nVSl8IdyEoJ9a0jCZ1ZlSEFWf93aYmWHmWdBsnhSBR7+o/3MIolY5VlRYBHOIfUXKXE
5EjvlLRAPDkLv0CTX3ZozeIeBX5IEjzB2gNKR9bjfwffxz1i7uLcRrXquu0bGB7R+HSeXvgLcvWh
jR0d2jRt2xr7mU0QbV7e2erN33gsg4Zbzx2Iz8a4ptZ/D6Y3ccVKWPVMWHFQry9e3MQl9Iubil7N
+yw84HUzK39vY1j9dZTn+ch381ZrSSA+nKKlLkeqo4r9CJPw9YJqrcn2x3/3DQa1ND/VNnkO9V63
VGLvyMkCuFv4l57Xoxq0see6DqcIXcSAjeStetdnbQ0QS43j91NF5rHF7d67bYMeGdrpSVfmsSQv
rvsgXkSu96dcVJn2gMBmBc0kO/wdBjKqJKE+xjCmQ9SA6fQTbyVptCsoI1U+oqMY87UR9w0OrKPK
gME+bSm0g1bNw5q2Cytpv2JU3G+rs+CNjg2fz1MqVQnB5k2CunjNh9xrVQ3Zc5KSTEuDHDsFIFUN
+jCLS4xEGbZCKLADVU35xK6KA7Mk+QuD11MsSvFjfJUyHlsYPjjRGDxSW5YIXJzqCu8b+9+fa84H
6I9nviIjfduKvml/yQ7DReN8WkCm5HlHpORo5LKgQ9Aiab9DiUPe+L1h80hUEiYT8foCT9TpUYB3
jTrvNBOPhXYGRgPd12u1zIvfRRh4nU7nfrvxE0prfoYMLRMiLQQ4WafJW1rnAJ3O+BB1TZv3Nd11
+wLsl9+n6IKanaO3hllwrznVL/FdLPILyP/gNzu3QJ2gVDw/qyX7LscmTEeY/WEHGNBkm/4iEnvm
qsAiTsysxSZiwaj+48fnkiroGgL+GNfpQXSInlOZBBM/81rnmCaUqDmhmopwp0Zu+R+ftdaqLcuZ
jSeJpZLSzBPG2uExD9Fx/hDo8ZA1h4vYB8MFUOFEwjvZXG5HB3XGMOX3mleeR+ym6HViFCMhRyRx
RVsylxI6Ya8y4NBaa9d2GF2At6Dru24KMpb5P+dRtM8EaN9OH6vO9JlnV0NJh+k5IweupezTFXMH
Yd0jbL80zBr3EQza1DyO9yqNyaIoCDW7rj4F4JwP1my2ZuwpaFubFKJz+lm6USZlJOT1sc+v4OXU
OQzT3D9kN6BPry58zRiHln4IeXHEjCvJnLL4iBCS+SkrEiUyCDTjBqDICqIRKrqWuHFhLrztg2NX
FIbuAN1JD0L9TjWZjpZy+L/Ow4B+5tt9X7ssKIQweA1t8ZoG14hWNuJWQEd7tAaOPKxw2dgz4Hr+
JOEr7ELWQ6n2YZYNcMTP3ENzWF2wKyMm/eO9e5RUlqtAs8biBfJCxvFSU8WlYCYS//vDOwk1/2TB
3GsLS+01hsSM9RXL/Yduni0l6S9QSGxG8IohDY1BENYT5CM3bxjhGHuK8ZJIDU84PXATiyJtuKf6
jTE45CGEl3BIsXNfeTmTm1++tI2yrUPg6RaEtJ8U2/Jq2k8yV/Xx9Jxbh++KlcPYRE7yR5FbQGyw
J1pwSfNTPg81V4+K4pF8XMGpZjFm2m6mcUSMuUO/oEZLx4wpv8cgF80PI0fkJeEdSlJXhBr2L6m3
cPAMk9OrUCKaTMGREbmjS+sCko/aNmFioFdJHIux0F0CG0Ios6AS9Fmt1jHFHoYD9P1AmdN+mFiT
GaDxxFek0zz1I1lafb9WMu6rvH9Cu3wT0vGGZ8wrJAIRXkP+5Qcl71m/rmqm18CYkdoco6svnSGp
G8FPaAcoRnrZTWp4P1+ZKj1Z2kqAnZ5pHnCkrRyYp85EHspZRsDloDhVQCR+s3ucR1RluhhNOZGr
yTm/r+b2edo+VtRVjhstoPM6sMRijymJBwYgt0cGDz5H/FMsRX85Feu/mEkHNZYimXCVIUS2IiCC
NI0u/Ec9Z/upNn1clcsWQDwzPB3sImTRY8h6riSUDCacP3TnVCBiEuIlWbV/8OGloZFQ7sEvdwSc
oJzPcb3fDcyPd2Y9Sr9EJLVsaeohvW2y7bRymCJOQyOY/9ohNR+hHYmY19/iUeZBnJOhwAvXsAwy
+NF+sXufxs7Kklo8gBI694P+KoCKmC2DY8u3F77xQCMQwQmsbn1E1T6K/5OuZjKHpobr0jswrglX
T4X6ZbnimmqBIF4+Dec82AKqihkEjtaG6GldFmavvfJaC/8al2bCPrtycR3H0qNnANB6CauJtcdt
z/5d6mORLVp1dWLJ8GEuFPg2jAEYiCM0Bjww7B1lbcCqybcutkU9TF7YN6BBC/Q6V/FcvW9HCAyR
AdomVzf+XH4x9eqD2TtROZji/wUWeVU/d5O/SK0JA9ff0aAKGj31dHAz7hIFaWJ5GP1tQj0kC9Wl
JuVHYjNfOYXFsIpWcELr8ONod6Wf6aNyZ2DZSQ9NE76aWn3/03EI6HfblZNCjGlJx93DbKgUY/W/
03Lr0FW9z5ZtMOREe+3ARzyIFbVaIaeHSg6USpVIaYW8+h6/XtIEGtgVGRrjSMCpelMjfpIsoxni
3YGnJrS+HdarSixrXSIv37CC5xtZPkkOj8AYlyt9kIouzTYni8rkTHWgcOO/XPdxCUArI4D2Mpid
+o0SgRpzu2RbRnlCf52AH+RgauXeEpHkQLAZOjj7WJhglUMYs4/vv4g5q8qxbpVg6Ip5l0ea0rIg
B7IBrrZ669G+fv7h5QPffbZCCeN5bn5lzLwJ+8qNYJeMgz9InJCA1N24yM8umzx8kNd9k7UlN8B+
F0havbOZ0uaDdP6n6WhlsVD2Ws3ZaWIh6F04+FeDQQvtm8EMk6PHL+kzGJ+0/pb5YaAKcDWhgfeX
VWRX66tLX7d+flZT+cCb9iMCvel6Z/nN4C3f8GsJkQaj5FtXoUVEv1J+mEn4LcBdEksaoSjvr4Bt
8TTv3Fd3PXN2vvvr2mQp5Uf8rh67LQIo7C1Fd9NbJslzcqWY+z6srVNv8DvsnAx5ZJ/QJU3Jg1UJ
DXSNLibsYAWpW4WDeGFuxDfDq+oXLGwY5rZNPAe6OJjA6Mnh1uRtXhBeaI4rF6frCMVse+xKVdQx
MJM8fC1twNfIcvAayruHt/cF2SjbLir+Pz8UUUOIPuTka3RufvYzT/INKzn3iiKMh/PIgiAkDDLk
J2tVmr7VsFQbbMjN04hDaxJrKxOzUJEvazpSBJbRv2WIeXM52IfY5QOrNlXHYncocL0kWEHt/UGy
CQZ8tOvBxDRoIuSrFBnbRG/D4l/PGRDr/8x1twrVPwOUX65tefWbciaizloXza7NWUz3ukJvQ9f/
ByEIE2l6k1cQayzh9pof6xuNoDZDWUEKRyCzqRMXx57pySkA0pQgy8DPq0qD/g5yD52ofavTs0AT
mzPZEfu+sVTMlQIKoupF59tRLmsQ1UDWWyAGI4KIK62J8VWAO3DP6dg+7CKks/tMDruDISVBvWEj
Lm6rmqwnh0dXzBNk1PtSEK1WllLPnn4OEaj3KTH5hV9XP7D6EySHufQ2rNJP5UlV1SVIfOxxRSgH
NULqQgj8WL9DjfZQxTZx2g8OLJXcK2h9LOqXRgjJIZ1SS/lWmYn96I+3ow/BkJDU4f0fxXEyhmAX
a86z/6fVm4zoy2g6wiBl3VXqpK6YEAB8pc2FJnM9ZHVRaJIMghjWFEM/65RiumTqVkUkpkgDb96d
C3QR4Jk4/utxHQ0CJXz0lfXOyboUgsXnwNjxEasxHjNNolZeYMSXYJaDSWz7cNhVyopPXbBwqaxI
EjcG/sKPyvTraQWduTI6yC7iOG0ua6bGILnjPWzltQ8D5MsszxYgNn9N/BHjSyIeJ1U/0wZWnWMt
G/Uhb7C0hq6XeAg3dQqQOnPVl5VQAS4+EZQA5KUNlZqVA/5p6P6op0QOUs4c0m+YkfZCvZSjFoF8
xmQmu/oWS/A2bMCBoU/Qq11Um+bVXepLrEc1MDxM3ACRfLIiI44G9DLx0xsu3bIzf+hwfJ+c3PGH
to4IDmZerM7PLig9Qj13FfAdd5wA5hPpXIgOYszo1dMTpXZqhnJdqTteuU/7GtwswIhdRq2konw9
tM0yoFAUNRYnE0EGu3+0COMYH2TkWxPDkw1t6CpCic4Atz8fP0hes9avx5TLFrEQ+h0/qq10usI6
BfJaT804di+noQD6VipPFs1+URJ4teGwO6s6Sl5a7LvF3rayynd8IxEDWaYoyVN3jQ2W6ydIaDkG
xUWdtC4boJUxrwkMH7H0hIDmNm95CKELR6ar5yTlI51ejqG0EPLGwHZdU6lY5BCFAEigZS2JsPGz
z4khiliLbuGjMqhbV2lIKAUnUf4akmr5fX0FReSjDUJKvBl+qZFGQ3EDvUwnjtaFAju7c0e3s5KM
eAvk9GBhnq9BJzhXE4UU/Vjhj3nwagYeXpj/eJoOM2apjnHje7eYpi6pTEf6mqREbs1MzapBDy/r
EPU2rEFOkqMcp9qnlW8ukDDORsi/nCQMW7BtQVNRDFpI+Pc4qy6Rnd93VBT6TKJDYqubBD9ZbD4f
QCerNIXAcPuHuxrO78EUS+fyP/FTFU58Dc4Ozx02uKn7hxOi7qrCKqa0t5wyuvhn15C/gn1mgBeK
GsrSqNOsN7Ie+9mK/YuRI9T4VGIq3DGWms5xO2BYAUUf5xuZTudyDTXT/cJaRPu1S6fDuMpjIEje
uZfFuAusuLs6zY4HP5V/SQPn1/N1OH+dVjZTs0Sh9I6tVkDCJj5Fq8cBDkX1uOT5fXNWle14+wd5
srYvxVZ7VxF6bewz5wuMadgVpsZk7CP6ZLRS27ueSz7+WvvudRFYSGHtVKYhxLtMXjcqqSZtJFNk
JAw9ht7rGOKqRe70Wd3qrOgKRyoX09ubux4JO8JWoRgimzbXLHdeuaZjt4HmZ805xoSMU9EH0clO
sHDaQlBJNfDlm2H93r/KWBH0VG31yITDoGWwQulWZR3D25/NwdUOb7e0+rEE54JNY1VLP81EqyY0
bNfw3EnlCZTJb0o9TElyCJF4nVgh0CygY4hv+ii+FCay/beYGa40m3Ldx7XkCnBEFWn35ExJEXor
QLy31VUqBq8gwPYCaQhT0nuieVQrnrLwEhPgLlxwDuQ0gfNmcXLT0uY/ZyomxKGbyBZdB+3WRo7S
1y0NSChvkDu+aFWGXNl6V9Tp+LFpEtjherrGLar1oxYz1QAXBpeoIVL4LBtxwzyAnQrE0hICERL8
FkxIFsmveEKBApTcQlIpTNjNkka1aCeov+ZyWov+mpy41ESIdOo3o2DrY+7tDaKqO6ltIFUZSMrD
0g3YfUBSEYoevMFkzfsvuMxvPBBrP2S1T9YgEjxpP90YOHs+Oy5ayc3QXqJpflKCB+jfYyhx9e0W
vkBDG25eANGJ+uhafATzJiJVzQqstIl9bBprfNR9iZq5kXgTEdkyZkfD2i0ZXbEQIKyyvWNMu9cB
HVGJbXJ0jxgWoOhwwahu/XaHoUFfICo6JhUHS761nNoWwiK8Lfo1RPi1hZmRsizv6iiGLx28rtCJ
Dc3LtXwSFcQvJkl+uZyUpnwDm5nYoDrN6wr68q5N9Eit4lsSFZOIajkD8oJyAZDRYsBf4VTx9Vam
YAi+hg36wJgWrsej60KYuiUpMBFTw4kDWuLuufDfTy6rPVVOIwaA4obZQvxdWFK/8+WsB0rU0J3J
jlKkARaGM/RIMgr3qJoBTrEWad5PlAvOLExvDazz6r/LnLC+C4VDYTk4S5RAFjjp/cwRwVErf2VS
ya6xz8GrQ7tTarafDYPBqt14e94iBXCO7PTrScBMm8tX6ifJW40wq3FKMC+edivvGghR4nXRXnTM
l5pdZvEIf1c3P/7KMX8M6buB/roKROyIOyq9j3hCi7osK12e5QgrkpZhGHz3rU+gdsEk48zmOe06
6b1RqYCmLWMf0qmVgJ2Ex5J9/BtN07R1Eg/122aTvdZvcPwd9KYPVK5eV3GfwAXjII3SuRMNmG1H
wK8OeRKFGIOqlaqfPfVM9siOYx2/hgqkX4vPzd6nthm0usCK7sP+YMlBNhgim8EHzqHvJ2iTxEqr
S/cNiw1/Jwvbu73VB9eC/7s7y1IDruKiiytzKvIAJDBf9D7AaxXDbnG+nZBKxU8NaonpxBZd9JeD
qR6KePfgFXFKjQKWxB+u/nSi7JXu1YHcoNw4fF/YluLTaUDONiIfIV5Yuz0Zz9l5u5PvHIFpoJY2
4xUkAwV0AQVJY/+qIPz77wcVv9RSk/MOslQBttef2cI8+2l13z7UqD6JLfRrFu+p+rQkFg8miXWW
dWDJGXgmTPWxuACHsacQyFR5cBr5XwunkmaJ9vdnXuHnKNOnakP723meecPpL6Yaajsc0vELp3oP
cgcufHgINffFnxVnxPcaBU7vo2NDpYwWSG67456e7bPaxxsVLxhd6/uND+MXp1uq9R3pZBcLeVgI
5nqvoqGza++0G/4dgvf6yB02m9wV/MtYZs2b5jdhn/u7ISueKp961/TTAZhectavHPQjBC6G2ELp
MvH2Dfjgz5hmYC1Fs+INDz/LmpXteHizow7ZolfnjxNTcEJn5DUPtlO1DNmujt1gePal/zxfJP3Y
M+73BheB9z/DnL+fdUduf91XyuEsA+5eUdHkcjVGsMJ6H+N0jgntNpklPUGH4dEU3oK3kdW3WW1M
7kEZZFKxjo3CpjN9zpIOlTxBfmvuHllXU2tMbvXZLnRXMPGF04aptjp2GaCBu2aQ8S5Atjcun2LP
4zwGJtxEM99ZihwT/QgBpzStrSaTfheUaf7fktQ+9QWDy6ipCc8MS3i14oj/UMAtXnREqhWCSx/C
/ODjccSxywn0LSx1cAHoedwfObju7rvgfn3zRWDylHvByQCSwWWuXND8ii0NW22k/JDjmGhLpRml
AzTb2coqeh+PBKgEdUC+JPyaClJkGiUV4kjLgMN4AqK17bXYZrcvgYBlBD6r1kqEPZBa2W46gDx6
Pvf7tveuy1Nsj/T1FIlDmRbQM0t0Lkn3g0ChoEMaxkpZWXNL38yOcGgc5HzQHvDwZYs4pUX1yiIo
RPigRlQkgZPSu/CdocaWV6aMKiV9tM3PvP2upLHdGq1nMu0m5S+1UCURsCkCjTUgGfUjyFQns7bi
CpZDauWWAB16F101xwOg00K5g4Nt2JpjWmjcCqnFvDEOjZcM1c0ng4OQdGdzByRMytk9GfC/vOpy
mqXM+qNS/w/0EZdjfbUmWJ4VZW+f7z685BQT1Yn3nGmczXa98Ss9a5/kqtzEE0vAdKrWxPZZvYG7
2wM+L14g8ECdlrfxJ75Iy8xbGnKCBwzsD2ZuT1xvVdCtRQd+YQCrZbrImSGhZuSLCGeYjab3sHzb
FarRbGHUxrc7f7ESEy3yky7kJwP/XJsy/vuYvB4wXSv2Yi4UGhzfo0Nmpfc9k6OEuCVyrnIY7OjO
6eFEaY7Qvehoi+V9ieaxtUofoi0WVC7YvBzqtpzNj0D8JQ4KmEz5Yr4GFUsGz+A6kNAwDLRKlmCf
en3H31egG2GdbJ1WYutkDOdbu6/fPU7SB67uDKH7+LsN085KkT/L1TXDBImc8gr6lZG0cDg8ewrg
jg4CjuL8TcyqOl61oCcTIptRf7SL/ONEQ8djDWyhifyuvlqWmwkf9+OEIZbqSqcpqoudibWhHDKd
w8dVexVGEe7CFaQlkZs3gKSN3JxaxV6mH+o/DiRitfFALHidfCn06BJtafAo6rHxRF6AUjJzbBoL
KNBtIhsvFGkAdd48vmcGmcm7hQnWgzNnzDKNDT8EC7gA0sH/dh+hR87XMvy3tZ39DcSaYM86aLkn
PqQC3Htq+VRzkPpfRY5zv7Hj+I88P0J+8SLQf4GdA+qJIMzlLchw1TdoLLpsYS7PPxoEjColAqaj
KyEskU3En6l1yxzIi3fSQNEZ6rlHBYSU/ACdZXNPH+3xKBz540JBP/Lq0iugeBR6wGtKl84+W2tA
N+9OACN/Os4ng/DyKJwzCKILw1qh1zqfEkQfHPtaapMPyQtKV3F5ACUrADkdzQbOu+IsVNWrnN8Y
32H2FwUG1fJUdlBp6CbKz02YeyVTEEWbAMmuqEnynvYleh3enLjupFG38OuJfK8jGYrUBqCpV01q
208r6BtxUS69vMh87Dd7QcSfpd0ied9BapMzcJd2LgMAhrUGMExkj9RbwXL1dv3bJy8obw4kdlK/
Srq75q9grKUWDjSNXWJlZ9GUoNWeSPeb3GaaTEIphbERvnE7bGpmO69jF8zGKq88kAutptlppOEV
yDA93cGmIAf+mItGwS9nKHyRUECu6L6zMuVvs15wK+0stmX0ayn31Zoz6wbmCyrpOqZLkc9RKzin
TfllUCDAJb5DCqSpaZfYj69eql72NA9nuIyCakUgtuCRrRUOFyLI8z+2XXXh/DzIJ053wfEv1kWX
zdeeviqf+kKRz01iwAVwxJYl78ZiR5Y6OpUdu49g6vUzxuiuLsJXitgAdn3aZDE2ly0i4MES9hfh
LqfqqIh+5joBkL2Wt6JFydkQ6jbTRM+/mnzfzhmtiRuhda77F1Drv0CMn0DWL8OGpzFRyk8X3HT3
wVJmBYD8F7t9EOa97BsCP9hsZWnNa4zn2OaBADC3aazO3KH0TBtu53sl/vo+6gDjxVUmIk6rzxXZ
PbciGcbCxfCEQfM99fgFzq7J0mUUysIT7v/Z6NRZlIBX3tZq96nmSvloZsR5ObEa6SvTIHJnfuNo
41zGrso1dGYAAR+QyGYcZT0DVeRK9phcI0glQFPolrhVXOfzxn4FFqAOTwJW0x3J1N3xPibh1DxU
PbND0ej4ilPk+jcxs9m6jdU3vQSfpKXwWfLfbDzJhxE29hS5k59Bgbr0S7cTYtWNWEycrbIcnQEk
3zf87ajV1Ng3416+iq0BzKbFgNm5ZX2EdYMLtV/yKopHRCO9OPGsl93OTElTKCzEkDEaDyd+FAyn
Ap9+ridap6xm2DgoqEmDu2B3fkVUBVqspYsmcQigUc/QV0N12c8aVPbSsgFXhq8ouDIeTd/iU+Oj
uSU8q4vJqAtRTpv6/eStz/kRHXSuOcLbAcmWICSBMgwHpkIMFrrr6nVwc5UATsVR4b0/C3CNyKJ0
McBrw1PbXWyOAJ6564Bz0yX36jimgivg4SBmg+H0QnyL41sJvylI8PQqxLlRK41lCafGZsYH/CHc
bPMSRFtAa/Wmtbuji6LfmvlxzyafhVurk5yOTpyY16rLAjfXVWHMqOzMStRpDoRSfI+vJL5xjmog
FIaUobCIh527Wu9Ee7RsRuJCMSd2lZfzjtj0/RTZm1gsXsfa+p+OR4MXiY4h7NqeAvTY4pfTTffN
F+3TrmTIlzdhvhZxLa1A1jb1Qhs0ANloEhDIuw07NbQ9Ynw11GnvlEG7c9wL4mc3qEktkA1B4QGE
0RL/iN7nWM4dQv/tQZLCVUNX4znjZS8P5X8qBsZVTIkkokSfYay7gGRjkF5v4FMEt7NzxZTz25Eu
Hn5yF1YLY0knS3bJtUH0mKXUXA5GSaJqgTLGZF2gSDjj6CbmhyyMN1JZC+kclMBEJ3P4KeGpYkxv
vPxT+bcI9Yg+RJNilGmpEkOg+kFRAXtfUZYeyG/7xO5PDsIRutBDdzf0ZH6lwAiDHrmoRxC7lhkM
Uddi+y9RJ/Jp0/wu/6hxueA+gHUWYLt0r5CZihEfq6OPZrw7gbRUZ4Rtk2j5ptDZ9nJt6dFmlrA9
oK9uWkAJMNzpawSXAoiqG8JdtSjM0Ly+3TUULbUKIMesodbH4sU9OSGsgSxaif/CKfI6zYo8R0WR
MgPZO9GB1V2MT4XMstyFOH2pOy7bKooAl/xk1KfDKyEEZxY+bNV0ftOf3hPAMrX566YaXPHvvFaV
DXcFpt2/yQJJw5pnLzaQ8q6zRpKF6sNoF4BlU03LmptmvvSzvdPr8ktPVgDlth/cuACG6whgDVeG
7nUf8MO9EvwPzyPLTOtV5uXu8S/zgX7tLfxvIOW9+1hUojKezqPg7ZPoOx1FPAKuIAUdn/p3/OIH
PeJO8ZAfLjHEHoKkI5Q9cxCQ+7vsu0V1BMkX15zK1OdR9owPiux7VIahqhUfJ0flsoYoRqVmy00U
RlRbMqax/SoZ/AWtcAEudD9jt6svxW+o+rI+5nrOQgVADjpBtJ15DF6Zq5luoq43G9p6Xz741dHx
xw2l0zY6fLgg8ip0Msj82AqR7StODtZRcnSPLX31y2Cus4ygHjBy8C50yXHE8kyDpq13EqBAmddr
CJ9e0Q9ZbVsdeJqTyAKKhr+88NsPicr9U5xtGeYRGgJ4pfSSUtU92A2CRFHZemIFQ1MbBvdAPDJs
GQxw879y8Gan9hRy//YvHfoZM7fEUgLWg6b4WmvroRsN3VH+gkNtaaKE4OOQq2Zc4qgLYmF7bHZc
qpLw+MrFZ7k7ekhppVHIs54ZGs4a+QUdBIdAF2VxdZlq77w4D1Vnx0jQypMbgDHnGrc200rpTC+r
2cbpphuSVKVm5O9AEnFsa386u6IHHk6r0rAWXS/K9XF2XIe4ta0bVZSB7r8H6L2J49BMuvYyg2dN
slFKrqstgVvsE5IEctd4GGtGuTL7nzNHQoiL9mCNjYEvt6Pvdf2jP6JoYB2/ioPIRFP43bh0y+jp
rnvBfVWQ103208K35Rf+51FSdJwtIGv/S8DHK43OmB9hI6UWXmInAd9F+lb98WXptQbba6UZavqU
Ha6h1010n2gfHut7gLjk2CVoFHTQALnJywTtUkxma35nO+CQ05jXMxrfn3dHOGdYpAszB2qGqXvj
uWDgbnmsVmQx1+VPfOZBq9c162PYtOstpYVbmH3Ea5iTa6DqrqVmx5C73YjSQpe0aCL8qrkYgoij
tMA+V8/lqA/4vEU5W3U33B8yLNCbwgz1qh0jS18RCgHs2/9TX+jlpFdqt/ZoUvwX8us4c5BSI9l7
s0l21s2djOa1K7ZxqTS8FCGGyH7vsWn7Wyr70UD5frHd5EP+eA5mYiS03r8LqHL7SDKAOJazjXjt
2UidYl9f5nfUNXhR+eHPWn7vOrgLUj+msVTwb7etJ0w0ydIGB284CYofJIwDw2e60XFyGWnTkJIK
KiU4R18Xj4MPveHmNSbBi6AEwNAR7CZXhAyyJ5e+lsT8ZjWgmlHXkfY/Pfb6zAklbWAQ4SHqWpo8
nsYty+JejgaGwhXBXoGeyM7M9vNqORI6ouSkxn+tPoklbM1JseRPIZFfnuDN5Af6EjMfbx2GysTp
gQH7fro+cLPmJTopXAh9ZHpVktg6uhG+w+XqJoexyqKfkXIOHUIxWwmNNKYInPr2/Jnhc+1kPsMh
H9f3bxWOLtkbTxBxjCZFRYAvA27gAshl7y08pDylCqjtDxsr8RNOuBQv/DES5Y2t52csEkhQWLf0
dQZmyWd2u8My0x7IbVPD8/Dynr5QidvZDo+vzstUNZKblATPe/B7LRuw2mhGH6vfoJkapzLuo8Ar
UqLiOX5Ak/p8mgk14Ls2JdSdoMKrTgoJZd47mcmEzW+X4OZXUFNVRv+A75m99QrxeUPb3G6Vasem
3HvaOT3jbSlhb2GZNjQH2NT355nCEV8ocIkf3Issw0V8QWSuZbF+ffbfCZUmKOYAE1jYndEOMHHo
bJ4wDuacKiwiNxZGYJb4sa56WMp1O8kOc/5EeXziPDaDcElfvFGDisePmdG83BfX72/mEqW2oxH5
aeIwfrlXkzFW4DHDefguIq3NQYm9MzAk9QIhgZ1HLjQFamke6W54Hx1Tjf0sJZ8TA71xW4GufHOz
IKOXFZBWc7DbUaACATriAFz2OfYkUUD73KzuwiMhm5LvAHO3q/UFGkIXJm7HW1jY2HbAZ5mDPKKX
Qxh/+t5Z0Uj2nfr7GuJUPzCiFprcJs0ea3BISak4JtuFaVjBt+gsUpEtfZZw7g6wNZdGQzb3V9SY
alqGaP9A3B0SaSG3DWOSq24gBiMM9gbHamLlpVngVIgkc5ipPm5Squm0ykul0mugV69v1pcl38qF
d9Zb/7/9nDJXDe/nqFbdSawnoIGWKlZo97KtAkjbA+e6nKc1JZmb1p+76JE5Gx0RKRg6aA9+2D7E
UpoHqY1KnSLKUx3LX3Q4D54HdwF3rMje3LBWd3V5TTlkPFN6TUBvKyxAKPZXHDOZ8Tq419CgPvdK
XsUj9F0Zptvk5GQC83vJv+ZR7329DfCJMj3mmEhn38mEw5SNjNFZaPFwK8Pn215tOVCaqDtKPf6p
X1Syk9RrTekrjl6DvAZXq085jgxe/kZmeZMPGoCHRzs2dvV8Z5RrncwHUJ5oRY/cyFW17Ck0zTar
S3leah2Pvw53573LJ4ecxP5a3buR0nihORJZuB6Yv54LL2fcMqXbP+SWAkuh1+3yWjdwDmzTvaKm
6l3bENuHoq9mudjhIs/yCsUysWRb6x4NmVDSTX4Hx3mXR9NjYFFFLP7ZLwkxlKDBQ+C7W7Fsr4UL
yiRAGccR/mdG0TF72ldwoOC06fYu7JuZjCexpgSbvYEx6HxZpI5bNCX35IqDFU+CHpFSCL8uf2Wj
cY21YbceFGLgvEdw+fjOo9dJXmS6KFp32t0JOr9fT4NE9kOWM3Zo5WPompPhgp8F7pMC2dmTzAUm
kvd5M4JC6PH/ZG5Nj6AfXs1T5HbbpSs4CVB+0dOiDEfunWq6Y7/ZIwR+YVgqQjgtrIYmUPNeMuIv
BZ/V2Ml9rF7dDqK5rTNAopzvH1wUNXSLpo40wCBuKVUElCQA/D2bV+O5yf6bYCyhQyfdda5uxpnd
qlo4gQrsD/m+koxbFHoDFCJrnSGEQH3z3muxxFmN3lHUYA3KsjKeeYzJjz0WBDNUq8yZ2zzJnZ6I
jNNREvYJxCNIF93XFlLq0PsiLPRFjjyOi6Vzlfl6G0Ypau95wnw0eDaarOEVEHuQSKCpioEkbopa
/WB+3sXci43/mRy/9WiHeJzbUQbJ2Z0aRYdjeOq18j8FC7c6S/rv/5NkEYKE48bw9nT4aQ4w5rjf
tfXmR7TgVPt834QIAcaQ7lISHG6tOt3WdEV7AJiFPtD4Yn0ufI8+jx2wJC3ALj7kJ01ZNbP1c2aU
JehgISNWQ6Q61Y/VFCLqT/y56rcZ94ZYJMr06fg7wlHj7M7U5dsiLjwNLTHKgi5SgUXw3BXOVciX
IV2cdinDcDebOesg7jkVZhHb+Rr94m1kR9qWVU5vYSqc6qBrBV4pcbJk8nk1vJEQPFH8gLxn4efF
tNbaZ3lRpcrsUcXsXPGPLs6gXOgphm5bPfqmCNzmDswN21rEc4WvwJquZiHHS2U5omh1h/BfSvYZ
mLkdIfega9EWN6nPhoKka9pW10eoRFD2Nit5Y71n0SG5SQTJYgR0aLW2RCW+OM6TmcEC8UCGegzn
zvoIr0zqUfwv/URKjo3HcDtW7zI0BBH0QnjUUiZv4jzwAjJlEfpLn55pWCoowD90Gt1WR/JAoZp2
OueHxR8Q6AcQTrS65Kv7bLbM+8/VqnhBXXN6Zfk/+1FEORHAvIt2Ihb2cf3cc4RpXl3jnsCBRAyj
xxpp1Rha5ALYi20acyJ4wRJDRzPqX+jN8WJGxF+Y/vxtYw4r0hCATZYYzNVOPqNW7Pm3XeHmqqkj
26IUC8YC4UEu5UhhmpA25egfoI5//K3Svx7EJRUw3KXCWSJybXXJhsjER4AOn1lLILIKPc4gQ4va
j0nunqZD8Yy44cOEPa9vyD0w9LJ3/RlX2hFNCDPHtrwatXrl6D5L4hX9dtewl/rQDhrfGbWDOMgt
TpydKi4ujsonZ3cTkzeqybZ0EEYEhC0xjMXjnCOaUIWHmwuDjmXx2uadzwycp80hFJ59D+EylZtW
kWDKkhQ3LiAvNgLRU/+H8e/Avuj9iIrC2psiUgoBMYd3l6sCQuwppR3HTSR8pFeNPwT2U9lQIOws
Gz9PvOYg2A36wUAveP6MmRTyo7zyeiQ8jGkCnZGB+Ibw0DglnAZ+n0eNsk9ARi+2zTkKT20GMooQ
mcv8lTM7rQo3Hb/nDq8zPqHko8BymcH4b1ZoyYEhhuaZvGsgUg5NVK7fT5HXTLmEKX5XI325lLY/
g1hoC0mK/XS5ipegoegWMuaU8fAPslLZonoIDHNX2V7dIqozRR8NhA57ooxxsXyZYm994cxvnQi0
n0V+SCloWflv9NBs/ILv/HkwCzy6tEFJ1J7nDp2UqPMwx6UId18c9OFkD/davlXvK7/iP6rmHda7
7vsJ73Hsw3QuSPIC9ofaDpc9ao5EdXx0hrZCquMM4s4vhT4xgPMipr7w+pPltl5aq0vR59XRRC3q
8Y8XfIqf0a5VnRf0YCCi05IbmW7RepSlRV3iMyNHHx2vJogqnuhm6jRzP9BhO/25QNhSg1fnVukP
7wO/MqWByXTv/SAt9L2VZTKDFxX2SXM7e2D2p8/GaslEEIrVCE81WCm9z1WmITWv5lHSLiVS2qIt
HLRk7O4IDinLAPs/VekgMCVhqb5BNlgykjyHX5Qn3bczMvVZ9+8ktatyy9pttLEKk7Q+PnnYHeYm
fvX//OG3/bJRRrKysLBWNSY8AUSlCb+T2H90H9y6RZdr0jEJ9/v/qx5vNYH1ceQC3tCfOEJpWr2w
X8Ef9QoFdBdUzorYgsn4Bpw3hX9kIdSTS//JtfWEFekLz7vo/r4nEz1eHu1AWekunQH1xFyecPhq
UoNovhmCcSMkMBdmM6+KEvZUwGH/hY8z5NfuoNneyKAOplrq2f01JPqkogU63Fdz+X0xqIs+dJE2
U6T+YmfrSL2YN9IUQzyGCcjTnX9eWyGWUeqoPMs5Wds8BmfpbYn2898nroj39M3phx1DSjjoi50J
R4XlXxmQ1ivnAb9oFWPJfOTvsRtcM0uec9iixljL6bWy32XJihzckRb18kF67aO//72QwHRsA9nU
8EixcyGzJAjIYlA3Sg+qIeGZMpNMRZiUZ6hGUzgqA4RdCt/qogtBT2K+IzOgUEIwAnyb/y1fVsSf
8HQV5Wpa7/fDMO3mQPIiykU9RE6lj4+I1Tpsw3126TVa7up3F6/5Q3q7TKpMdUFdcT/RQG0ib0Eo
0cjKbCkdrH2eP6/a/J2tkQy2bOnQEteUC9sq9pHL15gCh5VvFblu62rPoTeBt1XrkvejigcOqioJ
bjyJIdNXt5BY2P40pDV/zrTDygclrraw6lxW+piv254L/QibkitD9PWdoSYggy7Pu0J3Mu8+LAr4
6WeiU5amz4QgHmX4WNhGlnOYOPUX+ArbTiioo8tg0/6cWB+3NW05wPdo/esjXYMfHVlvM619UEAO
8yQNhMl8zSYbaEmbwI3OjReBtqhboW6t2zsdqtMEqpAikAZJCp/yGgKX5NA0FYoADTHBFHpaSqX9
nEH1nVHFTGmYTQ6mssG9vSpjNT49cMyOC4iucaq31naBwMeUCZzeTh8kS8M851yz6/5k5tmP0/bT
O6RQrb40JpEdMfxOwnxFUW5G7pcPzje4me6Tb4QGo793smi2Uod11ABHst0bhV9qJ0Tw1fp9rIEB
5wlm06kZI2bapxLC+ya3HKQTW1DzRGNGQQFmiyFIkUj6ZqlB0pAZ6d46U50LBuB9/ndKkikffrkU
Whq5SkNcChJu+5YXwraCX8IYYRk9ZOO46vKE3xNl+YEx2DbJep8tUBlRsDrZdfXXaQCxJKHlw2Ai
P2pLdmtMthQi5sMRR2dOOabislqObRXxO/j1RfQnJ2iLwvTNDCTPx3CMeOkVV1gYW/BDcryEMEAb
A3vcg3KiwpChJrUO2XwQVVONI6aecVsuxmmd0dvr8EJjQ03NIDkx8uN9uK95HdQ/WA0iNayNwNq3
KDWGOLzytpPhpuw3MtiK4vKtREySSFVktij6QZjbkxYkrP262KnFDQ2cY6Ieo7fMPIVLHq274tCF
XuYAafRtpW8uvoJ1UkijQ1reBjcVpzxLL0rvx7YcMyTx6DI11aV2UgtAwnQ6zcLfgPNgfAvz+drS
J75TTzdaLmDntxp/lYqYaQOn98HhqcIcvTlT4F+Zo2xEuacUB6qyQpLQVQWzyOtB+7sfYog+Ejeh
9kScvmEBY+MUa5uqXxVojqdXvx68+AkW+EcVUJ5gm23nUc5PUaOz0QbODMS9DRVrR4dZYI5SQEaR
iP9PBTXW0LpARnRk1kwxIpqUm+hvyeCnf70LUbqny/FhiTazcKZU4RSKXtfnIiaT1GxTCGyW60wj
43HW+zGZJ+p8dOb/BuxR80Aktdyl4ITdm2j5yzj81Ubg7oXVFlK/F+14sih200V+9nq4YbEzSOBk
i1/wSGf7ta/X4fijX+wH6yAlBY5qFApmy/TdT2EXbzpm3071J1KWB2WFtwt806+vovaZWuCzEOL6
9t6nHaLmf89WnGE+qghE6wwdjpbYougzg8YZl2zKgQt/bQfir2LKVALd36A+lYBcW6YopqP+XY2Y
1fQAZGwJ9BURrKhM4gJQluBUgQrkO8b9ReGfcivwXYxDL98f1ll50MAkHJL2bZH+hhSvosPS+pID
mwYFhWTmp/bXwRWD/kLU1TXH21IDDxlR1+1x0AdeaMNhFvK0xOcxkVxvt84VAsuvCvlsPtI4O0KS
VZOffXe3/q2JdhqUCBzoeCXpA5rn8wbzm+t/aZJVaQTMnjm0RjqNuD8WqxIW/g92SXz8YGuK+RRb
jQuEdOo/8rb4Q6NJcVChkBNbEHtfkePv1ldhIsO/hbDmyF7p1wHM+T8udE07T9ch9I5GIsKrQiWw
sUdDOOAzVP3KXz01SzalXUOTcXISuEfN2Sx7iLbyXng5fcm19weM1lF6Mys4sFZqmN+/YFgnCyXZ
hCwQhq3Kz32zlOvrmuIWyB2Er78UT4JYf+XwWwXJ8iNLfVPvMBz3rPe+rOzHho6fqYOpHb7cLX57
vIKJVvifZ7UhLtLhS+fhSWylaTgHzwwCIo1xW9SnV8a5oe7NYc4M8aqRLeiJKEEBaJlwaXyq+JwE
Jb2sLHSInsXQhbX/JnZ1D6j+T4y1bJ3DxDwQ3bu/VPg9kkcMKc184zwjfRj4KZdI5wBvW4wl9JKl
sE3LjXoEV95C54OC3ZuZ7M7zxsIhnk30IKbq48Zer80eMXOWv4Src7HvQPzLJjon4eYsiPtAa2Ca
GuF2f0WtWyME6iWGTdVN/eCSiw55PmZ6PqAY2+0s3m4bqOiSZfbEtRk+I57xAWp+FuQQeslFXg3k
aPdKGeNE6apj9sB4xkI25EaElU2HR1cDvfacTrofUaWX0B5yz0liffvkF6kCoWPeTyfCy8IUNblZ
b+j0gQJtDEMYimXiKKzqJujp6TGC58dvC2d+hC9IIMgbbrCAlBgODRnEEWrvOEfZ0NNgpg6BsvVq
0FBrtyzTsJW5BHmXT9HZtkEuGpTXXumXzZrIGf7ngaGOg+bALEHwzpg+TpBUR+h54fC64z/UR1yx
jFYsuYm3lcfJeqcQwI+/5EId0W6DrbLcOQC2AiKgXwBt36FxbrbTG1qcmzhyj0Q8CDvSX5WXDIpq
DchqSv8mF1R6dONBgqNYAa2mmvyJqrREihp/8PyCMiSk5ehfCpcrz7/gZ8AW0+VG1Q/ct0mRlHfb
TsMoUGYO/4JQPPbIf2QSr+yX7adIYkQQMaqKn6Gd9jW0peDKqKFG4GsK1ZorIhk1AH6Np2scLgvz
gvTrBM/I2DW3wweWhhDbp5YDPp2EA9bXwT8iyo3ftKcUH7plqGVyyZsFaPftkP4DDfBqWUZiKCoo
LsA662uBFga26Ft9n7kkdAbs6MC0t0EQMv98rpX/EZRB0HVvdmb+XnBc7Owae2lNp+XZ7wJQXchX
yAfHatg3toH5Y5KtGKRo9JBhFNOSJPKTiIs4Vio26yO0s+iVOrdtqHuW1Fxa4AMnsZwmdgpNjsTi
RRkAubVSieVp6/w3xxPDITQSXviTAkC05fcbQBdMFEYWC1Vb2R90VpMH/RUM5omPqi+KElQbZ/gi
6peH0frZZ/jK4Vvo4CgbfoAFAkA4TCcAGT8yp4T4qjkrv0Q1/YjKQSvBlmoL7rpQhCtTAs8Z2B6Q
Q1Jxtpgj2XHTGjI5R+/DeYKfDp9SJZWbBH/eRg5Dprreuoq5A9Xg9fGf8y4vJnfdugCsEHNgytNR
U/QgmVBf9szW85tOWGwL2wOSEvuL/hNIccK8SRaP9BLUWI7QCHWWzVZZjYAbVeFGU98RhcQRlZFV
uBveIJrT9Qtlhhg1AKR8nvhiTbOo4S6x8cEk33bRaSKXcm+GYt1s9RItf3+iRcEqxfOorBULBKiD
ExelFXultrrMcP+EwG8w2oOzmkM1ve3TJWeaa65ZrO4KtNrARx1C0w4bd4lGLwASYvYxE/ybFOMN
Mws9LC4iTb2teIdqjSNQIkM56c1vXq2jlcZ6NfkuAji3MxQD5QU+akTeAyzfXcIRaSROdQwi1NyY
LnF8iUNJ8qIlq1kik4VMtpyJuVcOgPhUE6cfHjd3690Lsl4qsU5J9vZRcvFX1jWWZUI5e3AxzMMA
vg76zuBCH59wPZ8O2eDw3kmrDjlyvJIl6JxjZ465QFjiNHkqpEUGEo5FY46gkxdi17cBiar9WKEw
qRKULKD7mGA4J24FnMiV4iyGs0wkStk8l8CMU/f6xObY6ljxAYPUmvjbvj1vaMO8cu1tUIk6oQHG
RFZh+BmprACv6Q49dSsxAvFihPsS+HTDC6e+PI9iWfM3Q20iY+d83ovr3N4tIeZ6BFCmntfM1u7u
ehyNOIAsATAG86PDDUqnOQKo2yLkFz1RzZ7nRsmbJQ4sOvHyhu0LfjplpEWKd9IvUQ4FInkoxJCj
oRONevrwKDgAp7qcuDOLuhc4rTwWN56YltpTA8Y3nbEuRU4xSgJspS3qngosptBHG60sHjVP8QOs
xvZSQINHQE4I3q97rbTsRotsM3pX1IEnuIYU2EuNVwSnlp2vnPsYzEVOyVA5pzuPGV2AsNB3dL7c
qRKbKf45JZZBoFnidqg1nqwhlae2kdQA1BrTTdgJWjiqZ6MK88hjxRcFJYLzcqAT0QSq0WMzI/Iq
FCEMcd++U5FNbBQN73QvgFOKLLEy3aJ6zmFGUUYgSq7LuwBeGW2MjijKMNmaPuYlUOa88qlKfRQM
dF88RCm7dHdVRqv6lj46uwXoUWhq/x2fo9Wci1w4XFMmG2BridmpWdeahhvXdKr1ym8stMF2/EKM
1NCYHPoo1D4oZFA4pxDYg+d5pbbY5YcYnfBu8j/wcdFWspw/kQ1fGzZoqpv9Laxxc50lMtEmI60B
3fq0RkRzbaup02eflPc0WPO1IMIM31sM1D1WQTyqoElTRuap/oiRjL7heLAKv5XJ2ORB+byQ8tAL
419CwVqfoYR6G3cQvt3J7dKaY6nCofJXEWQFZBEz9oES8F4+cImX6+EcCazc8AA+4vtDlxk9EYg3
61Yu7a/UWJJDMC1gnZL+VkYIOY06nCg2MlYCyM6MAYk8TAL0jy16oFPv3Tecp8u8S7MESQ1nJ1+d
Wwz8d7EIDyG4Ibx5zmxpKCBRPYGr+cTx6Ic63UHnkXEJkxAVxu7FUp2OuJHegwn6lbI9TsUhP5Lk
83xINhPWpAkuUsWCjz8OMxOAhJIJALJBQ5iG3WzOSWkJfwFXZFtzfMkipB65bdHPqbz+8Bc0OHZo
URXRSRVy+EQxCMHp2dndzj/6s62NYOzHMJ3m0j4bjlPdZMlqOMyzXI0P+0hA/MeS5EQ/HdkaNSQD
1GzXSMguA6GSaAFDIxOKijKMa6/QD2JxqinuRSpXO9xrRFO4csizJDfcojxgzzrY2n9MZvOJMk5L
Xj4fgn8Sb4GUjSFKmn7ly5oTqo9du1F0ZHPBaxrxJBJ42Ecu6O74WK/gB0E/mrZC1qg1K+oYvWyt
HSClhGI5zRktGHFPpPlxXxIItHwSxawpsWsJOzcjPMAxFCVUdeEnYXPNeu/w6He3mLiJYc0TL0cl
Cpnr0bIeCWzsoq78dKL7TDySpp52v5emnBw8XuZw8QZZTr8OZcrPsLjGjVjwUL/6wZuoZqMUtdid
Brle4esfp59+tZ4u5bauMzsIhVQZUSFd95mcN98I8Xjt4vi8zUh5qol3OIxtfFIbyfkCvIfgADQH
CrYgXhUcUp4dE/ZOfiK9W5mCQB4goCye0O2+oAamGSRn/L6B/qioKa6N6fcmf0PiGDraEvp8GAyB
Duoa9bjTOZmTwTBpqCh+QrVMzvqhQyCieMaPAHHUZVrXSvzOK9IsZ8RgCBICZYy3L/PbM5Lp84C0
f0D5m9a8euOIeNKznSXipG1K6zSrMAHPkS0ERMJIPI5VNdJGGvefKvltlk8vj9XiL4JgMMkzLDP7
VFiqXN9qvFnknaXPapgfJPoT2YODYwycnAy7yo89+vKvW1z76RICwozhyS4URksmPAKEGs7T0dYc
YPqxniHqkpzDiMRjfDibF8A2v051ZiHPEy+pI49knw6aWnz5F8OXK2hdfQOA4zcoV54Bc3L40G+9
XDMFKCcgSKeBFdxZUsS/cpR3hR2sGu+eWY07meUCECr4XMKWJ6Iu5drAOF0EsD4Px0pp0zvdi4kB
9sQTqcCtPBAa3nO84OFWMFAzR21rP1dmCO1N+wu9DCVfuaHDQD2Bbkl2i8bqVdYJ0H3JCHsJe4SC
susj7rYMAQsVsgBIC2lnQ8NIrwwPd3XLSqnp6sKD5sT4z0uxMW6Tadjr6/E1B5xf/8JJ4R9719nI
obYyrS1KgwgHurCd2cNSGo/AQx61kz2mNFWEtlEVEcczdkwIZDsMMj0YfB5iuLrjYTg51IUT7Mxs
TafhDth5bEgx8VEXURKQjFe2EOWVOHO88BIIRqRcyip2IWsmbz8VW6G2ygbr+0HUvhUcndjfSH9z
OqV6dcFctoweD0ECR2VekF1pvSyp6zMNEz1kah2xnCFShuRioMyzhZxGMnS39kkGegAtHMaTOygr
0StOA6fBZxfSkBv56xZW9IWerV6uw+6nHIce2xpo5WqyRUTaVP2Smeua9AWx3PI3FRb+ykV6Vql5
VFOmuGb8mbgr9nflxvvqhje2wYTJurcH1490JGn0ZgkYbWuUyPeTyrY/E+lpvFIFJ7FvZgG//JPd
DxCEeim0tEoJtZL6KjRnm9Enhhcz9/uhQE1S2MpidUfoLJjQb2vaLow5qOL46AaNVezbRjmJ+0q3
1h6u0ODq+v/LXlcz8LYOTl3jiG1xiKVo16FBui06V9FAp8WeSDSUWmkPDhbUWfwInlgP0O9nEmx4
8M58lU5SFifL+sOatOAn8z7FaLvQ6aZ59G7M0f5ShTw+ZOpb6gFFMToXwxQ2Xx+r9lHk0nRMPTkv
vDeWRiuK6NCNUd8Qw5YRHDugT21tmvLaMRl4KRGMcNHOlgTGGp4hYfrYUSj3FKdDxsT5Y5J4F7Op
xPpNd3zOLGeBCn1YyVAnDKVSduGRlSVn8aCMQWctzakTqlXD2gND2ytcN338ki8Q+pL1zumn6f9/
Itz6Qqap3p7gPMX5HEDj6Rx7LjW4bx36v1RXG8m9coxxSiSJUwa+qLEJVR2Sod/QoSMKY1flU06S
/Ao6kXN6xjAMUI6KE6fATsRtRkKfNnlPx0mPoFXZuaZJ0SNb3eQ4Izc2YWsehqbMh1GhL8WTNfNC
YrcPFzligs0fP9uKN+Q7a8B/7DXmvOD3XU2JW0w9QsfzJyS5+CsqeHTI6gtRrk/9p8snCqI4ZkmY
7eLgByAH4xGQtTIb0fjsM0ldK3bicySIN6NEwIXAQN06W8LwoHmcm0N0yC5pDEEVY5VL/bNGw2n3
XXC7fF2HZLv3ozJJ8SGjfmzUHWaz9Hm0nNC8LrlLW8KvJ/S+ISFTdmh8TCLH3dWBugUU9bIFLF7c
7F/2TO5h9XYIs3sAPzevcYngO/WRVP0qzCH+AxiTh7TSDc4ABLp7ZTtbDU1xj6mxJKm8ZMuZVAIE
vEp6G4dvoMoDvQgxSbt/SKoLQDTGMDEG4lG2ZlM070I2Qcq4MIHKWxmQ1sMz9dNRo4r0IoqUvogw
qdbb/FqxWyXamD2w9DC4r4eUK0erNveMbFH8OhZVdRhcXrXDIZLrk+MMfbjSP6RySmmwh4eyjSxu
B1/FFOPQz53hTf+0PUdq8xwU2M609nYXkPGsundmrEpJ7Y1/IpvBv19HSnjSRDMytfg0yxbMDIdG
IimO8ANKa4LEAEc8hV3072bYDJpJVtvLT+ASZpGDXwaWC7hs8wBS4eh90JOtBW4irXiaVvyh+qYs
fhv+WwmKJPk47XsHECQFLM+Gr/XquALu9LWrZcGZAcXpi7tl8bLhQsuObmpKK8yZQg5ImxtgEo+J
ntD4in4Al4agmYD8OH6Axze+YrJAPamceATc5GaKB1Fk/H9oF8LSIt4Q9F+c5QW4oi6I6jatrnND
TZhHpoQoAR9iGBbDRwLWNtQANOBeSBL6O72ZaEwcGmowTKHehU6tk2nMjtBdXECak+px6WH7MMid
9RnHUKvrYlwXsIl/QDZ4QpZ3EzBFaJNolmgvnVS55B6XTR7SdI3UykQUFH9w6JtwV6oFb4b3UcmQ
6v1OGtzw7LzB5Sy1geq2IafODX6zWTdatSK0XMcJ0LsW1uW0G73JB4KmQ/Q6tCrQEtNY/OzUBfmC
Kq/HbaXiH7Qv+ng5oexeTbGGYH+QxLoIZWr65Tpy57/PIidmO0AjlTSC2Tbe9MfxxY0mdH0/zGNv
tF+AE9XpXymZfaafoCk0AXyvwDsCo/amMV5AfzdQ9YZ8u7PWkPkl560u/kEfzOkOzeS5em21cHVV
5hIPB7jTd7yGOBjMPmAKo5YAGwZ3FgcFDy1O1wZ3rBA5pCFv/tsU4xSdj+3pAbWDGma1IEaZGsXx
TyimYGhq8utOjMYv2rX4UzGVRY/+SvhcearDGQZA7M+r+CCa6iKa0543Ule9L2vRE65Y4IRCsNh8
CZ8YYdGvNXaANGBhWaIkqkW7LO/3NAnz7BGVOXxOHtPAy8KRGE8PeDpYemhA/+hdSJXLKyDCFz6q
FZ98WJTaMbqCe1/LV19FOlAb0U2GClEY8i0gFlApCVHe2cENkYPu5NZjGYv1yZys6CDuuMDbBF4B
YXtiwWUKq31YfGa5KJS5+9hoiDVK8mIVyuEU8M91wa+RqjIeFeXRrkO8NW3VRSVjBiG7dbUFo1Er
VNf7z7kcJ0aHHYCTtUuCIL/Iy6eq8d0cJtIrCaGoFRbmpSuLy52Np3bxMhIiQKcQKCjGZN7Ynbc4
YE63bGwrx73WaNofu8AUktIEw58n4FIFOe6DAEAZbqR08II7jPOQb3xq58m6X2ad4LzMWSMWQhid
G4E2jStmCaW8pAhOiN/vJU5CFKtU78ObfuWbmcxGs2uQ5jlO+G9ubIkg2OyTUmXFR3/+Pq1NrTKl
bkym0d7HOoA6StRhV6iRcSMT+sst27XHGfmS/gyIiFiqZB+WHqMYOw37I3gcpSBMnze5cq6654xX
FzM+IJWnCR2FbXwnAv2zVN/ZBjk4pUJCo9HKF4TPizcxztdiI2yCLRRC6qiX2YhKYVbyDKK84nx4
FE53Qg862dHMwanAmrLVjjyWxnxjxrvWfNuhENkTGaCB2DpIuaJ1XU6ZsNcEljFnWhsF7dursVBW
cdJLRpE/JPzisdk/4NteFjjifHIPaCH4uKoGlBvq6CHsL17FYmuQR9NJxQM3mSLNI9gQKh6eKCJE
ANw1LQiB0xV1c7IIShzzPm7FlAWRmqFsA3v6CTjtKMo+PiiF7BZQWEh0qa2PiUx+gKt+nPv+1S18
o22Ed+o+ltmW9Ir17/WprsCFokH1qb8TRk0zMcoM2JaIvemsfCdwKeZqaikNCUVcv7EtzwcOxSTN
kpJTalfk4CHsuI8x/EpSZ9baPw/2eLWxKq4ZOM/8umpkm5fuQQ6AjNz0l3Dcc0x7oMi4zTRzhDBv
+RLQ82BNiJvtugie9bfR/jX1l8N7dxkQDDrvFiIb/TW56EV+z6HYuTTnhuYBdbrVyt3MDpbiJRqs
6/uCUCVpO0Gt94gcmMAcg2nFU/V1FUeFOh+Rif8atZGrtDyvSosNpuXrvnAEDEWQyji9ESZUTN2b
SF5VBd7ivk0yFM4UZFSxqK7ID76qbM3x+g7JoLeB6Yp6f6QXA/uQct/Hr3cGKzHzMEJwEIDmAe0d
wPq8ug4dQdCy8hMidnRvl3M/8XgjamPQ5oBzjRa2Kw0ozatCLXm9Wp3Lofx5x/Bi9LDbM+7gKMxj
Po+Kr/9jL1W/Gev4Di009BsJpBN1EhXr5Q1BUheHaYBABsk3oQNe7zCDh+vr35Ap0IfpcmEGfQ/J
4cTbjvVDFVEiK72jHMxwgOm3rcQuUlrJZrHw26mNpd0tq7A8cS4ZrUZLzd10q1sS0CQEf922Jy9I
xUPwTrVw79g+SLamIE+bm91trXcA5+PD2BVKlj0mf1KFlD/wlaXJ0Q6D6SF1ndTgazisRvbwfc27
qRF8bOVSEIGmVkT/16jZfuvpAzcNUzd0shVhVTGl4waWggI4VbiiYV6MeUQNKA2NYVmLb+ySEXBM
9wiaY7dSUwD90YL4JyDtutWZjEUBUWvCvjXAXWbjSUPje83A/k9KemB/eDZPxBi33qVfQ4YiO6TU
CEjhYJ3d9XyPzMExR6qOHlKUZddSuUxuGFr7CkCuApDMbIQx4PI67jXrhA4qjx9mWW+Bo3ICm6FB
a/N42b8dvDpuqXbQP9tzubA1LO8+yeCi7sUcEopcci1PIPA/6ImtFOEJIoFZtYvADMF8+tRtKDbY
qDBGi9Te7RQ2Dovp2OvJSAq6bh34d+FJ8ZuciOWIeU/U0N21Tyum23EWgklCXdN9YGKi0OVtHQGG
tWnHivnQFoalvSjKEw+vJCsbwHiSM+PbLanD5QByPXDeH0PCfCa8qYJNMZNzrILYi9A59g2Y6qOY
M9B1MDHCZUwOPOJHeijU18Q31mNreQc69Jk+nMNAkXUh7kFEh0DA/4G5Zb4rr4qsZknN/c8zBo6G
V5DE55LwLrYwplXdCdoBxZZiABXLxUADNqmWhK1vL1rhRh+wyqcRZjXQNlMaTclkY7Bq6ECo9Lkv
wh8B4cMKntiuxhodsSZ3WsqiI1WGA29Q3QiJ6IhrzqDWGXD0VRwxhkmQi6Z/9qNaEPdE0kC/FPx5
FJaMauW3Kl1OYTKrjuB09XquFzXIEoJ6GAjgTIG4pNE+VsnPGMGbzgE1HXwrXTVRgZ9nvKr8h2pj
FIxbwAsd1BD16Gv7aK1XUKpTPThSrnMSfR7Q32lBUqWhcLxq7nBuBZOhQzLYNBB+uEfdLkPhf/Qe
ruiRZhsWttqDARW+YqQ207WjATLjyR2/5d3Wd7YKbVklEmp2POa0Yie9+6pdjb7bWnPj4iFZJfIO
dYnreDC0jFIJ+2qM2vk73t7KXsHXOMcu6CohkbG4/wYR0EwipUgGOUahFuD3dhNgE/5NgeuSESA2
gRF42cENOu7O/DGnzM+Q5m7K254XVkRN+35b0cZU07XkK2nNNCZPR7cLb0ewOc5lwE7a4BMUBx2P
ZGyVMCJgEU7SjNobylTrB8hymdoWXfvItxVC7Qj7UABURzlMi8uKpg9V/oUjPSAtnSKDfIuNEzhv
mEEl5gT/jsxyR/IoZ/M9NI3gqFgvSBa1UZluIblOnAmtibg1m1/jGZVKsk4PrNxzlFYaYaSLirET
hIw02ey5N5Bhf2U8Pae9ZPc4w1x8buR0Tc8LjAPEV4/cXgV49D4cnUFSvaJtOnenreVPfQyiA+uW
nLirBbPkGQo+ScvpmhJY1gLNFIr8J6PZfix24ppsloPX5iwq1qlbZC3rQB7ZPJP4flo89M7aV+/w
Lbfy8dgP53DOPsnc0W2Rqx2qKm72C0/AQYkHIvy3ZzUkxYueJFRyBUltG98KlvUj/BDtuyMDivE9
q2u+6U00b/x2icmZyamO4pauiiBL6jUOiSdmUq+50vxnuSftKf7m/9UxTiiGCX9b2erY3wUTTpyv
hpMzuZeKwdLkqqasNcONB7jHpMWxCP22TCeGH9BB/Agrc4WmjnUKfKahkFKhovq4qtL/IundhT4m
T58SHqJfOn1elCc5Rd4Mw6AgWAvBoRNvAHNB7ahR5STjyxha1tdj0YeTA7ULipmXutC2KIq/sNbj
kANBUHdYb8ae4pqIR+hbo8+3wlOl/N+3qCJXGUXe6T0AYcWZp13Or/V7DzQhI1ROhE1gTkGhJvp4
G4CuBPglBH963shexB6Pb5GkDHGENCr79a+seQmtRfxtgHUn+EpnGtqT9HqlWSKv64A7GhVTMIoL
uTjOYHeUOeP95u1aaxbJWs1MWcmPAawYU/ispOOPd1G+04gaYJiDVquAYkSvNUYU3KVUe6kPRvsy
YNxr+hO3JjNxaz/Vs5ncwXSX7TSQ9wf5ldeU7G1kZZHJQppTHPaX1Vj9nVEU/6ors6PIuf10pZpL
FzRie1NjB01mKWO6L2JxOBj2f/5Dwg4VKEeqA+K8IA13RZacT5C+zAXBqTukF//EiMIi094orTFY
x/AfYvfGhapBmI7IheBdrlpwsNHtl4XVV0NX6yitp3p6UeDHQPpTRgnB7qLORpUnTZo+ZoQp1BLi
H/RTgzNHmYPfvshvFedLMMHCI6Wy7mesfrSZWI+YwyCNHth0Z6Oudw9Rlx3WcOCXcXPgm1kriOht
Rl9JVDF1h3RcdRCuwBtvLpMmvy8HmtVcuqV5/MXNXV5xoKS6kZntY4jtCgxVQC3Fkey5sPIO/qCY
CukKUtQltiRowttOa1NrJRJGR1axGs8TyySSaFvUexkxp1fNIOyPQFkZZO9gEQPBraWCQM7vNL64
cd7xhCAQl31PJD/djAwJLOu6aSgj6tO3j1+oCsO+H2LBbUOfeJjo1fAHJCxxaHkvQnXQ5O4V6AKZ
pBno1XZ7Bs93MXa6lKx9sS6zZtAeG3gKno5xiIRdrEE9Oo8u7MTbBtVu8YHzjEI7Sd/48LqbgplC
m3FL5FNy05fsNtTLjUCrHQ6BahZ9Kf6ozx/pZaPIw3O08W07tH/4c6kwznXn1ONnBCZKnzMTidJ6
2CTHUDFfB06D2ZlOsTG3whKGDvurlAlkdERmWwuKd/0WvBOEFQ8wmSU2bhecHlmB7YcP9lo+rD3R
n7190HJ1x8TV91qHxHhNrss6422s7NqNS/nFMk1sSstl8l0RaJVc+2NJvc/QkZpspOIfI9C+DZKi
ETq5Ol8fMVfPiie2yXCbTpYKF+vbgw3w+Gbny9Duu9VkSEgtWFJcO6SkmhaiDUkkGR7W/q4LYlDJ
+CRGBlq2BBHPtVuRHJ32Cqde4zzjlwUaZ2qPxlolJ/0vUbFuDaDoLLJDae8WM4MLj1C76Vs4cDgW
Zi9ES+tSjB/4X9RbbomeluSnnsRez1okUlxTMJresxRyzakkwxkyG4Y5Ao7G1SOB8uDfWxwBVYu4
ljuIqkdCVh9Iq0RHr31nvA/tCopLVC0yHApmnDm1xuPGimDBIJTLHJ4WfL3ooaWBU9GvtmKIeLFx
Ozke7/NezMHa98wwPXrBRfY7JdP04s08yHNA167yu30H68N7tFXbaZvWNz7EzC0oX0sUw4Hshjvc
gyujY2acDvrb1L41SfIy1FLHUIxBDkhv+8rmqdIGcQj0nrHlT+N2pyItT2Z2LYqVKjJnCHy24VrC
cyzOMbPvRxiBLeGmnsEfVarlENMSwim8PHZ+m9fGV5WLadrW6QS0GAhz05Dfra29/S75/6+X+tCv
/w4D98IUp8GvGL85fXV0KaQ8HaMbrjmBOvLhTMKHvWBH7SgldsH00BbTjD+u1t7T/TzdQNeKHD0L
3h6KUlpxfZQmlSbFEWF185dubAzAmw7Fhr5BS0c0UFkBj2y7gOurPtPxj6S6DCTGFzXyzjNk+JoU
y/LYGKLsW7DQW3uURlpwFjGHLLKUhxH9OVDuGmGnQTKmejEvcNTaO71rzKGx6L82Ufy7BExcZIjd
KyvOMe0giBcehFCkixaw5TJqpUhra6Gz7MNBQncdpY5wON52FtJht6PNyERZWHDfRqODqMSXxuY0
GDv3tTN3wdFv+mAVBYzkzFZUqK1pkXpX4+bTX0pOuI23389A0ZMiuMaCJLpTnCVEwJnP56/okbzX
1103dX/nyQY7+PdNFlDOERW/nyZqqhVj06EFiynbcJNWlO4WRGYcdbwPDcCUetDPgnBqDNB45cDQ
bX9vEKckObfhqiYr1MVEsA08KwIZUqUdNfko/rhKpsk+/MshmYiV1iIV8HJabpiO8GPGmuroHlrb
224kXxHZeNAZ1m/peI29ntMTLAEtTsvx9TmbteWluDuik8sddex3OrJ5aURed/0RSnRh4BAAa5H0
wq2x5b78v3kNiz2M9a9zDElxpt47ggO5aeaI1y4buudLVt8X/cwJslmIxBov9Q38vnb5ylFU9ZtV
8hp3w1p7eLQaF70BCJcQItK1Qj7sxWNKlAEIpJRRFCyLBwPgNxGyl8eVEfpZfVlzks1kba52LtJB
aP5/rQctXxjWgrkxsFOvnVRN/G+95B0/x8/D0G2xN+ufiF+eriTLdHqfMdu/if7OHSJlIk4rqPzS
1muvqJAXyVFFXV79eG+gtv5aNea6A3lK8hTn3g0yjFMTJWaz0QlfE8tC5L32I+e/21/ct0iLfYff
JpKb0o8S0YMFlE+13l6DPldhZGJD4G+Da1A3XGyIPCw5duKI9ZDRvZSOK+V2w4GYzabqCG7PHM7d
EMlz0ZGZxiBckYx0dy8sHMuWI+A6OH4Vf0xP5zHrkd1HbkE1ovy+BZtzNcoJQoTCXhVh7SdyK5tg
jUZQzuoto7/5oNHBigD1GJ85xPqVPFye5KU44hd8oouSdRpLVYjlSeRTvE3ZH/9sR6rcsyFwzMsJ
cgYTxGSGAYH/UuPSudI78eOZYtRtXXj6D4PFZhS2TdOt60nAW/3wgzqz2wy+Iq7lkBPZjzgoIbZi
ThACTPYF6k1aVFB8MTlsrUKEcY/VGbTgW4EepEEm6osKbrNz1hB7+0StyC0jEhk/EVhFwD+HqVro
IvjU//hrIyaftxRpTQUB1+4/GZ0P0r3o5/SCGuyBAfBryrab3yJxZ9bKrFIJaa00rAi9LZyCKP1T
hW25w9htzEuNzadTdUbuv1zjilaiuhWUH3rZy6Sm/IXKaooiRz+ZyqGcOQAuhjA8mB1zbIod3MnN
dtBcGNG/1dX8oKVp7Sj1rewFcPjigfNwOuzQYbrRYPNUGABHMftqa1hoqy/TyQqxXWu0j+NHx811
nWxMMkGgHr5JLTIoxuZw5qFefr28gLfMfv2a7TTFK4IxCMkdp2pk1V2jePg/5oEffj8ruQSMhynY
VnebdKVlU3unF+efUec94vu9hGiFhIpNGFsqbbV6RCUGpNaGCklx0WStThTcPG5tdbIRtvDcdopQ
ESgijrDvfDYgd2iyjVNG1Bith8w8jmnF1pVXZkSR0lmdaShgz1IJgVWxmi9LvuuD6YZHDuSna0Et
FuAPMUwVzk2XrgT4G7DNelnC4f2bBkdbqIpUPOYb/NUpNo9swi16La1m3OQvoUMeHieV63GyG8/A
qV1Izv/Jaux8HyxNMyDdmoHWnG5ZK8L8FDVRS01Z10XD1078jB8iyY1IIWba8hDO3lv53Xf5SAJP
6DGIQXStfGz7FcocBm/mUPmYBgUGu3wNbrjTzY06+de7JBH2aI0CdxlcUxAVH6C1grQNNkc9rS4p
0z/zUR1kJksKPMjnYnPXCD1B+n8cZydPa8IxhJrk+stzZdVpJPvYAiwDVFd2dnSsG+yadU452UpE
Fu650X627yGvfc2cE8jY9pCg3u4tAquEKllpD+/ScmAVjEsYHCyNzSvHGOzmX4T6Zf7xb0vUrI5e
pNjg2w1c2mTLlWaYsaXnB3dJyFk0xaOz9IEImYy8hgc2V4TOwCgigKcx7pdW19tiIZagmPz1QKXy
bsYYLHi3LakdHW9P6C6dbPrnxnwL82zkQ+awQrBCZGOjKY1uMHztonHD2ItvB4ZPBtCxmdfkpdY4
2i8+joUFgCISaO1h49a3Cwi7OZ+TjkDSsBRcvayDoD1ZyFp1mskF6Wu+3ks/iE+dFgWnFxUqHG+s
eZnoVD42dy/STTvlP6korCVJhloNluY0ZPgDO/OcgBxY6y6jIH2BEHJbbKNmMO7zCElPWrbgY9/e
Nb8cn5R3RdQjW9tVY2uE1yF0jmE0NVMoW2SGvRke0jkp0fINeS5vC/7GIAMbl5H5lxQWWB5WmDqJ
XvE/Tlf37d/6EyKAZMdoR4XJwwVlEZ+qd1CdYccR8nYzK8Kz78dYYSwITa1thAXMltuBOXIS6Oe6
DbbldORyuf5juPKuXQQGhxBr+vvD5iHmU563VmdpKInuK6WnYEu6XtO0+SyCUEChSLel3D2QogzQ
Fc2s7U2z9tiSF8hBu7IjVz/vhfx2I92UfTkTs07A95sSFV5ZUsP7ERIYriyYFNxyafbH68XBfBOa
AQsCMLcQhou5ptVrz0aOnzTSttY+g+WmpfKfEAeAIW/UPJdodFkuII4bvQ0loHgKUOqbUTaancqu
5LtwayTSksNPQdT50QFVNGvrtKY8e3OWFJt74OZWr+iIIAPjAlUbN/hvubHxyXRRN2BjlcojcFSf
7J58nMpeBcPcZ9QizzVc9FM44Ji+JBwWnVaqQIZ8Z4Sk/QSZCQbnZRCm3jevLM0EagXy4B1FoxKO
dWVkQv4/WnpdESQ6OTaO8i9bwp8A5e1/477hPWbyxgdoCm40ZZIRnObglGUTwdsz7E9I5L3ZkPub
rTHp7YTVGd7d1EAdNpd43jfBxuizoHEWH6BoNjMSTZmR9tetTSOh/k3Wxa/5spO6ve7f7bX+Gpi6
wRDFxSaulydzk3E10Khg3mR10kHy00pB6B5lbhmMjwTtn+5B7/1MUzooGzSZ/ySFuT+VmQ9F13js
kZQpjjnIGqId7muYExIe+NyprjlXUG6/Q/PjlKVTGndQDm3H8+YqCLs8XaNltyiZ0A/J/X3WAzeM
Bt9YhI1ilHuqq5YkC8FjC03Qsuo0I9Rsg1pO5pWMLba7yGValdQ+0G+8OXXwGNprXMbAa88wpcbv
J0ILDa9Z/I4XhivrJspMdFd1rrZvSJeEVrlauhfnMf2hOyJNww+iCatbFOavctshS6tl+l4m1uPA
F07JFM3DC5kRqWyRViYLdByrOs+FaC8vAUGO8JVkyguM4+C4SmEDNxLCDcbh6W0JvcFZvzy+VH2t
cidi9T3ybLdXlfOJqNbbsAA2XtwjO9Vwt6OvsQw2MxDKsTqUclSZR5yRFSm2Vl+TJGeS5OSscypf
ZJUp5n67M746/tJLy+6it9ng89ck35jhBJp4YpSMaHsFsP53ORrSISxmFziBQJIAF8xMmySDVc3W
p06Db0Orh3Z53cgzgnZuFZArZPhV1suhPlQ6nkPj4yLY07z3o34p1vO1rBBoj1T5wm/HgmFkWpif
2qhkk1+SWjxPsjs89rEpWfATL4L2kQ/7rMGa0hnmJeq0OqmvLprj/3PcMMV5Z3VWQ2S2SCeayfK2
MUtFOyVLvcGCHo/pgO1AcTqPw3e6X+QNf1F8p41XdN07KFRV58z9nqEjpBeYIhUAudftjftKvxVx
X09oetlhDxk0Nqr6cITwIdhRWhKRrrUuoyVNBoGPDfUr/g/mDjgDA6+LWtTK6yX0Xy6ME4LI2MuV
YhsnSKvuhJQ4qEOsGfVgN8EgUYRucTPEK8Se4p2IK9Cjwc6zGKCmr5Kqpa3VvQ8Yb5P8VaN5YOST
nZvv+9ovUzZ60UsgEB7tCvccJK27h98Nl6Hr0Df97LGPTrW/rUnzl529KrrC1QPX3hTLmZYShotl
8oREyK8XWbnOVmQu+Ep6vO3dd7U9MoH/OzAtiC9PKlNCTMMAhYiFzKx6dRMDymIy+2eNF2ZtqOO7
HYXCQ7VHPRSJUIRyPv6hVRnTFQUtmN2ddzZ7r+XbCFt/toe+PwyklMpOS6TcqfOkcmwOUBA8cVbN
UHt7H9lQwMhfNmsxAJG66NjDJRaUZkzExPwKiJQoLcjyJG9lXgznrs3ln4Ch4pKohDNfzAV9WuvE
LeURlS1r0h+mInkWLBWf5Ie1pUlI9rR9DDZBtfavZ09XxMP8q5vUsGFAXQ/UBaxwfAcl/Di1GNEp
1qcQkmTkkJW6I/qBqfBezhmnmVOAaA7s9d57DKjSLcmcKE6xX3bntclT3wLEvf/Q3v+2KsNCPnTm
N8QukYVuo7tohTgx5LyzKaBOzev4iShSxaEnS0LsnIvOW3CJSZ17/4vM0hFXlngHgjzGhwMJPAXP
Z/by0fIveAdDyDfbpsxPgDWmflq0NAxbkRkzNVEYg1/OgY6H/Cbz2NIo0m5wRjrRt3n5OZ+kGy+i
M2RcZAM6kI/1hXq6tl+CcNmYm2W9MW1sXSRtIR00rWj6AGkVF1olCL+QYeJK3XVFXIM0ovs18TgK
E7U2fOJshj6nYwMoKlqmBjv9u6A0A1T7YG6HA/MubSPZ5HHVUW0G5qOxjBWH4IFg1ZCVsehR9RH5
aP1JuJR2IQnhdoUxAJFY4SzZpQ1f1jO3MKaYIs6sGZJO1VZRIc3s/rCxfpDzWFcENrdiQny4zs1n
pCKwweiLPo/Sa/YT/+P5scr/P0oQ+59uu+52a8zwW90EPO0glvKQ5coQQBu6XDTV+Edxuj3xJDTG
HDFFmtHc0ktBeQh+hmx9cB1Phb8LBC2Qpl/cxBihlbF4D/MBpwns6HfoLnMEoER/E8scU9bNgTR6
jEPRDxRWHBooVNQutgESIozy+Dk1TWBQHV4Lg8DjO1m/PLOBWqSIt0Ku+Ox1+DpjtiI8A9xY41x4
JubM1i4JOh2jyIKOTyMd9hyW479XmkDNiRhRNdDkhOOStI1vzA/aFdS6Hw5iV78dY1QutlfWCehS
svzcIY1c24/U8bLCOl/QlD0vyfn21dQyb1opT4+x0A3McZAVg1hh4VFWh81G1bKXd8g0K59SwENG
0ZkBJNyP+vhdrrRuCRDjjhgAXy5o2oh/GA16ABw+2BoHR1X5Gd0v7YEUVGeLbI2uGkMKepJ+qdcA
bMY2ZQNAPpzn6jorHj61apXZ23cfUYJOlHwHw9Xe02OR+YSiBYwgim07cEzLKP4ctnUjCqVIgRQU
CCrz7JzHQj20LiygXGStk1vZfHy/EV+LXuzuBw9L++WIGvkzV9zVuU2wsTARaLmnjfd3VmsV462L
gQ58B8uO85nO/lCtUsBKCCuEXtU4RMA+ddkugwX2YPGurcmVgYyQgsLTZ/nB1xFyU559qFntFpvj
nCUOFEH4Stm9mLtBOYM3wgDZmWLrqIVkTR6cPZYLpVrzmi3FNjXzguFED8ix0sbhgrgVvNhvm2NN
fGgP6FQgL/4tsD3Nmn8/oWFPafBCwKEm44qmUJXHueeyIbA0CyXxhE4rQaYWX5k9lUmE9UzX1Vth
MUmy+sLCs1zqpb+4vbyEt8++h0wfmgSITfT4l93+ubdg4/4a1iLMANzCBy/5k/TlMkKrieTpbXE8
VZeGGEn/hZLOiSCVodlOX8OaTnhEdza2VsV+FLxg5k5VO94/V7eXaln3O9eu/syT9Coa28Y3AnTQ
pASyn7q6Ay32FuISh89cNJDfoTYWN/trEXno9EwwCgopwbcQA7B5iT59q8ddozB7ZLfsPsmnXvj1
cmdDTEuHVb4HvejRGxa2gc712/H0vFfzPD8ztCbAWmKfWdrf5WxFouiIjzxMeY3QxAcYKZIt1IEi
PJQZJeVy8q7Ekca1NM04KklI2QAX4IOHIpE2gaeCMB49JEBmAU/XtDGLiN3kjQFFLc5SrnXn73zA
hHyTzzK8wywGTNZ4MbL1jp7mZ68sZlon/xIl1w66s4EflvceyfNiS/jbKPchD76FS/owlhOmkBtw
w130WfMZe2jDQ3/qPkNdLTGb2wzefCOR/iKxtcMao75Zix6hrSHvJsd6NJfVUtT6de+J+xWNEQP4
f/ecZJGuLeGbWn2XKNuN+hjhcvBRj3FXSzEQjLM6pVwOEuwaFbEmPVh26VM0TfepLadPqhjtT2m2
gajnnBvg+lzZM2V7CJ/hVCNjuKckPj5PnxYaWPg+lP4O6hYGvwGb/5qS4zNu3ZZxftXTwjxr2n1P
Mw6UiOVjRc7b0FJWXgRyyEgoYO6c8LU3NRjd12VPmZtQbts+rM+MIC5t4kLzE4wHrQU2BjIeKXG3
NOUjFBGhfZAb01UdA2/6HiPlf9rQBJsv3+9DjE3+C55X3fo1g8g5Looc50K8Uc3IYg+B2fqs223H
+0jcPOACyy25X8vcnzQOnYdBk38DmfDgNEwN2MPY3w/+CVlzRY8u6kTuAh/u/MOK+D39HUkOwDg+
lrt38Aam0zlxN0rUwxmYJ8fq1u/OTMz9hv04NuF3T3djK6Ogp160wAp03AVqWXGJJ7A61UfPxsSs
vzrGlV6S0C2N2k3E8uUnvqqIvDcvJV7HY6RcRMeRURzeVEQJnIA0Eq5xogE7UcAQiNRlX+jQ8rHp
GtDhivk16jQaRZEVxCOFbqT4PuT2zO84WmaEwXVgDJzDXIPfIZxpx9Ze/HN0zTvTPLY3NZGbwXZI
NazAZe5AAaO7V4IVgBfyFdMGi1o2jbK3Dajbcl1xbmUrIoEqjX507/+zwz3Jf+HkJNa9Oz2aHpnf
PwcTG26Vs+i9JvTlTNFCbBMcGb2YzLHYB4iFiLrKmJD4m9Tq0eTgXewGPm1+IDrwpGDm0Y5FlmJF
wAGGfHdyyfzFMUsMFhT6yVC1hEQS+hxmffAA/+HzIg8ZeSJZ5gFc+RIJngrAgdu6/NVUQ07iJIa2
Yw3Tc+aEBRB8J/1LL27HOiKJ6R+uJMqlv0eG1R+nDdjKW6zwHYHBihqXGfaNjQtk5zIBUtDtr20V
ZjtCrbsxA+r/Rn0uBv0rhF3w2a8Ye1kjkRchPTcucRnkIgc2ecUpB2IvFcsoFbX1/SzDpDkbiYWN
vcVGyph1MCl6urOWD3LPn5XHr1KwwoFlN3lX3PF4WZK8fBKSqluKYMeep73KFZPT5jb8sD9nK99C
mA5d1d4EL9l6iSfts6kh63dghZ80CExHl4qGVjgMeIncv9yhIkNWbDMWPXstW0kj2nOLZn0U8X0Z
CU1SRe4PipVX+dMZc5QPQhuFnz9O23fMIF+IwD9MhhT3DRTORg7RduhYoQ9J900FDkaYXd0TQgTI
wVSn7FmFYBqnAHMI/zyuv6gDyccdnar5r6L10jR31c2X/hQ6rd8aHJ5nPEnCRfjfAi5jJkKp+3bK
Wgr1AKDr7v9aW9LlgoMKR16n1abcaeL4F0qleSE0ZUsLNVfSpNhUsfTR2NctBhGzpSbf+N9kyehj
vd99EuCoWxaoVAe/7RRB7u9G/g01tGyz0DXKfSWnCclmWz4y/HCrq162AmSUB3p30t7crMtqhvTe
ihOQsgxCCmVLPLTf4wu6y/NwzjZ88x7qgYC6wZtR9ZU12ebgA1Fxlp9noR9smRUT2Q4td4xsUFO9
Mnr9xC42HaP+irl+LzZ+VYJLmOdvZ97rurnS5Q9waXybpyz1KZJoSESnlQ27lWMfpz6PlDymLtoS
yU/4BiJiVTqn06WkotjbHDRyptXd8KEnrUjBkDp2vjOyhC0AuRfVw/yf98VEpQpd7Crj6OU1k893
R2RRabo+hPO4FjGR7tFgoX2WwHc/AkekPHH3WdplWD29WaVeclPof0mldvDeFFYlgiUXEYEDjnoJ
SeI+VrOaUya3tdqGgj+57vcBmRdPlbdYnvrfIDifw0vRLEEnsb7w74SklG9Uf9qr1NwzgqJ07A5i
DeEfHjt3P8qbAzwJjnId6ZtoVr5ljwlKWyHCqk5DQYQJqWRmJkowY/3DSqijbipseLOcMsOSXQoy
W+kNOOIc30nNNFkw+BsGO/pq7t0NpzGx3tmW13mWdTIreijtjKIHNq60nKKXn1ZgZyoGZ3H8Jutv
wS4PbCfIIdN7MjrUg6sAqw4ubAt+FZv0bphjFkLVfADqxyBHeFSXS2V0HxfsRBHkKTJZTb4WPL3O
VezVcHiwiI064Jxmq6X11lMhmlOepdIZQLBaqbt0fI897r9NkXkaRGA9/npmqSzXnu+il6cCpoBH
PKfLewA5cl4OHwIjQXSrCwC4y2EqSHGXIyTuOVYSafJHhHrwKyVvChRh78p0IMnKbm3u+MHW62g6
EELjp/JZzO7ufIfyAMh+qptsO9ccIv4UrVnSlawVkdbzo2/GUgRp9pfMEgaLT/9zsq5WXUWE+SxJ
U9cgGwmZUaHpjp/Br55VagfLy89GCsuZhpRUB0SNtjLs1thbOe5LdlmtBqL8HFsbLSEbW6bTJacq
WPE/rpoWBX+DvkSdb1MSuLC2w5ZaNj9P/P8PvQPtmeTDMcZxXY+yFpHVUSLN48bKKA3ef4Guvpzz
9NIkXmiGPNdhGCokQ4Io6crZVk4d2XOsraenAdnrXA6HRn0942GUZYhUtpHTe/7ZsdTylcjrhBgP
lzdukzeHgH8XxEUYpHSxMR2fv2Wggt23t2IynpaMg+aG9ziplSPud4+gPzlkjRbtiFEPFYd7poeE
E4na3OmCk1wvib7uLG+eZMh2eUx5Mx+CKJPfnpE14CUFsrLSDPAZ5SX923nmuIilmH8mF86z9AIl
cHWIXOxPDxFcVs5E4jMhfRJHCRxh2p2sFUr2z4DY2P/0hoGcvAG1PsKboupT9oIjZennGwlw1hz9
LoZ3XwDuYrAWj14+WiPTkryfdmjVOxh9kjeGLKZfDS/gH7E/1Bt489q0tg39B1oZFmwqSmmzrj2p
AZQ5rIaNZMQRNW32hxuK4Uc/Eit9EF7LArluRnrPmG+zYDersLAk3Zlvs3BNmP+wUuLPdT1RP0O4
BYM2bv+fdN9/kyU/BSlSCl63q7wgOAEZlwZOUTYeSgKXEB+UCdRhIPXUFyH+P3ErwMgjow5crpes
q+a1yJZD3DHpdbrrG9RKKE8kr0pQYP/6ha+a0bAElSf+VQ+vxlmZ/4Y4mFzpdCtfC/gpFvGt9bUJ
A19FZhT/b6F5aPnBdeLRJsf5GLozCE4qX7/5LlvGtP19HmnhV3TOilHqr7zxcUqsyqC+77m/r2vw
UgshGB4kA4NH4I6wT8aZixJCGEZd9fK3RiWeVwmcf/ngXLssb5dX4vwqtmfUafsLxQK9kKm7+xCU
65M/BayhjAxLfUW60QOaIofrOm6Ba3LEkBmMSYxyLTKcm2bSyCNRnAQUBjhzM+CycWpVLJehvpBb
/+c9y2hmpSi1Ov6+9mHaNmso/CSPiHZ8nurUsUGrjWHWD0x66LCexv2btRTr1AsHn3VzTvJ+wxgr
4/YnMRJWNayD5BDdd9Fcy9yU15QWIY751R9MPLjAkUwtDi+7Pe4kNDt5EYgV8cRbnn/EmboVCN0U
RkZT63sYKXb++jUbhlmfV6HCWdaWnhqzxtCGQQSw1e1se9Hndea5KmB/d74ODkYQxSR3gLq4RV0E
8LMYEF7ZCQsFK/xla4sHkp/eTMGwZM4MTjYIOmJH9jL3uJ257k7k1SccSSSWke5V/CwcsIfiDfgi
GpdW9/05bTPIB6FZFuYI/FCjx/6mAO+A6FD0F2YZuHzbSkyAyj8s0PuvUNC56gpnUHag2FklL3mj
7UA//4CeGQZwJ15NAuymW2fHvqpW+ZQ3atEnVavA2hbYajKxTjdsbKj1O7rzgr+PLn54WoNEx8b7
thTP2wcuSFnRlCUdpj4agpinhpTQsbfyOg45wCTXSTGOxibR9UfpvF3VbBfLLUZHPhYGGWhvo4LO
SvzS5aEHJNxFuqYDLdW3n1JDzP7++38BadLaWRXX8ZIrjnlwwb1My8J7Ev5VNEYBf/9xPaD3ogCm
zf8wwMJXFClIUeUewxeuvf5GApZeQXkrpdpMPU4r2D9L6D+WPAgejKyj+zHlvk5rXJmtenUPCSxV
9qHhW+WMxsmi/uzIP+IR4oLgSP5a2XNnB4x4fDF/jCYcgwsXrzFKRCHgOW4e9gZi9+EAE9HgfrEQ
5W4jIgmnFnxeYUPprhm38lRQ8eo2lKyW6SK/jnc/xzn9b/KUVz6pmwHsUSJYrNSn1igjz+3cpYA3
PZ5m7r8w0RUEyHRULnU3iRp7Lfi4DthT7NZuA0YH8xxyTSAya+F5K1uNH2omqRtFTEFs7MQywPfs
7MXyiW0tTG/nK2pjO0jzOQp4+Yj8A06uedHpwMtKxgQxNrgjCtmmX/MgV6DMLJUy4g2z6rQfDMcO
8mLAV87QBgLZHFww49o/TyzHok7SmyiL+/wgm2pqw4p3vZg81OYnpfAhsEqIY0Y57vSNXuLihmDc
JSY5voNZJX6Axvvs7FHXFVMjg2e+QwO4hQ7xNslECvAsI8zHaoILnG+Nazd+wGyvtN7LnoP9rWuV
lcRhA9luVA4/6k7Q/nMVIi2LY+jeHHUJJExLvqgYVD9HqKm00unK0VDUVoPCzdCP+GIn4blagxzo
r1P2qbMuFhkHRLGJWUpWvnFk9Vrnvn0+uRiNG66i+KAwhxO7JCmump8EuM5V246qfSSeliBbSUi3
dyOEk1Li6OF4ct9Y+CZuOsnwEySjlZOw7Wi5MRO/eobXyKakhflDYxNA/fF/9InYEXhdg/aJOHWk
Gjysost9mtKfnjZwFOpiyRqivxnWkqo8qkRodi/q9INE8nrasP1NQBwtxEW55V9WuhwSHOG7GKcc
H0wRmX7ZZKhR4xib0vLyrk+mjTGp40RuEhoAcuViw9siwDPqfcXTqE5AQ7cwM9hSMBG8spnoLXk9
35rH2Y2Nc7+XcyeBizIYGcY4mBXv2qtdWlgkcPM6R1vCkWZltdIMh94jdDWgUtuPyuiGKJ+eIP4L
sQOlhoiPgceEHR1YF1nq48AdrBjlPO1p9Bl6NlIJoumQXWVKdIuU+ePBf42CECuIWb1fVLJSpWpA
rsWJoM8ftxv9XZRTdE4SrVt3qE7fiSSW6tgDJVQ4KbVW95FyIWiC5TWKvZRBLHLt6qBhY+hwT751
L1vZEB9FEeU24Vq5F2i8j4fEaYfUtnczHeqkK9gKENNVj6vMRC7xGRUvjwjkVcis292XSiuO1EgC
KqQB+Ey2/rO3jA/gT0A+OdDP+CCE8HfdckywALRICR6IeeDbD11YH5PBsKZuKRkig292JnaKMBan
5rbEBDHLpvzjBpDKKtMrTjGOsc2yR0HV84iqD8Gj7K9v6LGNSOzHxgSt/s2T3Gjo7ZEn6ZVYedTB
7RC0U68U5ToPuK63uM4FOvGe63oAO1fo5+sJy/Fz4CxJf2AbcaE1RasWj7pg3LN92+uejNLYfCnh
6NbBechSllRisCtlylwHKb8ZmURdvf7DCGMaot7C/GzIt9mhwPDDaxicNwGKVFvKB44BvSHG6lW+
8i4tjXjrZIuPNx6jElw1ylPUiX2YQK++0zkfZCf9+LMpaRTKW1pPzdc0rTfmNMu0oDp3YYjCLLlp
deDEITeouEI7BDr/S3FsJfXgly/PC+T/iZubDxjPBMAmXOrQWSvhxXEufkvbo3NQnSJNhhcdEYGu
CAWP73KmOrUVDHdAyHVSjBDu4R1dRcDcAIcanbaE1Q6CPWlPFdsQwHvwcYRUlZ+ltYhgsDO7kmQr
nAYm/0Dfs+SZfhugoJqAoC1nxLuquZgk7mzjFmQXuTlFh/3vnPYcFNAhthSX/MyQdpTJg080cc5a
M4/MRRJkFGmt9ciXpUOvEy0Onc/9toHPxh6OQSoyvIqkK0RF0ti4x86n7u52Mo+FwPzL/6BwEG43
ngc0v3ZGljabhsoD9JktgBoi8BwQU6u93TZvf6y32htHtOlaC2RzsLoXg+VvsBQFtGWkZY6E3j5k
bBzbcmuMyXmQoBmYr2Rk0Zg7ACi1DHu1N2sfq8fEyVasJerUiVli18BnvgLmgTzOFXRl64IMviQc
6cDEq7dDhqFcR3RhxP8D1E+LPCYeaG5/fksSWoxwxKlY0/ifV4Md2yd1QFaQc2PDErwYj61CXLZR
J2aHJzYoAFwIKMXQEjrMEOa3lBOtESaNYhnpNkZ5q9vkFsswNa7nlkXMFRmw1i6sO4JUjaL7PEtS
QOlJ/EkMasbqzLJkNyksUZIv0wvQM9pef5soGZwo3epYlZ/5vMoOGIxkiGpsKxau5a0STfOPNKDu
oonmnQsXRbra6RrqqgRZ5xqffc8XHaNLVIQzdZM0UNdFdoCeIvYhTsyGHTy7WBXq7cz+JRyV4EPc
Ot9VW5lPKm6GDTyjyXBKY8JV7t8Z7ZSsvtYrbTwSP//0ygaiZl8jNP76c8wB3faK2oB30bYZg2f0
rCzUKJV7lHrojhadxEvY3R6tvhQIsn4HdnMa+ssp2s1RlKcVtcKj4wT5enhGp1+syHHnCxqTH3MH
VLpA+ysHjIQlxzbY3HTYGuKoFzR6UdigyW+2hbX/8K5RXKI1epdE3pMjGK0uOBodU81AZJXHLt7Q
5TgO3cCV+S40bUAmLfr/HQ74M4eDzineCRkDnCxqu6f/HGpNNSkETCnHj0jPbeQRqnAIfUCb2PP8
IIgB57PD5+5tSpPIZE6wAYrPzhV6wk10goixOsl9ZD3ISp05DobeEJKRBEMwFOLFh4iO9uGTspma
nf6EXS/R2uanTTVKwhDC5qUbWNtaI1J/mwxb6RAqDBAZudT3l7POU7+xZ46KyV4Im0PVSP3X5+kE
d19Ky7qibhwFEusd6ka4cQFq11pyHIWn6nCJGNk4ftVkFJwqz7VX3G72C81Zhx9L+9KGES5GiZh1
qFsMabuRIT6AdQmhOBw+GCNfQYPUBJb6jDTOK7LeIb/bIwY7FIF22Skn+clAl4toOr4HwpH8Uj6F
LnE/ior/JbqAOquBQ5ypDA7Rfu9Ddsw2sIDhGsxxR/+31+/mT0qyZxPiyEkQx1uf/1AcWVdOArln
TVIf0dYhru+ydMQFasYU2uQrQHhczKd+jPAdi9L479CgBl2ugJOvAxsJl7zxRLu2sbE8WNup0bxJ
c/E66ooSpLLIyZ1l1j8vaEzxg6ZF/xl9EdMU6wi0vwMElxFJxXqKSqNPVgf+6D2I+yrGJWHh2u2R
NJO7Mqb68gYJtPIhWj86HiYf2srg3B5UyYGL8l3qtwQ67ZbXNNjwphO5lZUTD6j2A7oIbI70q6Sj
28/RldyJk3o5YLnxD+A3JoebyWVupFtp3+lJxwf4KemhVe1tzvBdqaZo1gdEnCTXSEPWRNpj++Wb
YiRCiPuvoqp8D3MiSk5z1K81bH3TwRdJmlSCqze1JlYwFJ7NS0GO+1SKlzi5+cZbGEFq3oK6M2SK
g1s4YEjQdORTEw4fa0LGYVLmFm5gVCbwFeKj3sdLPWRWrNDCOcXdCt/YaS8Go0NbvMygM4XHJciY
8Gp8VBocnCz1IQChNTS8rRmaLAqUa0I+m5KjpXr8bD//HIL5XHMrowjL2qkxYZaG3ao3JAf0Nhdx
sxXR+jsSTTMIHudu7J9/KAZym5QhtBiT7RxpgdYYX0NZSRuVAxFJelO1OYul5YqHJ5i4QBVXHN1m
VIMJ4mo/Mk1EqoWo3iG20rRxqhngI5B8uJdW0mqZnyTfciqVsMmDNCK0npL0JRd+iudn7rCWtw4z
n6l/SdmVh1xpD22lWPBbwlgA0lTyYXgg5gfFghFOIJN8Qswe+fZ5pVDFuKXFzB9sib4Q9XBLHJL6
m+40Nh9jg+j77anRWsE0Y2bURQORKXL9qsFib5J+W6t8WvgI/dQLi92BysKxd6aPMxf+LgoNTthW
++wF2fxNKL+SUwPnTofsYYWAdtZr9lV4Ujnym0248xYH2pwrLSTcJLbPUrlFCkLs/a7Jn8pc7Y+s
77umwNK2s1JZxEuxU5GVEsITvz4zSJWPAxFDHbSFwcpnKpxpD7VVYRjWzVkRRahuueqasEIKv2MN
sc6pIASOoyRpJBP29J3nJztdS2jqrwrf3jTdI4LgAE00ph/J1n9XBjoYGlXVpSKflQv9NuKEyyyR
eVCJpWQNmNo/pyp37byoWRwbBV4ZvhUE/Fu8ERVgu+mLmKRJ6hJQtyz8p0ID79r6keg2/1QzCD45
Qz0EXIxmo+vsogHobDWSWFBVlSgE9gMtG6a53BeqbYDlDStWNtSXdBD8kUCY1yctWq5mEnS3xdHk
+125AJoN05VrH4CtXhXK+u5vefQYPOAjNIi+hr031IW9uw9I8pe6x+D/NzgqX5Z9scNkH+7yhaGU
FttKdjV4J4H973tASUE5RnkACFkcv/kc50MyZ6lidKFY6xOK+aMvEkiO930DkIp+Z2nGhdBfzaAP
yQCjiVEGIAqEfjQNdy9R1FDQGHnPJKU63iiO4TZL/xe6H3FjrMPu+E2awkaz1KQjbKORrHuSdG9I
Iokz4cr3AmFg8Gieg8HHOofFAeiL9qlJTKLMKyi5nxUDNj+t06M1BX3W+cPpQQADG+qfzkp95kY/
VUlUKhBxc47h5Ih8y+2QI6Xebli8tJslDLXjbKwK1z1GAp3JpDR3Y3ABdqMzY1/WyOdBGLqcveWm
u+YUEbmhDMQIDz84qQVgMbx0CrXqVu9oGWm+s9X0WCV7H3IOKkwFI35bIe9ah+jScXiznRnGuWLf
E+iwDk7o4XvRD6Dk1TfpYPEc1eoPwURdbpucemjagoVcuGNM3F3GflKB6sdaKZ6Pz8Mc5kyw1lxZ
AWWR9u4Tr/vUlcf8dTxsocTO/yI8fFCD5HRwxKL0p3D0w1As2t+rPbTuUdHdeQPI5XoUdXx7EBjN
2cjq6nvXioeMLJzx7BTBnQIN0iRIpgFy8HO2lBL+1XAXN2zRCjgM34W8Z2ijUpSEjU5jl+Wa3pqb
uORbFWBegiszpChlDAmH0pVUBlN9xBNqBx6afl7dmwxI8lIuQNogaECakmCiJqfvEE2rOpYYbobr
cOHhPE1YPRT78cdJ3Ioki5cp9j0XDv+CnmKax95fiC4opqahvQGT7qCtrMKlejKyeCPSYUHtbNn4
69fXEsvCijkMEIQh6TjulBEPHmCQATbrVZQQvU747UrRlNRhbQ2DGRGQyr5GGWr5IYyEgnvxVJJR
85PgQg6/E3nRR7zryQ0gz7uwFvkDewbtUy3hM4sNhPjxxEFAJMatvSQZGJrxsh7WNM/++5GQCrp9
1BTe1zflC6/OXveGgjjbxBYAAje62RME/n65OF8BUfnCAChCXAl9owr7PcvbRBumdItuUPmQNCIn
b2bdCn3rqlQKD+4dDNw7p4/wKWvNcd/Oxo6QAt4JrPbyOhz0w17j0PaRvzqAMBfF6DfOMmZXaYOO
ycboQUeEZTeA0YXQ+CI3tSGhhQSXagusDsFd639p/kumPiN6ZzrssJZrygB3zJuucvrw8VEwoRyT
1xMi2bDRIWZLjq5CBJ9hoinH0QLXu6fTr/Torn7H6fV7broypnL6yvjpWjcVZn9aJTo5FkyorqM2
AvJScFvOU9DHjJZkZmxubK5l+4bcqHkz46xAtEE9egIGY2URyfiidMHtBtRZVspnH2sYQg1driNl
JoVKKNt/QoMJ+ncdwGMQGwG6d6exTeqeWCoZyx9ayud60eRMTatniPatAgxYzhpaw6EU9CJWto+G
itpnVucHZ7Op68VzRbiKCMqsgQ5jOAlSrwiOySQvvcz+spNNwFNKF+qcfgSQT29U7VxSlihBJeg6
7LBHiOjJFAIrU39kdII+QwmMk9lpbmAMLiV3ACfbr5BC+VSpnISv1loBBy22XHPXquGz+ZBEmE9+
qVuXysvsqgBUScB4dRJ+IvKZqOsqH/8eiV1FBh+i8wbP8oY5CbK3MU4YSjlBiYx8QUjUPcTQLju7
yIyg+HrA6CpEPr4XeQ3tUZ08JZK9gLrqG2nR2YP+fT5g7tN5qORjzoGp3WnmyIzA6YAaYshCrj3m
NpV+mozX9aHXw5ogTqFSDQzyBS5nX1ytrn8Y48AtxIXNj0XP9m5XB7Pp+oOVD/sa0eltw4hSL2iS
keNhW8BvcpLWzwlgwzmtYsD1BF6YarHbmtgq5BdENwAXva9qCdp6NQCivgCqRnKD+VCI1Hg36We4
ajJKxZwjZsYnJVE5/jAYl4ITmbAcHaS/uMjROOuVQRZRQqwqsf7GEYKBnpSRNizkaVgawVO7TBt3
SgVZVPOa7EiEsIuYSkUfCVIxF2IxdwUp5rzTLkEK0ME7BE1dWHeQ0woI3HSdVhKXDI7nS22bUzDI
6H85J0fPQ18vFQk0U2J+tSnPTB7YgVXubWE88xVll6q1wCYKQLfyDwPou2gWLPptgaTY4vbeUY9k
7Fiewjtd5dFpB3BxRXvGmf3HDMxjnzx+hKdDJ/YNls1PVZrL2sWMh3UrNQNMDEvdN9Kfz3bgqoNg
1PvgRdbPhAHPYZEGinP0iTHP9OWuIX6/DiLRBg9sO/GksMbU1n+OBvJQohi9RMmQbZfdSJlZbIu4
ZjMPu5KoMhP9Y1sOwllge/4r9Nthq4QRrf+zKNjRAzmGkwcBlZgo2d5zztzFdHQchqnsbdqau4NK
7If3pR2RPwWIu4nzgDWWDe7oP+xY1C5SLUV4EJPb+Ms9Qih0C2PTB804dE1heczPJCeJFJiOQsW2
Yr+tTljC/q0uuSSe6BmjFtRA1lTQJCImxYw2LIGQTcXeAmIki5jQFzpLYQ0FXaY4IK3v8uP5/6TH
/laZ/k6jdRybW3DGGW4WVshaLXZv3sbSeV3EMrlFWjUTzx9PKsYjegNo4d+9DIUna4jFx0sH8058
3MOmOIXoQEvejQP2ihmRTZTl0pTI/gdYrZ3xqJ9wa7Z2UjgfGmBD6KlZZPBZIulJn0i5kegl2Gzg
9deblgS85nubSop8BuFaFxHGJZHQgfJCkbtyWW8VNujUnxI+fK5GPAcXQGtlFOkgT+89iXlCIF4R
tIHeU4D8WIIeTD2Rg8GQJiIhhw1VMKUU+k676b0cctsuIDt/9iQU7i7XCUqmua7+K+qtEZNSQn3d
kbfXq+JAy4aI1vXqh8qgsGI/4J54Ns0c0H41U+PqbuMf02WdjTPJ7Vpq8X6HISEWS0sMDmQ0LNQz
IaesFSE7LJGQXJ+ve9uxm+dMih3CNs98V7OJJ3Q4CLrUDM/FwFkxN/agDtgdxzPGTLHf3jeagWDo
EjRDmINZOxKA3cFQpRMLu+3b+oHNlZ+c8YQNiiczod9LeSEEC9LRgmhr71WYqNUqHyBIFdGdj1Wt
M3X0UC3WquUL/F+xjEeUE6B19Tye1CcrXYrcd+3CD/HE5bd8athq4ZGOWKYclr2t+y+zS4+drAtn
F/Wgd1oh8tbMNJsdICySIk59Z1Em5e1Gg+LxH8Dfg5A8R5AvGklGObtzO4ej6ZfVI/0C4nCJ9Cm3
daLLmWKu7qYAXSWUc5n46zVflV0T4VF+XrwTQ1upnIFPl04YGOnXMOLkdAgHt2xEW68pFLsi+qSG
vju+6Kd4JONl47jeR4v42646jn7RhVrNWFGPatZrzNqjtd1xwITKWHgAF3/CahdQLI9DbnndVrXB
hbJ59kQ7BlWqWpF5Y6IeJUZAPlJRtkTCbExnTELDfp1+z1caUoRNmXiYcvX+LDHTxdukDbUg+q+J
qOevGrIfsdwOOZmf8V4fXIU915zVAiYi+JaeQww8mOnKV6UFPP6Au+iPOTx6b9rXE75jT5CcQbui
myFtSD/2HTBTiAOWp1QITjdW/ioMaGWPpFPghVoXY3vrsypbL7nD4E85SJZB4/W7TvjtGM0h27d1
DWg9vYS0vhSiDA5kySkrYzx8FeoBUSaVnWFaqLiK0RY5MRmRI3Dspjc4rFd2mbCi7258LGD/o0Nf
WoqOZANklh+xrEWRSjeUqIKsRUEAbSunHDSX6+j+zu13GZJCsRNiEFqzUgiUhmL8fu/8YIXm6qON
mOn2fVTcxYQRpt2TxQkIgozdwrKyDaSAAJOYBmRAVdJbVxoDjjiahKnb4klv5PCgloYi6jWk8IpW
KxoPFcJTW4+09U+sGYfWjHCsYa1WaV3zAikg+pOLzE9gKc7j4SACBzz5KavNXqVztVK9FD3DlTqR
gVpVjQ1StpJVsX9NqbkYwSPXGShIfQA1cuzOERBxZRsUTtkH+ZDAKX5YZaBtegWN9N6V09UOCGE1
RJHkqXBjZIPqW34dsIdPvfHKXkMTUuEgTr3BYPkkCjvCdVkUsD6EpU2yUSeurlZSbxQQekK5JXaN
UA8IPNqLYy2M4LUwX3Y7uyKYy78boaWu3T4gOM6P1gTz3HYvAR1J6mmvq4IYAKeCjqDGv8Ph+NMJ
o7noHW0WQrolNdfA7fhFu2ntbOUeaNoee4TTsgjygolNH+ewRP5doahXa7anKuIWvo0EbsHum5p6
VOeIUIAjxLMq55TBbeGQZqIo4ay6U8ced6n8I5V3XWExzMUphnDtirLllnWjSDMVRgv90YwTNosH
SgiKpSbskilca13SPyxbMFT1ngf+TSfkEnkD1wR/IuPuMaOeXRTRP2peXBZkR8Whe0CoZcJUvZHz
k0chA8GtjsRDMkH6z/u/od4AvAO/gtwH72crKwd+42/WxnPrAhFDNWXHtxaROAsSrXUImQeSIqrd
BEEYV6MOORwaXRKwFNnQVxB3/ccI+rINAOnOyX5M5zMGdtGCZb8hlRCbKNw3eQmPFnpiGJ0SLbrl
DvFg4tqtIKiQwV3YinGvJserSB1CRDC9SXz3bVUwxyGNCObMp/wzSLwLPCSrmtk3Iw66VAtiP8MH
ZkZrZMU9roZq0iqiE+NGwcah1gtZ5DD6+TrfeSEOakNrRPwBta5T5U8aRhlYTojEk1ObSsgTqN2H
SGKfA5TinJn17uuRUv8zOAKVbH9xN2MTD21RFgrfJNEentKvTQ97XriouPp+NXLDReWkDwf5a9ZX
1GVRMEtIndkAui4q8n0/RbY39d06b1+1oQH/ESgZtZ76vvXakTatuL6YhEbztnJZYf0MMaPtLK2h
JHCZ9O1RivixtKmUM9Z7MWiWGwDS5ULpdKw+2B2Mkw7MIGxiQ5WhOC8bdU+THb48QLpZ83MWAepS
zNsnbRL6JXwQXqGvWsVndwZCCPsOQAPUN3puMHyyaN2ufqAEN//RAefTP88MaK01SMLnOfA6Pd1+
WgvHyFhOvojtNJkt4lyXi3W5hk4kB2gMs/t4Jb3uSynNiMRpgoJwgxVX1Zs4kXDEmcKPwnJdmkAy
i9eWOtJYf6OnVe27FOKAYFbjIfHSFsZyw9PrwFXkN5hXlepTINRnIjMFboQbOLlcGe/argDTcITh
OLlyOW86UTDUcl/wvFfXlhQon4Cma3foRJ32caHebWvsLP9vAE+rRwMAEjLMYxSERhvmfNkm++Ab
3zOqEhQhJ3PIU1t0vH9UFx85/p8DYrG8I3geLyRHD5fm5LqTRtnvNpGVEgOf1sqMFTfAgVB1aTMf
PigBTpgDpWl+nrelUZ34uqAE7e2ycBOjgjOKPMAmgMdM2MBdinL+0/Jqb5FmRdhbhqqnBI6V2BKq
qreWtC5e0IDD9VUNj2ARkjvRlkIv1cyzm6j5QrLFc/FiLJ4dSkZrrHOMR9fUWIBUMeB2rgnj2wG5
plVXwK8o8WXNr6B8KD83mHZSQQaIbgm0D97tT1nQule/xXZFly9Ouit40XSxJs8WvJylQhAbAE6D
ETo8OVFzUZ9Hk20mtzL8FuCq7ce04/rajaXvhZJL+wUKkXgGnkfedZ2izgW8MWzwoSsNJbmZd9bD
I5OZolZWpG8Q6e8lkGV14PrO+9EVujIyNMX+DX0Q2QFImR/R4dG9cje+XXe84Luk0cF5/psKJQ+j
hvkZpLoOL4KohMTceXLysQciJcZw6EsASju4mITGRIC7FYh+41UHS+UHi091BmXc1R9TzKl0Ug26
qZRGsKcpJK6wkS6ytmhvoRvz2jlEZDJFpPZIriLvcaEebj2WjANLHw+a5RnzPbVr2IEsxuY6peLH
syoySBwYXks/k4U79IlNfBS1Sy/8ZMdgZs4+c2wGytayHHEbhSQl6FnqFiPtLLbdsGI9td/VfbYv
/T4L5Vq+bNcqB0vuGQW/mB4NnsqaLFAL65xXAPRXNMtJhH69/L/2zzst8IkrPlenvogahZrKJ+SB
9imlGyaJV88tq6T5nahKP1qFeUsCrFpKcouexbL3/tJuyyxVTc7rQo4pFYc/FDVdErRhtUT609pa
gyvtKqqYSxXl7HSBEQD2vJ/MmuFesmCd4zoY8xTcisa27ByqZJpF/fRdi8JrkJbhaFMhvU9M3lUO
5snltg4VJdOJ4fWJRfBUo6endsVgjlZPXuKgE9N9RY6k6RtHOChvXl23qDzjHwBIeRacXrAg7Kq9
5rGvMmJ8AWZC0wn0Lu+q8L2DBM/SBT7WeDKdsddPBaMRpj3H11nlTm4p+lvmLF5fLtWdfc3pRFmM
pTUcfdvkSO+x8fdO5mnm4O6jOTRizzB2cDItggsaDqW/7yFn8LGXTxl3IiIxI+aMARhrgvavO1FI
v1DlQ4csgHeLnQ9/xCXKAGf9YQbGhAceOxGL7tc6X5pwoDz/9sRkZKKV8jGvb3QABeFTjLBUgQbo
r4mVP/OsZ1jYuJklLpQtE7NmwdiMTTJ/9ZCmkxt449dRi/yI223EMMPh/UfcYAwIonCS90GRISrO
dm8g1bBqWHGsjDNDiPd1n2tytYpOKdXOc42wXAYiELRMrP3JLnneSF/UVXjkXtnb9jNStZgkD8wZ
0syIHRQjlcFG3F+3ZcAowgfjY7IxFyDhfcHv8BfFzUMMA2pNT+PpdrgQNRAxr6tp1F5fYHT6AZsj
AZTDOX05JXMLYw4V/CLBnN14sRskMakFcJR6Q/XLq52k1AOwD2nAWBfoRNDWu8vnB+AlJprv29UH
47lMMn9btx5X9BEDRLQBYXDXZlWAuK+u7yFmd20D6G9rxNxtG3kaZsR1D7alMKo4FrDF5co2SXXB
pXEVPeUJcJoCNYyf3B7W/BiUPH9P60h94YJCLjuh7DruuKUJ0viHlrQYi9v6edV0tsCjloZNC1zA
56qP/f1M8UmsLHx6C4pMlRMO9mn1E4c4pgJismq5cSYywBiCXCcTFrK4hoJyxNUV2SN8hQznGN9z
7NURkwIEEb9IDnPtEu3N2bhsgFSGfl3nj5tv/4lObSDhpTJn5Ij5H3m3WcjLKsy4Kw6Uuk6bydRc
qpBO9sMxW8w1C3m2rmOnHXs9eotOssb1XQbA+P1hIqsgUyq6zrtnEJrHlfbn+Cwm1U363lwsg6jL
nfX0wTD+n+jev9UNc5CSIxjVJJpF7uMbL48z/qmQ60tcHJJuQq9EFiJCTkWVMhM93fPQzyAGR8Z9
lCldPy53OL8Hr4qALZSchwU6LerGQUnMrr3Y9rT4xx63VwwX2w0zM+HBJ7/34sody1y1VpsUhrKP
hiE47mGCiIVSHwvxCy5apN22BKYf5zXJLMttCz9C6vlwnucCMDtxqRqYUiIijjqRhGRlgxUptEzX
4XduIHgFUdhYwbuq0aUb/NVNpYnCohhrl2FRBpWbR+c9WyPZaSv7jwke5DqsgtAVnkAVr/xDEA4f
/PJriaQZHExVr6VfS/bAvfXUgYIEJR3B6bzkys3YxRssNn3ZIwzy7jQ8HcfpZJCODTU57hmMQq2h
9b6wItfp4r5FdTuEk83SDchYPiMh+hb/XgA10s1DSovdpS8bOe4fXAt3ltm1yFccmQTRrQxvLW8S
iC6G9vnjodSnt/9IGM79T7CFAUN7+9GpiqPlPtQjP7fK1DCEFtdw8m2Qw7h0bB5iSpi6YfOaBef0
atAYeWeBhl70RUYrphDE9FhGwbhVi/bFmO/lay5EieWKwN2H/btkNqeZ47qvnH2Fo34pO/V3I+Gb
ShpSw3H0t10/cbTGt1wplGivYkydN0i94mez9HihMiGjWF/fsZmvngDl4SJjES6tzmh2G008HvA9
Cp/Bk2gNDtaGrVfqleZNRPnL3ClfMQfSFywuV1lk6J+bUaNpjyUwFy+NMWuMx+03eyn7bd05Gw1G
o2vW2xV2DkhJFV/2Yfqwaqz99kZcrWOvfh1dnTonAwqZbhTZWptOSBdTsbodgCfnml6diRQJZDNR
/VC8NCUc9+0Xa6svHEwHyygOR6eDr5oCvnb2RmEweSSbi0FXjFD92uF8qTAhbJ6lNNJjcJ2vk2JG
/YY8xuPDG1MVfEQxp59xHgFT1sH8xgAYnA6h3YmEPSzqKYG33X158eBustakYnBhIxMpQoucY8gt
PUL75LF3BfKp59Q9xa7+Jvkbl0IfQInDBhAVkWzgCDXGaiEPcM0y5IxuZmjN1BGVofariPwxbbqN
2NvorusiJ7LLwIC04O3ACsVG5JUJ41KFmtMiU22RhEv7qNebYYbxJ5PelUelR7wJl7esTj7oxFCW
6o+wyklxtcvIp00hiT8yMesqeb2Ia6+qDXet3CWsNNFw0MzhWuQ4pxuFsq89KNSF/kwi8+NWrPiS
ILLpDHo2SKTxwV1quPWrKMJdEkUIWqSWG8TG5Cdrto70F0vZq2+IbeRSzjewd4jrXm8GIrfL9UpC
1yA8nbm+6g9Ipu6HGpDccjJlRCfCX61s1BoAWSz1dSTlbfxdbgQ/9YquDW8hKTDy+dETWFz7KhSz
DX9+oSc2iSMso7TuJnpyQsn1Q4vtVOYa8JDS0XNw3F2dmMS/oH3V3lcQA7rF9n8HYw86pafBd2om
5WDdkePt9oBIXM4+Pg53xM+a39UDWww6DeSFBy00vM/3HDGFUQegeoUsLd+WwUIQ7sLdMQ+4V1t6
y07CLdy4A1QBsp8wMAr8StDWuse6Yune9SudtvHSSYEkx7p2HT8rsJVCuoH7bUqQ0LW08XLTuWY4
jwt7QapcqMv5i4CG385xo2Dj77GswNp0wpIjw+5w7JARi1Z29VvvYCvMl4Hdol2j9YZr15Glenjt
VG+NGZ1TQZZC95MtPr+X8327ff8Wn/EmMCmIZUzPNbG/0OQ+rBeF2kyeZcHud3w7ozqg8ncKzSjV
kPBZBwpkYzE8x3atBiLjRcMsj8Yxxx8eENUB/uAKQQhF29SZ21QuYFVt3l6TXTR2QTlwejr9ljwL
sM0mFIHdSeJgPVNBBDdvzMjOvHWQn4RCE0ccRt+/2bSSesAa0pnEVQyLQei6yOaOH/j3uiytYosu
iH22J3tXR8nf2LbcgPfeoYAHlCtUQ/Woudex+vh5+JhZiTRaSqm0fomLtNtO3ATZ+w+nDxRaCZEo
RUgso+el2h69pDvyenMbKZtZL+jLkU+B95Xp6dqB7XjwUr8bTRrXhf6OdvPe3+Hwwj757Cp5JLVX
Oyo0DxJxtkV8O6L6HMsfEPOOJVs4LPteUGvAwewC4s7lKluf1c3lap4X0BuPlyjarcubkIcM45Ph
xZRl4d7qJ0ydeqijfS5jDXFx7GBBraP25z/IDDuhILGZoFPh3LZ0m/clrDye2ZwA57US3AveT4pO
o6fsZoKqxE2dBE4SZwom1rVxwOZ1B5DBng1h5rdJzQL/z/uvMrIhu0engwZB5TIx9QtgNUcfFuri
6rXvIRkfZVzcXwtCeYJ9cHt/4FQuVn/+WpDndU5nySuG2zg7LY3criBK5X9arlTZToUvjKOwzvgf
I++3Ket8mTuBJgDXaltSmi9wRRtyK2Vx3TuklyALGsXQyVdoGXzAsut++bKlUq5r8L6aIH8VJmAZ
31tUO0OIwdduq1SzjnitXqUZwWFp85VzEmhx8/jw8UgB8SiRJphFQ3OMm7CePIg5fj5ppQLUCpeY
xOQOp8tjBUpmsEVesopcKxfhuSvhBlnaUHOZXOeGi/QWKYYEJTY9YANBhG0IiCPu6V9jKZDNFXk3
S4pEpdgJS0siIQ/Mtqe/YSsnVb3mDGD0P0VGoe3+vP41F7bWd6MC/HB0IEwB+kLTgdWNShN30/Yp
fzzFnaNJ6yKwTocy/lU0Hs8GlEv/JFcxm4TKBhi7XTYxIKwWMF57ah4UiMQXw7vWzEuLe8zJ1U/p
jJnskEuIW1P0RUuvNpgUCDE+AcOk66/1UB3xPpFtDyTYIAqTyKqp5AO1InC4HDLMwDVwRz9eqGAl
wf6K8JdztkrfP8IiPVFsUiM/yxkjL8w+MzAtuiBCeAnqOkX0jvsoS56lTw5MuQjUFqOAgz8FQ/N9
1MClh3JCtPP/1plQTO49QJjTlCXBGBTLa97q1CAwFwfTFJQgGM86HqNihd1UoYvLaVPOVuJw+aJj
sT7JwgtknSMk9Z0Twb6vDA5f+cg9lEzLXwAej16lIbrrNCtZR0ffyLXVUBapNXq6cBMLlmUWjnZX
3WfsnyKyRV2IUxXJ8oJL9ySydHC4Ry5qyas2y9nyIJH6RDUGD5WIIC5rJRAXpxbBk+4/AlvjkEcz
kWsGHmMGVVWYaBzM5h7hjOk/Nq/Dblnf7UXgXiROTyGm6Ei7QMBiVrLL0hqVHMaoUXr3tdL/LLM4
SnqZfZbufqBLcEI+DVWGG+52txIIIpMgh/GqW/EWl9jV/BxGkAww+lX/xCdv4f86UXR7rVPvx6lf
YoweKnbvlLymQwRhx4pt+45FQROE6vk/H6XlAa9HpZKsmUJcxslkLrYl6n2qmhcK3T+nXFFXQTZQ
Uj7UYC04PkdUAAwWtjup84maFvH7GsdTxNqnmGtwZWYt2mvV+tc7n4/GvDKi7K/lpoYz+rf5I7r7
J8nz5r45oR7gGBGT6TfpkZ3QdyH2NB/hGSJIKN1bEceiKuxUiZKORHwzFqmfVYueqL4TfkcTehsC
8YDq+WIqZAi29Pq9OgifywiJsn6iMlYqp/TvXQaivVvaG7g3NExk7K5vE1Wf5ibzNwTk3Pssm+jZ
QqvQKGHDRzOU4QRyFJZ5igbfEmMq9MuDDZ9/BMSyiPFqnCPQ/doX7gxlYNtofd12MWbufj6V3uK6
yMW7e+KV5vN/FTfojv9H1E67XYZah+LGdYQRXxcdmwKhZKrVH7zCr/F1ktc1zGEikHvPfmn+EPZo
CLEk85hdOG7UwYSnFnOhBG0rOsUnwigqm+m4YPazdpwMc3mIi/NFIRFk0RTe+k0F8llVPenMoVDx
hskn2fVHJT5xA0AKhbQ6T9qkeyhOxDg4X3WazgwV0oE/J59KcI8x01u7rD2Q4BoKjzWPnxsHcDxf
XQ+BwqtpBUuQvyna98BuEoG0zi1YqZXCJx+PQ4qb36FuGSjRznvZxE9vtcbQiUfX8V+hGehN1m5W
LZTB6HpmR84Gp9ykb8AYCAvwd1MgLp02ovN8BBSNj4hXTkeCZQ2Dr8MiP6jQ8lu3350T2KU+kMl2
VbQeP++ZUJpClcLZDs97Fz7FfdowOXLFec4HBUJGprlRh5vJ12ZjK8J8p4NDWPR6g2A6rs5RmZ4m
5Wqd+KIAFLD/IUBBmFXMypftRcp61QKfbs0HyqiOjkXn4eZKy2ZCE3x/M4W4k0CZ1CTxGuEy6aqs
zM/AB3iNROTsplTlIxl+FvmEtInle9KWA5mLKXwNH8G/5I1+udecThFZhe4/qV65IkSQs95jVOCE
boOjqj5qSbM+lZgtTAcnTSef1p9DbBKjuYwwgnpOX4UFr56ThrtmAvUPAzqHKfJNXfitWCB9YNux
X9yfm0jx4FTyVCmSKydpITBQoqQcCXTLRDcBXmWI7tUr+0vkstQ0eWbefGTAkZ5UI/bRKSgI5wWZ
H4XUT3QeC+14DUkruRLR9rw4ZQnDHB0ZsUCucnIQ4pOy3xsnEjQuEzplKHN6yYJJ96Xnsq6kq/Cv
XYxDkzcEdo62NU6BE6hl1IfTg3nV/wcJxmdd4GQJISpKVfqTpNu+5WCaay9tZOvkANQBJcasllQf
hBRYCDlb/WnrEs7H0BTtoDY04wNN/cqXfMv/1Y+xBs38aO7F99m/xFoI9XtcOq9it0A23rZFu5vx
tCzl/A8BriDWsVjhz5AZ3IlwL0tSNnErKfC0teXP5qGvsKu92cZImObOQilyuNsv92jLaU3HnX4J
3R0anY7jTmWUzt7PEDym9gUkVEQLOKCH492SNESb/yoF46kM6m1APj/Xx89j9gOeG8mVDdX7WjLd
RObyhgQdHZRowsYLpSi7qp2pANc8+LRg/OP7yBJO2RzNwDgmrTASIWPhFR/RnsGwtRIlVsTI9BDz
iMJRqhl8Zcn+AmnTFGqhu6bs1T/xdR8hh8aKJzy+MY96gVQW7rzrg0jEQRHuvj1uWiMPzR7VBede
pBb3NQ1kjQax9hEiJZoH019OVUHQIZ76VIkBsES/Taqo6yAPihT+cyvgbQnigBd0httuRVZyMla9
nYbFQFxl+IlJMUDkljgR/9zv7NNBHSz3TQ4uyPYiOH5KftPKvly8V8+nPS4MksjnOrYgjDBUDx1g
NyzYZbUMStmEEsTmrK9Xrh79gtSHXMhIo9dylHYIVlSqAnQ+rK4IrAZ68zXIH6aWAwYdtSbIbifk
hsjsNRlYaGBvSsliTAdnk/ctrCizkpPYKVHb5URV2WZBll3qtRsdvN0GIHroOnEM9oeTEuXxfhcy
7fBHUBb4vj+24kxsIB0OhDyjPrTdFZeL4p7o5IPuTCANIRcT35jli8W/P5nB9KXytkAhYlGvUgMw
FoB/KKiXRFi6CVwoPubPTBBErtjmU8HP/6wDwDvB16RLeYqFvGKbLQnSuEjFVNN+RjV7x6gvn900
AjHemGtgzpVDDMGXKnt+hJBD8SBI9QmDsqTICc/IYA9L+miX/9rshJCdzHMSlaBIyG1Qt9lD34iD
lVCq68sOit2UdbSsk9oiZ9msQE0gMa7iIF3tsRScTP8OUeAvIGceaS2q7ql5JIT9n8iTA7wdglaJ
laumyae5PteBw+ztOE1SYXkicKzDrqeoHLXR417JJqIow9LRuj+OG3+1w7yWKpJaf/W+3F0KGwWY
q2yaMXCr0FRUxzCDIll1hYfTt4pbum8K/gPuuxUXQ3XAVMu7+VR7CAaMyLyyMiKxZNlT208mO3aZ
sQ923/8o6L85kUL9jIOrQlS99PkAinDmIAyhhdJONWc3OMEw4wsV15UC868+V3x9P8l4+wiYUlwQ
ypL3P9m4jWQfBlYTiS19mxOBzJhUE8R8ncmMf3fIv+vUUnr+wr943Y9kiKWkv2+WggHgJmg3V2wS
OxaETiEhhIQGm35k81Ph0kLVFErAn2GuQNHefii+Qf/PUO2fYLfYvRlFOaMPcpxxhxr7uMEEWJZ4
lc0xxDaSKnCqming85qtOZ37lPvf+9KhLw/4wauJ9+tANl9T4RccMP/Exie5dPp1u4AajJ5aLa/j
I+kuNO1E0YFvTdvBwK39twV1CA7EVrkkUG8X0Rut7TmXEwen+1ZNkcBBTPPdUywGvN0IiHMxagOY
WqhMSwnOwhAXNxV+nmsqIyOa18+2ftnp7CK7Wkypbt3M288EnwG92hdpfiOiR6BneIa4KBK1ODqf
PNQmUoHPfgcXMXzNYKxuHpOSGEJnq3M7eD0gQcoKIUJzu+Xl8dWCLXrcnjMJecYju4+48x1uXrWr
gJ1ZmMszeY2fo0j2pq9Ku0HhkD+hWshGzf/uB46jmJoi9hEs4bCZCK+76q2i86SzQtIE/ZGpTtYr
rghDXzI5DAQom97C8sLIUdwR5D1VWqvsItEPIqdnrVaSiT28bG5XEp80wACOHiEOz6Xw9HkXmzxl
72K37Nv7Ln+6SfbL5/0qJsdVNbeI4gRPgBmmfGjY4+9nKXoizJ0Y1vwsAVcWDa+xG7nYsYSwn/e4
JGlMbIez1vZ1asGJ5Fl/mOSPtp4w8AzvUOwL1hBEtD7Lbh29mbTP+ia+PB4lf0LAe52/2fIzOtoA
rvYTH7Qa7ovvJfGa4ZOakvB7i90GMKksIs54xFykarWHMVg1/49EzD961DxG6vKcfvblYKYzw1KR
KRZvhrfldyzFalu6du+agObA+zArJF9sHJ6HsUWJs0+rQKoPn63kyFXpEuaTd+kVxBNuUXFxwGLU
d0Nskc18nWgU9+e8N0KSV5PyUpsrP9P3d4lN0QfFqErVhLIMesVctGQHOVegIK/hEP9c6cj4xLHm
Ba6t2ZSQPTfhGAmViYxd50Xm8NEogBjW7D/NUO/LumzAmjCEIUY6YY0Gx59AB9M3pJnyzIvPsUN3
kuc+6e6ejP/3AED2OCb1RTe8gR/XmuWUD6MsYiGSPctPGxsRwmPHDRGWxLMXzKhBzkb6P8jqUmAo
nPnoInI1856Oi6pPSdMibXCRd6hHApP1NCg28cLRLujJtpXyJRive+DH3r7xZmF48iQMJdAZDuNF
fhw3KGathN7bMjIoSlVPQuL0A5XVpcb3CZaSAsUBfDTNYqRGo0UIbYTIKLr82C796az5+EiT3DOI
L521pXKtqS96L3J7wBi3sh2+QUAUAulsqjCEL0dEb1iwAR8vTQeCgVDSgendhJS8Hx7qEQ0Ugphp
WLWkZia+Htl+zhVBPvLp65BCQTQJsIGxEoDKTayndsyFo96ierVmtIf3T2v8azlxWBXiSY7ZrRHv
D180HbkWj+7HxKG/tFQzinG+9EVEk/hU6Ks68nrDRJuRPO63L4nsMyIjY9RUrYlN4oTW6JntB8kR
e0BZJeS+CXt+1pvKn4VRiAPGdPUHbwonyoLHygS0nlZq5RWwIoe6HXIP7pEtkCkBFmcntV270RM5
Nm6z0JegnUyO4R8AzklHMKWUuuVHCiOj0N+FqHcwnL68N6sQC52MoXsk5sYBttf5u4En9Vj7y8A1
wtVIpPlbQZDnrtGmNNDfrO/vyH2cd6yMoN5mwSHNMeAoNM8K+tQK40fswWtVIjitj5jKgA5yNm6U
wXHpPIMBtfJkWJOAQQGmU9KSGVCZl9BmsT95o74b3KiEasZF2Ksf5QAT2UX0hucEa0kiVUoygn3F
pbiBDm0Oy2F0mCUX2BUEBh62o4j6g+Nnb7Li/s4NRNNPojy0oL1f1RVAUJXOJcZAdInv1585d5N3
maACkiOITb8f1fPYKPiMgZY4ADHpgiXxz2I6zZQF4SiKQwg/3hJKHAxFDAxSQef37YyAsd5gB9Lg
HmkppNXZVp1fO+xo7IQtRtSzFltu0cDqVnMF5JmNMjd46cc7XIKMJ7dMGZsUh2V1ZybCseRh8IVS
oUY0sfili9kklox3hSf0P4rQ7jKM6s905hub+s55/TwqPIrBvSev4BadyakwbxdQ1e5qurgDWZVb
JZU0muxbid4Slsjd4bxeGvCN8aKfyKTQH4Lui8JtkrSLS4km7caykB6NMLqWXYjHslz40OCDzxtz
yywUC6k4jcawFEnID8omQp62RhxhbGJmq4G1Jgrd6/7BGW1b/D6EqZQktKeIVw2O4F0FVus+kq0z
2J4PoSEtmwE7DLrvPFNQTKExhlVeq3wPWfdvkJc4LsE3WWSQCJM4eKBrulN0fh1C46iSCCxpAfC6
LkBbcPspxdPdEeUxKwRNQvYAhNVcMHOCh00gUqAunIdi/dwCyKzS/aNdCob9PeHCGA2GniPrfWBC
T9YxhBSX/nx60rzzMy7fCD9g2/BknnCzfD8CTBU0VaymowzhKnYJWjGQ3E7fPBh8bx/8Rbe+abI6
adpWXvnVMgT5fnVI5kcuWPpILxJ1c3niPOZ2XGSziPNpSlsPV5wD3mSEHbjW+XCyu6+mQZNPZjdT
2IVpQ8D6ODr47cxcfr1FmW1z2LBg+U0At2OTK38zQICnFrhaUxgLu8q+JXmY/H5CCj7oHxdecBU2
6JbvBDiWWGu7bMZbpKidGdf4KvNc6ZxO/vw0EkKmYTrrWCHXjVz9AhnqJ/U76DoUyjdqyA+W/P6c
OA7284mqSEJOqtNKNUQ8mvZyIWTU6Pa2uAd5QVxude7s11llntQ+4CAw60jYxeiAAMC0jxMOEyc2
edc8+cZxFoxgUPSNEm2kPzPNTQhC8Kj468h6mGPcdKXCP43LcAimss1NEI068beuaRv+poN9eWlz
ywIwWtxv5iTjVYXIb4l62Xu1Wb0MbXmvNEDAsT4kB+16yBbKj23ZD7Cjsz1lhyhVYuS5yXfNvi+4
oT9lGCjUIQnEW6EDgNMLKU4KV+aRdFXes+0ZUO1BBg15UlrmkxImAmjza39qEDn4iONHLBy2RdjG
wKM/WW8Q1ptnhz2+F5hJ7C8URj4gAN9oveduVk+YvL3Wv9HaCaLQSylD4SyWAn4RFXVfAmlrLf1P
/+uhgUth99xmuxAf6zojfd0IFqlMdQpi2i689IXaP6y1oHX9HIE/tLgC9Qvo4NNCs2f2A1fRir+m
XthI4RKKQW61o6g9urDLSBlPCgiYQb71ZEPXrGDT6Fy4QsfeC7R9G459RUuP5tuJFVyq8kq3U8S1
OnBHvY1jCAPjgWRhtOHU+J2lUKfgPTQ0LFwKg7sqYDRk0gxqALSWPoDj7wc4mNIVfEHBIj0BruAC
qQ7mxY8BWJrvf62e+sRsynJrXzzfnyqheflLEkS4RPIY1Bsj4ig32RdfnaGzX+hiViDDnXBnFLVs
uz6VrvcIALFP7vDLfInj6vjKt8Mvbb+Qntp8jdmwifvtRcRKPgYoDHvdt2YE9vcB6HHyg8YCb8up
evrf7qilVqqKSfPIpxeqAvaxsqnB8aIbwbZf4sEYle2n8s+ypwrq1UnUmqTeednU8Me2RzwL/0VI
pn80gxAayQnJEnumpK26thqkNLV9i5W7AUlaHfdi80NmWlEmtFvDW2SqECvh15adtrC3YzzqPhfG
z6aY/KG0jkRGv4NpVnc9R1yoiAk4Czp5SillvF4fVRM0XVMNknFf32vOBuYdIH3rolnm8UpEPbVl
72D1co/V3hsLAMgdWC8jEnqGpk4b+jP6HosKB6MsHiZ+86p//QNIFxh5ZX0Mx87ubZitzN0/0ScA
/yvNlWvAlSdLKvOwe/31nuqs0HXap82/pYStfRGbTOK9gl4VAZcKo2wqACyeRXVAlDNRMWBIGv/H
GxcQqQ2gkT7lImuZLv1E7II1Ts8PLLbPUll0ZaLGSGRvwNRpFpkJaNdhtLGE4t1YIoEpK9fy2PT6
8ma99od2r5LME0eP2iSDGMOL+UxWv+eoTCWYj6+HM6jUpi1q3G+ktFFFeTVYIvjfTii3g2lQ+/bL
b/PURgL8XeA94tYqTeaAjpBDobVkyShgLOdxp1omhwNq795rkhBuyhAzcE+btow/DfgtlfmpX33Y
s4sVvkxd36QfYDYLurn7I+X3O6sW4hmcHmiyI0PEg0k6rdbkrxjTx2dAQZBbVMqloam1fevbC18b
PIPk+OwIUWOLKJpIaubsEUfcjtZsfQ3QYeVWmw1ToAV5FxOryH+84TVlvHv8YRLjTG4BNR0q/iza
zR3bn52rsLOCfunhvcrIjxHdRzQps/c7Izo0ey+m7iD09mJYKwi9YkqMD4s8+nHAiyTRNG1GKAyg
UkP9qPl9V78nzWkMi7cuxyaw9JgV4Npt/rdTFmYdmbjtXhGLp7yn+8EQHFU9JF6H1bRRLUaZGD6k
pjZBSqi1zwmOoyDPCZK83QwU8jNKwnOncibXOiUQfSeLw53ciF7/siICRTZO+Lzk2ZTcbExV0BLJ
uVVmTdara/NIW2UM7gBnlLFwXyDqscuJL1vEJDk6dgweeBTt9PhBralQCYl1TQQY4kVOPYO2+dkm
YNh0ZP2Li2aX9dlah8dlx9KO5Hmq9QupBUSXxecvGrxERchxhJfJVhYa4srUW2s661iXHr3K1pcs
2loG2x/YK/9HWsxAtqXkHNw0ldmPr2DkXgNNybpiUdWzRZp12A+tMNvVEkhAl+EKi5iN1W6NlUEY
EfBdzoFhHeyiYHEetnNaKDsI6j7DA8p3sKqRRGDUi8mnst+HgGr2/9tgLGERGI/wh9XH3TgYHQP/
IxYGazsrOtDyKleu92Hm5zp4bRD5c0JVaJSzVVOrqbUU1hZCGTYW/+nxvdOQj01VxlE2uDuBlyY4
FQ8kTYfMju6tc56Y3NYxgX4HrBA8iUZqz3t+2QzFmn0MZd12/Zs/zU+1I+2aLpNk5aBMLcywDH7i
jaJSjQjJhofM+s/NVhEaA5OdEQ6Td2ciOPJllWiI5Al1oRKaPfumml2XsBRprmq9VIFzqnlk3zHD
QsVCOp5b39HXsjAHBZOc3Crm+CmIyuPG+FfkzLLJOHKuiUJFlXUZQ9L/SmoGCIbB9/7Y9biL9CQg
1yWMYKjD8OosUY+w7Ir+WhnkoRyIKEdltWTGKSAfeOeOCT5d+NvdoM7C+FMTPp8RFF0HbwxLwZ2H
YeiVnfNYZ+FF/ZznSjYg+w1ebl9CXLuAOeTdUVzkY3ajnIlflihbpOYxAjkt9NnWmNtnvYxFwOIi
WVUiEx8vk+FC8TKLJlZO+sHJkgWln8VwKqXz9QBeBV7GE2MGEv4OWdFP+gwu4qaDUDHwb7/ZbH8n
R8Cj89UoboBiQPoc+rbfKLyWsvXMxeuZyms1DKW2Wo1TpVbE6Gv9vMB2pG77ybP/8GSBDDSfrkW2
xpfUxCWGy+z411q2LtNNb0aTPg4x3TtfXaA4/GyftjtMq+uUj2F920YRZK5LR65y69CTVK03iHAH
ddYCYzJ0hRyJ8RU2kH04Rsiv4+CwUwJSpbYOdWBGt6DCRJCbzjh4P+6vO8jePv1zFu2ZhTsw9i6j
Z2HcT9QxOtkagysPncxnHjf0xTbkLxjo3W2VboXCy2O5TPhiXOu9TA6FZSc8ea1uBTqtb+ZUy2tE
P0+uu2wXchWF60sb4f0jRzUHB9hqMrPrTBu0PxP2QpT1tgeBXEdPxkS4RlybEzhMpWOgHigfGEcc
YqMdj2Tal/ghYmTQY3qG9dVBC97tt5AIJzEHmRA9MPlTTm7dQ6hyINdim7WVqsxD43Dz80VkARJ+
fL0zbqfxhLw6/vWzySqmxMp8JHWiAGpMTNyquu4AJ4r97azxyMmSxu1d5um73fkH/7xYAJN1+OWv
HXyUazviBjek8/zvBdfYD2Yoty6N5hC9+CxMkcmyrcudducu5xAcVIQIICTWoTkAq/c/M3fu8Ult
6raukHwhaacaXJB4F7GMLQBiWL1ezQXV/lEW/XGySnB87CzBZwB/kDnBI6W6508V/6RCb7KmKEHx
xOwS7RA7UWlkjdVGUphImiMqTVDBf7pr8zJw0Q8jfmmLY48zZYRWieJDMvNbic6ZTRvQLn7BZHCR
S+qJ4+hT8fLvqd9j9qRFpRqLJVmyHoWTqRLp6tCpL8tU5ZQCCfE+QqOMfv0uyqZ23qe6s+r9QC+Y
9t2svX1o4JNUpTK2DblM9JtuQUTtHOb15toLCjU70C2QqboCr+tbHKs5ABEWxCypa4AjM5XAINPm
YuTXVvp7AJIxiQ7clapc1FN78s5e/BKNiLJS+e7HpiDa+t2wf0uwkgqcgABsf62Oig8tReOSY3a+
o0QWzhpza939I/hT1glS/jeF9QjY+akCrpACjdBKG2yFsQsyd0NXFmZAlFdm/oXHbjf6tfvQs3xs
k5phfbdJpSEy2QPh5BFHl65cC9+e742ksG36rOWdnguHn2Q/V+2yRSXmZcPT0lMnQPx0ToyuSJZd
HC2Zra52gYvzkkodOmLlZtzGQ3R4noeapq2lKHNgULNwsqF3/KwP+vSkG24C2nZg2l9JdiMjpJUB
6dGA6cLZIBV70ETK5DFUjF/eiWMAqf60ivtCLGdmwGZnjE76sygLK4J4S33bVilheJRJbuBaB+4x
mOGoYWZXm2N+HZV7gkHl0pLfy7wLrTodWuT15l877IP0+SGAYPciY0yKG3LjuWM92a76sITvYfn3
VE082obA8BEaKENGKRE1ieG2RBuQLrEMP6dJ46ErhSDUmztln4Ws/kC65VziDPmYd0xokJe++Rja
k31LgRX1uYOOLyq3WYkYfgckagqT6/JLKPyL6+p1YjZVkqGPJpduWZwQmT3Li8Dzl4uMyqxwQpbD
pDn0UUo/GaJxoQ3N6CNRG3albymrMXA+GhQaqfcwMfCAzX5Q4lB+sJCP05EOhjzQZbzAxe/TxuHm
pBP3B8iQmjn2e/lxrUJ4eeuMivqtvgU4kaW7dTndYCmQn067+XgUivU1eNdV8Iq3hzJMeM2SHwKZ
KpI8DtbTDSXc6t4EVDk7yd+T9kD8sr/1VkFPuka++CFlkzSrI5lAS9YHKmFcn3z3R87GuvQR+NUh
uMcfV2/FaGhgdh+zuGyLWjq8+2bb/aE+XbJB87WwJ4hgw3K0QMLKKcbEPNp7A41kU0EyQuI9n8KR
Dtzx4VsdLsyHlMnf0bGJ7I2YPoRoXQRWs+JRiHGDwd9J5un5MNdRYDDX0htslqU1FPEdLXdk9UBn
AX2VpXFOoHHGeXLUZy/3mwB+9lsaGlGH1JgXflxPPdbZ8AdIgeFZucMt+YDVGcIUrTqhv+btNHI4
JIyLritDDJ6nzzb82oLDxS8PKTf2UXkfVgo9lzpC1Y3dJn9w8Mfg3FC53zmsYHhRbOQmmU3Y7fsI
8ULCowt9Enc0mJRer1ccUBE7YRoVjH7c89bO3WjtRbDAjkej4vgBeWqYNpY/qMvrOF3z+DSGbCgW
PCBW87iC4pH3PWaQDpnGC7DxcXjqMp+mfWcUJwIRYWm2H3XkBgmv5+5I+shrZp8hLf+t3DU74bDm
d5CupKtiGLR7SIKWBXty4jF1OE0xutyd3byIwoJ6POkGHcbFv9hugrHqnWIxUfZjkX0b60tA0Gtp
M2+k1vOay9xMRN9dpebL8mPsB5iECG2ZJG7E1mqtCiLoiH9KSaBtDadfYyTz4Mw+XGRVwTng0F00
EwCr+lhtJjBG1+xos3tcauvIqnjwzBOI/jVbydKKfL4pPaAW0JKEEgJPlKlDTjvcs5QMvtReBy2V
N1TwIARvbuiDpNZ7bBKYiFa+QwIekom4x77hPA4zy6fYuhiQtpIGz8kbS2E7awLaRapZkZ5/LjX3
aq8ReSlHgj/nLeMpPpFaRF4h7JNNKY57uaAa/RyNFwogBSta1a5kaVbllnbXke0H/B3PeMyP2Tb9
N4bGPzmECjTbVAT68ij+BuyIevQ2t4wM70rueQ+70N3fBAy8qWLPA00a8JReZ7auYZU4z6+RMsUQ
xv/vAEcH8hfcEt4caUcE42ABn/UtbbIFjuvQC8RlD+K3Fpqxzpj6i6IxXnuARwMDq1XfdSRE8RYc
HN/T/0EzIFB6pKprL6owEJlUGEYJnOGjZVzlyrMBjtY3fiwq239cQaAU5v5iFMxGR5YNy4ZNM60x
RDbfBxKM6ivjl3R12NgbaN9y7sYR0JeZ30Rg2wJg2LbX0vg6K0CygWS22mS3urdMx4/GX9Mvt1Ro
Z4Cq5Qs3iNW1XLxrYPLhOi2OwLJSlqIY+4YxFGnx2vwAGJtb2RXjy6IBc8MkT/ebQnC2sptUAYk2
rHNNJxm+3OGpFMDYAi5WVPcMTW34dKWIXs3Wzb3Ah7fG+lYaVpqLf3jiyR6i8Hyf4MMchfvJzUg3
MvSQzYCG8jziHkCRMj43ZqZ+I6PK1p1UxCmkwkB7zBlVO4bsx03zQ2UoC2vshixa65RMhwiEHq13
3r8/uMFsNA7vZkIZG4HzRUCEk3cGxrMOPkh9EBSpw6P8QfJvJJLArhZBXtoyx2LoUFSXy7boYbZC
0aPTvEG5Bui02zgg6Y7CqpbwreWXUJ/uMT4OMHKSJs6goDw59OVuI+xDePlMd55jMdXmjpwM1vQL
C0WbewV2I20SvjvD+JU7o7YjsUMY4eQ6TTbtTUdA4/zVCy2ddU+easFr97K5AGWUkw+HhqDnPRI/
nvEL4tKLN+jDHcA0RK2q85tfbIJsRyfiWyMBWHKHTmVhJAHGI9VMIOaU8fQSQGfm0Sgt5qn65F4q
IJFOL9nXTLNY31ziwPGxbdZ4f4+vmCqw8v0NIVmREvvhTuEC8uHUqI+kudgcU+4desdVYDdeD5H5
Ksqac5Nx6QTv2sL9NK4biFNQ0Q2csSFHzWVfn4sWJ+S3kfNOYcAPVE0W7QuEunIzcefhBpjbRw1Z
hdbMZDncvhBK1d+4F7IsCWk6zR0QyDiX/vAamfbB7TVSlfy1HGrpXg6TXvCkgagJf8IJ8bwe/Sa7
RH0YLWwk877GzqIb9MXvw+FpcxSS6ClmaBst0Iz5R7jfDtP9GpkXL3hImGi2+gZXzsc1ii53aV6Z
GeSEFbo0GjzgenDiMS9mANtrx5bOhxv3XoFVYpiFQwMyJHPFny3LnFO7YCqKg+RR/3qqgFEsIt20
izsD2O8M3QXhtmo0JiHeTFgXqps630VOiUIM0q/8hsYLjiosQjF95rOrB9+jlGoY85JWTTVrdgN6
7HHa/rrEf3FmnomillB6lzE//7mqWwcEbzezgU7LPsdJuUTWtoueF9YyJm3vpglyqAo5Obq3mpGt
n7bGDsjjf7+PMzKCIw2rzELR+IjsjdD+ATV0jOTCMfPv/dBfXdYYBA3i2wdNZPRxxjM5KhvA9QYI
+v4y40CQlhfp+zyiqafjtizL3Y5/N9YOIzMxn3LBAyGaSGBIjKxNEunhfJ+B43wSzrnRNLDBZwzu
P6fJ9JrYLR0m/+XzDPNYdNugqALmUHovvPng1jrRh819j92mMbg1VqnQDg8C40IZ0Y4rxIVElEd4
sRTIUxwkExKCN24b1X64AifvDzJsCwYeZJ01cLsDTrrAdbDq5pw8Ov+fQYWZdED+xwPwUiyA/Czk
SrWdCKLaFaHIhHnAlfo/Ydcw2DjUo99Bn0kpnlO2gOvotK2N7qnOBCwv2BFtPTKCZKODtrIoC0+X
keQOl9N1phJ+tHhuRQLxBzRPmVmXrwxdmWQEaLKcoEAj4lHympii/whMBg0nNmzLPsYVkTOXXwSz
Owo8h0bCfIGDgfq2P/x3tyvaVMyiTXYYe4yrKcRN+SDz5zjn4MfDzVqgXAD6B87I33xCTQ7Nh+yG
/3+dxNSrDyMs1G/zKBTazWANYODRPr0InrIl0cV6jKrS9j4DctWAXo+4Z3UTaYla2QzpFMmbNGe/
z/pCaLreB9cLSy0s8lyLcdkRSFNJSOaEmNelJrPfHZfPf0m2+PsbgXJA+U3CQrwMNxBihnOq3vKf
cx8jCZNhqB7/2JThIIrBWCFFBl1bo110KZu3ho/z2pQqldESlF2upy/sbv5VXsbh2ZpxVE0w6cZu
MWd4kBrBH1l9fhaulmpIu3TV7m5foU/cX3sAcaP52NmBD/p/MZZlYN3XWUDw9r8qAoFnnEoLDHl0
0esU0sLziNqliqnrkjlQQ2NfEYbbVepsNYITkVjWusFS7f3Z1YMtzQETMVluns828QoAuzHtV6vk
YCdV7Pd1gl/cX0QOS+r/el4Llu7LdrQVP614HU0F8ZnwM05js+4FVDlgI88XvD5wgNnh1tS3ZBfH
gk/uHOFAuJHZ7lYq21U64EWREL0sLIOp5NhedmLA3o4e22jC0FjiOiAmIM+rb/SHh/52QkBY9iQ8
E2EDkofKOkQ1M6YglV13PW/kqGFpaAdnQ50jDImasEctWIPgNq48PnJ7gx2H3DZEmzcatJmXJnAY
jLt/lcabVdIpZH6nX7DAzOkl+ZrHxC1dfRRqR7GqoI+1cMym+RHXGrcJeB4WpLW4y3aFzfdJs8B0
0JNNUQ80kYrweJDsJdaCld0ec1JNoDFZex+fBhIwph/T0VD6GM2ecW8a6RFzUgoLNcNq3mdEe7fS
irjmd6v/z32yBrT04UobwWPQ67qSj4Y3xPH1PiJ4TcbX2LH8fyUeSj76RWYcx+QyTqbYhjRl/Pj2
29FhzafqllbrnI5exZGuuBzIQqJ0jWvTPqROYnsuMAku3PVNxN7H1Q7WEhjNeTlSjehhnst5/SLf
jLDOc/cIbsKUqDEq1md+plAy9k+A0I9sb/CyggeUwsFAC9m1Q6baYHG1bSYL7osKLBDM1ywHpjCy
z2uObAw6bFcfj2keLZQigf7At3JSdVioohPwzuGAWfuyKrsSjiL8WWwIrr7L60JZFagBeqr/TwJu
rI/Dn3aDClxdLDH6tGVnMqEUnhlpUSRwjqVBzSYrJSm9ii+MqLDPxzyWnPUehCWDiRT3UHv7g/4W
WsYit4pysrwgXhrLazAn8u0hvW9BD7csZgugGiChOkYqKuayVf7aU97lYGjC+EIm34HfAdSgq8ei
x/o/NfxF7gtnnY7gyJFQ96mMp8sOku9TRHoBsa/YMpiEZ+5MnJo1FSaqBE5FLfIALfmKeUlG5mMm
EyQ36aV87eJv/luVTcHehiwQptWmtFJk7bsvkPo8ZvYOHHQQ0bZ0572QJMBrf0rNL6Qksl17EnQr
FSRXBJlrRs/3MtJUwo0evJyM8usAp8Hvr/ByVe98zM8IGjy5SqA1orbn3KT3yykFZVGKnN2FYQkN
OSwJ3dtpg7QjZwQZ/8QsMYmgNfnK9rDfN0ZawHSZUmeMVY9g05MOMSiJqCIXUO0cdU/2MSdIy8+h
6DSSWoOXDYdC/9fJzHx6u0ttk5DpB39aYCx0TYlWBK2nRMqqeJTTVTl8uf8MOfdTSWmXkoMGwlTu
5xBgncJMgmuAsihAFq9+UEKvB6rXOJ3h/kaWMAu6q0gjEfbzwnKsysXs/8Ych/02JqpxiIcxm5HQ
ZH7/+pGY4K/lOnEvtGdqhHDpuF8lzSwpJcWj2a95AvX/WDqI/2Ky2jqH202DNBwuLnZNcT2tVeLN
aebzMhipIIJFy4Kc0VGN415rFG8sQCmsKfhm34WB0DTrqol6qUa0+tvcsn8fPZiUFuYRcy8FPM1o
8HDca+deoKiPNbAuJJbujnaqZWDHDdhxHQi/VvFdl26A8UFox3JgVXExZmM43e+GLJ0+ATqQW+QB
iqc2Dw2U9TB2Jxgq81xdpNeomNcwxhsdHPum+mp/ves/HUkIjKK7COblIV7vZWaToYhjc0QOGCtH
a9KXnIx2vwcZXpgHXIT3ldGRyJhwPRvElSczK+mtLZH0niIGozGZh7I/dMXbOeXfC1fSBP+fhj5f
CYf+RfcIk+LnD/k3J9Y6yTPsF9JPvIj9fkZPVvWDyPmKkguJsUDOUwQat+8Gy7RdTp7F3LI4KazS
1hQs5aM5HphJqoad9ZGCPi8zQk/1fJhzRrqJFxknTVjo8mh/XfvT9J/0UTC4h7Uv+HfUesKzdTIJ
YVY+LOu+rlA2LwDmdDFPTr74R5/QLN+SNNvsRyrLTaDz+DFlD/iW8NCiY9HgMJ5BpBI6BevTsoAJ
YVWWka9GZNbDayl0ESKS/hZJs16SxdMuvoBs1v961vKhPzE2a53ncrPQRmk0CeMl69LqzB9OYgcL
AuE/8Osy5awiLDmFmEMQrlouMol3CURv9vucsKfR68RQpqNzKdKk0ggosMuABHfN47VbCK+Uxfj+
p1HtgTztgswz41nyIifn7YzzL0vluFPolHO0K3qkDBL/QMo5vJwqXFEVom0/sKDbGev5SeIqyLqE
ufQttkxdlQowGvYDsT8oOH7YEaCbDUXtIXqEUQip+xPXT8OncS1DXNK0BXbe+ckNAZGCNHOeW3OE
alZTxKVr1giyyatTDBnwwEClGshTwI1LobacPFYpr085gOOMcWAHeAQRqVVWsDVjoSP4lwcBcNSm
WZUpWwHBXMLd3TYRN9YWH3Rp+kz41xKSyT9XI+KBFCHbfUCI1s5SKRFVUn+KKVntoRzjAuhyp77B
oNGJtRL1fwVcmbNwpQggRYYh2wyMa9gy2ZibKUegGjn15oVB2Hrpph3q92nZUCC0RCyFTk1VTGM6
YoK36npfgwas87LDHnyUNwSClBkepULp0GhRviQeL02atFCcRlB5CCKx+o68lsv00CLhp2OLk9AS
zmrNXuwhfug1+TNENusieHVBo82lmBTTUQRzgwcrxUrCkqTFnQC4rFjRa8KgbKgn2euVTWv+L3Sn
UEuUglPAQOBdfBVIJ4jjNe7lgkzh4bFmHr+j9eNF0gBbZfmG1NXVrwINvrBUsLBnH8277YZKCltn
bB9qI09ZFQwLST+vXt3ye8b36EfbJq5axWCSoUpZt67T3Zm0ZKpfeXrRfDjaFB0RKfiLtgT/apVn
8apjHcFDCOuI7+luTGSXUsWq4FPVoLHMmPWkAMx9yRhLA/teYl0QMjNXovARJmEPmkuPuQ1hQgQb
Ur36w6TnQ57XBkHfl7PK46YnSJWieYC+ytfGgV8Bz6/BcgO9yhDrTw5OrgRY9DHp8ayvLIZSZ/F1
l0mVLtoQJXu/gIFAUQq7vmwixILxZKdCBKK+KaZF5m+b+NfmitplyI4XfiiHsm54RsSqPZ23Q7nx
CNKi0qpS6sgXJNxTJTfRTqhAHUUwv5I5+3qIzoFEuD2OvTcUo2XxlRJeo5j/JyIMWyPMiAgHyAk4
Fz3PAudEIZrBdWvM4AmQNaPGPunvq1G52u08bfkayxQfo/kUjZXCad6HGoHHCLArCrXsk1Vp1wUN
oKvaHrsErpOQSnMUn0fw40D7pqRSpQ26L4KPj3j1AUB0B4clBXhar/FgQg0cWswhY8yEqTtfmm/0
HZHSlR0CooHkcS8bpCHNk74IRiqYIHNVNX/g22zec5mScsNkELVZkzcgZjV3dvyCB2968OFEjpqP
E2XA63MADp68YSakvpbLzgZIDkhinn5mgXLsRMXVDPWLz4n5yEqNzxgsVTHivAS/Apbdlelnat5b
jF/0ki2sflo3hN+aLIbumtGcHM7RdCyZLI//RHepTyVOP/1yvCQVkcib8xH/DZZucbL4nuJb7X0e
zlMv+nWNXRTZeA/59O6no66Kk4DZWY99v3V+65Qu376pEos8+FfzMGZWsnRwiZRpJ61VYsAuCTDO
BUeYTaPkrOG3QWzZBTk09oN8YR6beKwJYRFbEICvMl7aBMavBpIuCaSW1ry15AzcjhPgBwMkmgCc
hoE5QuskGfDqQQG+8rKdqgYqow//5LkUua+kWinI3fRCVrZef/sMyzKqLf4aonPeXz5q/WjiAe9M
2IcczgzAVBqWVsBjFu0t6m/RmWe4T2W/9nl5xG6I+gLTmBveJC0Hctb3kk4BLHAyJDctX5/x5PFs
Mwpjm7njmi7Au0bHWmxtFqwYOEpB1BNwDav5GlajCY2HCo0rKKiVXmAXxwq3JcECjVbK8/hQjswM
I4uiLFgbEl6UVY1s5ej0caRh254WIdgywEJENCvHvOW2ck+o8udDrPF5AxAE0S8t9mya5/vO4YdF
ZKhQn/y2NBDhLWI+GcNsUSe+wl6bAqhJpA6UWFT438dFcYCwGxei5C2pB7Ul8OKHKDsSZBrkRo8C
DHuAyki6w1kXTwGBKyRJKrOIZ1aD192dmL9tnSOBL7KOXPcopRBFGIR79M3RsEdXJYYfM3cbLh9y
Lt2TER+odoEN2UFkV/6F7CCww9JcTbua9jOnu4WyuDbuHvibr8+kFEMZQZ3v+pZdQ0JVr/VIWjjN
EsehcC90a9XliYqnkI/Gsub2SN28n7JalJaUyCbZ0gkPIxIdBll3SpBSG+25QN2AqYJXBuEpRvbS
0xi5/iVuzVagPV2q/wRayZ6yWU8WuVB3MFnDMiA9ZMQdrE2qLGXFCxxSB0QYu2v8l4kmfre2k6tP
SRAg8khHwtAx3b95E5hnwBE0+IHh1AVjtbtJII0OkG6sZB/TOe8C5brgxhn1xvwxEJjxxv2Hs/yv
LE6fUVkcxJ9MAXLxHlLglr52GUutvR6pyijChW9zuHMi4+3CqvMOY5NR/XhyWs96q4kQYGPMxtbV
bTkR6SdZex0ANGYQnQVKXlUmksq+NPTN/nN4GRmjezfi4AVwK1zGWd8nQCCGW0b+qKKu1k+FRUV7
xZLHLikZyc2hMMsQCeHHpD2aFsM5KnJsguhwMT8b5HOfozlB2U6pqDoxyxVo01zePwfm2YZ4fI5t
2u6dB3on0sfm4s0fvB01RVzXXznBA8LXL21LZ7DHFU8xoJbbz3+pAbYI/u6erUx+3CSscN5butNR
2Aw7g0fLQ1bBB2KztsV0Rz7TAL8nwKUcAciJvlTcozMOQm5SL9qDiGknlST9VKZ+ZVBoMYtU+AGm
yuXC6MjvH+jUIwKWUzu2/DE+QK6J9k3iL3qvU5pqFq0NBurXzhGmkfY3Yn+Hz9lA3+pqan8rPH4v
aAnjvn+z/PI1GTK2BHdBJBlqNywTfYh3RdzLcfXhZhbs72w5RNtcccbsvx6op0/nMcYHtB+KUg2d
7Fe6jjQ31WR19eSxuavRCXyCFSRIa4Cx0jCCqOQLPxbc99Gvflb2rm/ksmn7SzzPy2fmVgJIVHOZ
bzHryV4QJGHVy1IompHJ7wrVYv8pfKjB5BGF+KeeDmrOO7IMhWje6YNtn2pnx689YL+vWmj3wQGh
VTHcSOX+FyjsnpRMqw7R7B+S/quY17WfWJI/O2RpnnkThgCnTbVaNHLRw+6xize4slCi+OmqwEMk
aAEd7XG7Mg6+7L8UUfDBTlBhg6GlWrH+Il9k5631NkVKrOPMwPdFkJ4REE1tgDHqU/W1ZTWw9IP8
TQ5JgwaUdhqcIOmBNi3lMuc9rboeoZpk5rJH8GrFEpbIsPI0db3sBcOYeaJhs+5PCaY02IKYrrmg
eKy5XYiX4rUYMF5MELTx69I4O77LGVmAXrMoLNrNT6dSVzj4Y8j2+s5Np2MMP7QLB/DWTbOMXUrr
e/wwxnYyEF33HQM7gfUq3CoXXgN++pnGqDmfZ50J3nXtbFmevaC2ZrlilKTltpqFpBxd3yyHy66h
yG2fPk/HkmVurAANe1630NblVNV94bL5RDF2dQ8GF8E0n969yLmRRBHHo9Cric+Q4KpUE4lOCfen
j2T6WI5RuIV8YUkomU5xAjX1JWR49y++u6OFJtLRQD1vhnmqOGMx7pw37AL3/Jbe2BswK3WUbr6d
jt/d0gv1Oy6Ygg3bFrMYJAPXHx+WuJ3mEBc66BYl8BW+3CgSLhGJOH48tbaNNl+TnJPn4RTfzq2i
757y5FEvQDjVvjmeLpKSZSUdYHz8CmxoybsraEAwgNUqH1QdSSt2rXMzhJioNMQq8xzwYdmoyvuK
Ec1Hb9rzXoOxBjXMg1EXJZAGZ603/V3HqwOEJzam4clk3wpUfXpWjDBDJifpwvAptD7hX0YP14ii
g3bcxtuD2TlznY9wnAQszkMEfK1GRvRRL4ExXZU4ZWsCNbGnLn0YmrfOQbgNKs8ZQSmCOtYUx8Pj
hU6StSfTdC6wLFl1RBnrqxrB9DU7dYCKqfI64txJW93yCI+fk1Tq43TFwJhkAwOsYXA7arHaGgas
P5o7TZe6x36M+AOQB/dytyCCeq8stQUgzemihE5PRU4YEPDdEiQpb32FxR7cR1DQ93ZFgS/e8hK7
XHFuRjOnQqFA2dX2RA1mjDYC7e2E4jwaGjCSXmRtNgapb7aoItLvdNlG7VxpB8s08pDTUBUKJLws
ss2QJY/una/iVYK5PogAWDPFBxpR53C1XgoA+lRuypUNEOY3yG1IaseWXwxGRBj4oGp8VWGsWFvd
zk67UNyQGKIkwiDnjaHRbXh3q8iBMOH+mlPPpDrGSRSpG4xH4zEC5Fikcud641sS1tFBo8aKu7Cz
fORfFDnIGg5H5EFFBApPfUi4DerJkGr4nOVN2k3rm6jYNNThTidwHT5wqiQSqVHKbbPZa3wvBt1g
ndnqwGQFn9EKzX0nZHvYovpzU6nZzD04eNOx8CnViaFNzqkImfASMqN0BJodwVmkRsxjaQBwDOOb
ExoOlBGbKPT/pW/U0YYlS9TPJpcrI72p/9rf/Uygp2Mb3Mg3DpxOnODz36legG1cz2NL8gNWOkW4
dLAKI5ckpdbmf/jyoGUSlOSrMbRPslEZDQ6c4ZcXtR9sDZp9rNLcT0ilYVVZ/iNs7dWR0AAt/+Nd
RfHJq6/4Y+B7PcpVhzKThtKaWzfIExg8sRGShYi51M47tDSm4lo5vuElL1OvnlbzUTkiBIjxNbKO
R225wU5jqNBOsfJ1//CEkfDVFJqCeXdiXeqSMfN1Xwp2NFBySaXhsLPxr0QFHlh5fbbTppsAXWq5
BOTMUt0W9bStCWfdjdLnp0SMYy7wePZQuse8B1uNzWcLfSUWbKWze7F04h8/6x8dFzX7WTBfpFBs
c6j+WCsCTrcZijUyg2Z7ULwAmDA4dpB4bZP/3fx+rkCy3f5rRhZYNpMRU9fphbySKlxKndKNAHe2
2W1vXkWd7tlpxM/jnH7c8WFsy6sbzAR52kfeWuumOSnuY6IBea16YoUCkO1Kds+Oh5IFpXaI+WqB
VqAeh71yrCOUvuisrQ4XSbQ3wdkZ+XDLcm7ioZ194j7cTM5fZ4afTLYzJah5C7qrTKQIHt6sFY+G
UFweKckWXOhPoqIsJKKR3B+zHZKsMfsGsmdT+bTI0OxTBAU+ujkW4C65pRLzU69PfBatDUZui5rV
W90xQAgb05TM8br7ulZJpHyr8AkoO42oABaaba/S+AxnN4Z2F/+aJVRe1hBLGANA6LN/k/H4/UaO
wrR19cZ/r6jfW/uC4AS6523gpWrzRWUAHX9WHvKQcuZ9y8dXNiJiG846vxsNwTxQgz85ePLmvViI
MwNtSplSF8f/WhC6N8euPib5Kh5/K011hzIBv8Z7S6uZXw/NEsuyjFN3mOYM69lZB/rnVj4ZgLwf
rlee4C9+cyTTrP4myR3QV9Frgk92l5Va9thn5Wh8gT7khaSD/LwyW8WMhxVADWug6mthuK3vBO2K
B+FbzmX2Y6vhPzwepy2Nw66zFlfsvd7jFsajWEs38iFvl1QMpol4tRvT/wf9tbW0PGhKSg376xkW
Tk7FmidNZrnwvnfvp1BxSuhHG0ClkW8jNtiRTGsQ0zc83B8SfrPXQwUILZzj7ecq24vUYTCGbwCy
AN91EJJ3M1Dxca89CpwV9eHL9vaRu/JGpyyEWgPfrbXIZQ0QgNLVcxaPMMfiawgSIRplmLtrnNQ/
2HEbJE5V6qrQcv1dLXUJzqB0jmDPNWxM5fneHCwu1vNTyx6Wzb7dpxlpQttKlhFEr1J3OHBKZVDt
IcsZ9UcoTgTsqgFhiQKweG6l3bPquXZ7srQGnDEB3esP9Iy/+0E8AC1T+b/MDLr7XaiEGiGh+sk+
WhXFlRPy5xT5z5XsLA717/Tnmsk+q+0pEii6zmNxTfoAnDPD9zT4BLVvmLBMDwkXSXxtJq4WSrLg
Ch9xxf1V6W6fqXBBhUjwGSEO1UmYQO83rThy5mMunS4rboMSJoiMX2WvjVmVFSruOQezFodHPPaJ
ds7IqjgcVO/OkKjdeSFecN72ypCG0vN9fJRtjsoazJIjopssx58bc+3m50fS91MKPZKC6oIa/9zD
pSX/WDYbZknkJEn6AifF08trjVjce1ugVSeZEfp4VhKV4SSWwhCiTcYz+WBDsIpiEm0B1LW6/BIe
5pGyTS3bLCF2QFH7hJUUzfxSHnlwr2v3DZUik+BT9lEtMoebkVVBvatFu4YHAtm9UT3WaGFdS9Mv
xbNhN0t7vw9jt7aM0uHVC33oTkS/NACcfaoJniT7QMsEtgdYxC9yC2PS8kG6a9wldrXI+4AtQt7L
8g171k5+EwVIYDd3lbxoNbz21aV1EDzWlceWpfmEzOM95Upm/eOwJ+my/Vr8rrphOp3eHpX1g6iM
TdbyRt3RJ/5cxncV1IRS2gaYDiq/nOGgh1SUEltTGx+n5K81nneSe8AW5woM/9PlsqEWclZvyQu6
f2gHT0kPHjH13yq3n/xb2V6dtTBsApsw5Hv0eTVskL4Cy/m3k7pY0jaTQiEH1LsGfbf++gCbu1yF
C+tPOoHm17B7sagxVIqvX/TYwDSfvlzd+ve9obBUrRCxL8TVV2fJriKgDIZBosB1Qp5AK/lADFjP
zw4CEc4OotHNbleFYkweLcqIJkguv6Tr+9cTl4BGhsmrOGsiXFojOAX3sE6EV29E3ZeVvDqe6sX5
skNA1U6T2qSe+5mGsUCj0O8HzuMoulJx8LIAm5RY9hvRsfVB9dqYkj+FhQSVCOQezAKFGy6ib3xT
+5M0h7zKOi1k7yD0lghiP6PVUoID7s1x9DUU+OhkRMvZg2l0COt4ih8CmKrK+ia4gDMum2AwCX74
BfA4oridVZhTSyHVaxZvllXq5Vl5V+HZAvT+iWbcwNFF69miISR7m9j/CEQYrLJet/ECalR9qQqP
bi1h2qzXErLBdzhKihTpL+Xin93ywePLQ1vnQsBE0Y3dWnLCtp2ReKhXAJKWE8rnl6iW5dokNFCR
IZz//Ixx67ZPoIP9qE7GZ9Lpm4mUGhLHag0HllU3UaOeTIDM8GlfQG5yXQUWSFpyqAsH0BydlWf2
5yY9VcgBv4PgHrHb4d0pWXukcUxt2kGlU6QpZ4VYVBpFwYZ2RZfrxauTLKuU9Hv0VfHmA84PtP9o
93gfrT0ShZn8tbhUzTJ67VkwnwovB+51OIdCiauJw1bZ0jtXEKlvOFooNUZIOC8gwEs+tkYoSYo/
p3iKhfbBdkagY3vzfluVzyYz4BomEXRJS0P/4CyusbY1r1PliVPgK0W1h29yqHIiR488Wzx3I9zF
mfF6tk8iJVPiHV5Q3+wV69IzNWEmG+eOYmkBmEEHbH0LZkCPh0F8yyRv/ioroO7yCamybXx+qrm4
0qjMzBFjNHr9sfs04qZ6/qTx4LOJnwGhPKVvzx9PBgqkImSFSsEaZ8YwFQhQ4pg2NZXY5om69SZn
gphs6VHQRfRAlyBAjEe9Bugjc5330hBSAvmC++tGuSHwd0q0Ay6KIbNBdfw+gde9VY7f6my0j5xI
MuFT/943YKK4+6qClUttHnVXAA1/g+22qA13JOxNc1CBzvD3NnXLXXp4d9zZpn+51nllruNPnIQX
2d7V7iCYNO1hkXaj/NQcF8prYDgRUjG3hO5DhZqo4zZ3yBNIKdNV9XGBr1TXOHOlRz0kf69jkc3b
BaLWm2go0Xura3RVbMTsdDlJMVU8kW1Xxg4KlU7sZ7CLVKTcFk+akIyawQrLb3CzJ2xIZQ20aTyE
OzuoFvYptdT9dPCw3lyRsvaxAIDw5zfcfbWN6cf5aw3Cfnmm5Mk2Kic9oHG5x81jvBsChm69PZfN
JTFxViMeK08i+8zYJbXU2EZhrr7YhkYEdl4IzuBcZ+Vmn5YkbcVV14Rb2HVrI0q46QeoHh9CCrAv
zJQsdcSRt2CnF40zcwLYdTeF9pndmkhJ9BpYsvEcTY8+iiAiKb2tmDahyhqb2WF94fFAY+OfuBRb
v/Gs+edEGA0tqxeIRmUYmVJwPfsKYSO9E2M+LzMrPMYeOWmm0qTe8UnzqPepIPJM0HzGS3rd0+gZ
dGoYM/z2z5Clk/WGcEhBlm7UpLcrlEo/2PwayIwgaduRzEo9DAtT/fFDmTmX9ak31meykY+tYS3o
LZiBqQD/Qi2xLqGMYQTQe58VSoULh2HI63mtLJz3G1NyLEZ4qBhvOewagH9J+xJpG/LhZNDL6y5q
Rz3osfXKNH/aNLuVMhUqf5gGYap2cQfPGcaLFrc/xJCdjp4Q1xBLvJtkLhWYeqKnAKBQg4zu11ur
Mvlgp26H3efzbrXZxpnCM2ovK8QDNKuUsV+qWEuAwrlqvDT/FKYS/T77q2pWrgxHKT1SfSGKUsYo
DmqV1y5ASxVjjVEwXldKs1gLjTSscqEoiDa9CGTkpB/JOy+rPWuVwrFJbv5/MHxZGgZBWXYPQWXM
w7t6nSXZsSBuYW2wP+rKNl494NUZUAnePdn+EVcA4IVf/FIJJos4Csbs5Eki5X4eyHFuw4wphayw
o3EVeJtTKswKihJG4o4TajXWLdPdTYkksOYDzSSa4S6lsX7zF71atjK/QKx5pTmSgt+hUZ2GaS8G
G8/TjTd4MrvX4+BRW+QFO8NTx3t07OoCnPsK+ihgM0JhGQ0ibv1bN8g53wIe3GUsp0VFLGUIswIs
/4CexLdidzg4D9uguYu63eKnbuz1QSyKSMmiBq2iNpH9NoswruLkUG8PFVDYANf8Ers5qHWT4IA5
PAt/iN3DwLi/tetj3yTNofyTt/jfRWXdWwWZAev+8uz5oeqFOC/88lHokT2rA+0OYhLkdJQg4uFx
kl+Wb8f71OBKXhNy+RHvLg3GrlbZKOx7Rdt7ObH7+Ovh/BdTkj3hFeos2RBN94Ln1fz+C0I6ZQFy
QICCcJLgl8F9xpkuZYm9zTxMSpQNyVtLPqiXhQSZlO9X4kFm0eGkJrC8DSjKo9AubxEiAB1KZtk6
OFKMeOOiQfpAnQPlinlKvcRRsfOQV5IwzeWYECE4UAjVLFJKW5lIXwY0KmrCvRIU6rbY72tbsGQm
i3v/uuBYrKCGgwcoqM2e25//oDQyoOyzwChTJXvi2Ma658C4tYaooLEguorY4XRUMvlBO6+7fvAj
XFXngGEEax5dilF0HYs10QBWWKPu6edEvtF6qtkYSSqajTBBrzC4Hatw5SLUU7a9KGidbFqGdyV3
kOMsI3bemPiL4BUpnnJfVwDYYuiJbYXyv1N2f7NtFGQNMUeyoJPutYlesuXSKDDrODcAFwVVqvM+
d8BiIQvvvNch64vvDc5VkXfNF47YU4SlsZ6B/UAbfUvDEqYsN1EScjIvPrAgDVXG/3MFyslgq7Ov
CKTufj5zxw0oIcZX4lqU6ldF9LsbR+zAkZRvQG7d8Zcsf05QLcSpCHl06BvY9X7TYvyryqKQKBAm
Pt5QnYhbZLD5xMN4qyLljutxE3bYyFnCwoRhVBI7061Xfca+YUO2ZDCNtt5ddMLXRYYYN2uvMURu
HjSboDuduEu2APDQVsqd1nT7CitxjA9Y6ODaDfEw8LF6cC1dgQAo6GumtcWcto5S2m7Nj5eQN7Hm
lcD+s/+G9Y/TKHP9VNNLRFsGpL7W0K/11e+8yXBb1iYfCBlj+73HDJERlkFe5H/jr4idqMUE+CKq
CdDl0yieWSjHK2bzwGUodzIle2ZIPimSwsG9IQ0+BqAmWtMTZiQqo6Y24uscBqg5kRq1Kb3dTdss
z438jWUINPzk6Yi2yyNDSXAiByN/5bZfGMrM1k9TTr9na2NecYtz+eysJL+0dkbRWaekGoaPgE+B
D0CRB73m3FYZ1o6wUUeoO26gmJ34e+A/RMlkZ/+V1VlltfhWG8y5vBOxpzZLU9eKjwE+j6fMrtHQ
eaoOYDkk6eeuAhzPONcMEeHpgci2OBg8BSwPeYPgXos+S254dvT/FwgDhW8k7PnthTWFCHqIjHM6
zIVtL6R1K9CbWQQwfS3isuTk5Lfu9jPfBCGcEXO9ldKJ/dnXplThmnYyf25OIn8+mhF+2H8GOa85
725Ye0gY9ly8kriYDjdPOi2Ov+h1vz3ghOpERgzMsp7JwqJeTjeFRK3TX7//l57HbD0g5OokZz2G
LBGaiAR21VkSk4yL11GsAhp1xRJMKxZUFGDpBHw8ZJXPe80b94juoYSUyL9c++evwWW07omcdSBZ
RUQXnkdsgVTeuavKxwUuS+ND8gIlAtLEXqWEY6TTE7pGp00aul3YUAOh8+3fKglrybfe2ClSAish
d3B5zzCFIPiLtdE4mSwz7c5i2im6E6p/l4JpRJzryUl7UQmRqE6W4FitqyqUm35lRPIX67svrhiq
3rFv6Zz5MrFkl8vRv3SEeJvJkUmyKyLOvPB2TAqpV2iMcQK7VJL0MvMnS87SInzQ5DnDZ47OCFPV
KXCfft76Wkq/Cqllj9RbPmCa6GC6sAdxMD8gsH9AKrmQqVNYnIyjUjWjczieNtHA+Dn0DaydEHyL
q0gf+WGHnDguasB/14nWDD4cN31MmdoaDVpkA0s1McyKDBNWibu2/OuwF3sSl1GRlUXen/xC72D7
/AONB+TaPuZ2lCJv783MXKeex3lpEaoHdw4qfQqHrNI+ePrw7ngXRkTnWhfGmozNMK+EmwgHVh3v
QKR67pwQ7DpwmhXzxnwCqVOBAuKyqt/NXO3Zizc2ulUx6acdbIOFijrOjweIW2mOkv5foEU5mGIj
84qe/lAvLiUZkbbKGmS9scbl76MNwqU3TNkObWeTw8XInWBbwk6nOEu5gKcVSHyKm0rUNDv+o9/g
nTUp2Beqj8q2XISZmYLMwnWLqElRwSvNCY53SJJ5z4e7j4Nw9SU6OmLd4cQVyNXMgAw2tjBfnChs
EEpKYt5j5RY/mHJnY6dWHkyPz3IeX2tthVpr4YV4S6EyGO459JY78rqKT9ClFFg9/iVrzDFE9/7S
WIYr//lYPZ20Od/UjitK0cewX0b20I4kNf6fAiZGKNsaaDrjz16UnUmWnGcPtV0NqxyW5mopyPO0
suzQzzKl3vlggKE4nh0usM97sSE+ieVZe9Mw9RviQqtJ4ZQ6Ric/JoN6ayorukMr5Hg719cGnIBs
dqV5KPI9B61vhV8CkDZ9RvI1JAR7KBJYvNK/sca3yxlWxwrilV3hAi2IIfibvd8P92E11mSqZAuY
4cOarvWPYqGBtOCA3AbqmvlLab6h1AOordKQyHDvwy4YofqtqOUwAx6f+rHVf4dncZFD94SNxrCn
PzL65rH/Rxr2MIcu38sxZZNxlFFSbVseMWCXNmTjL2FPMxl2vEMPyqn+EuFykIC0PkbpJJ1GQwru
YvWGTNGpk1IQMemDkygfUnJZ1oEe8+Pisp81OMh8wa35tAg68/vxPY0qdA5Avh5lJF6Nm+eAcg/P
W3CJnwYZeE5/PLobj7vN9N9QEEs5AaxuEjoHB3ZqD9NtfICh4RdhMFOPjuFp38V8ZgGQI7YpOCba
m1zMgBO6NNDhZ/gglQsaMWLHMqxaAAKr0j8biSQj40fQe+ggzuhvtKP0d1KHmwDaCCAAskXKZ9H5
vnpF3dyiZzrfkgv5qVdDG5Y/RP2ZJzlxYhLbjco8PVlDoeTK4+w9LnkBp2QubBEN6sDwV32FxLYe
P2y/w7eNI1vhgi97GOU9GyPMYhSRYS+5i2IHiJuxGcRKIXp4poeHV1w8daw0PD/XpCmOI0vydsgf
6mig5HE+ev56aG/Xxl0iZW3BQSRtyYCys9B+3jqTanXrO9j75v/KkP085zUKnLsSrRfZlE+BbMei
55PBeHC0NcfY9AXa3bKKpxLvSyvp3lfRrLopgxp7ySR+yZ5qgGF3a5HuNb4La/O21rtfs8xrZ7Az
it2Eo+KkG9tjy4lJY3vNWRQuAEMk3262T8FtQi/KnPVEBoVUI7T6S+uSBCekiTEsbCeF6upuTBne
GkUXiVWqq0JazeQJ49jOzHruVmHbKmS4cx/hZuqtrub23WsFHGiCy2GNIVQgOOSfLARSik3g5yfs
2q9sgUyJL+cStlCcPeHg48EKeG69fqQV9mIIiWvaGoFeQ9gwCaXmvWnNu++dQCJlFnx/4Cb/i4UI
XGnvnzSKfSmY/mwemgc0FKm1oGtxYplXCquLhT/5GbPXWS9AXsbekNkM+crmMO7ff2cEUEUb9EOH
vBwnAzapq9dDvhaxA6+qKeD8ffMh1P3z9IufMn2G0sd6CWjzq/BvYH9J9TGcrzC71u/dZ7fHE9mK
e/NRG8rDSMbb7FDDiQdbSaUgDDUrzD9oHguHPOh7mXoaJJlxg8K/xvWrPyA0qdhcE8T4I3Y+rSPj
kfJZhTIuWvx+0yUKJcuXBMR43XbDHO6zPMR8R1bpWKtmOu1x+6srouMu9b1+9UglhG9NOKEWUL7m
c4+AeQvrLOiOHnrKbB76faf6SNW1PDwy258e6A2tvtPEVLncV1eLqeRfRqvJpXDBteFqs6xbu1r0
0OhNY5JWhf7h2QY0v0Pb4xLkfWuOKFXfiRK8lpLit/tUSI7Pl4agu3A/BPaUYc464f2v3S2NHNEQ
nQkS4dx/xaJ/SBX7CUSR1En46TgiDH1jKJo+6SRJjG30KYCpUprdZYegpEzpVdGJVyilF5WB87cT
W+Klslgx7JIT86DIxMqlRL6O367gyiltEcEliryqJ+/WmQI2WmkW5txy7PxFZt9BZDQDXEUQ+wvn
C8OkaIUM39qCX0EsKLBnobNXYnmbIGsXPYVdelADDKGocxZhNwDJcMRcfCupfKlKf0UEPdOI9mKB
9vm/G4JgPz2PjwAxnUNFaLA0LYzYh869N2Y7dMjbRfQeRCPv/fdtZz7b0JGP4RJxXrgwBo+8t05N
HAaynX1P2K8GGrRpzQhTbS6rH/tdlcbEbbikgKwT+Qefych78uNArqCPJraKXr71rfdFJ/F0OTZl
b7XsK+beT6akinKSP4G87zgIWC6tHH01K4ykVjAZfulPvmGh/eKgSZXAXxC4E7/VSLMd5TkMCzix
g99njWQ+iUEp04f123YW+v2S/09y3AloLnWrVMjW6qWzGHJnTzpaQnqtiz1fHCXelRBjF6JKyjPd
2Hs1E41b3EB3wGLzJ0DmKDLRq1lupsHHqgmw7NS8vOLiXgpp42jWiYRnFr54IU+DT33CFsjzjD7q
QrLw0yaG/OHBjaOJPsf32OznuSiL/R56ke2eHM83zNlbEZ5xs+KnCdkB/YrTfQslU/lOmrZHfbeo
3iw0KNl+ylp9beld0Gti0fBbectt5erNRSKBr+xP/UekWS690LrORrIcAz8K3wkC+HB7q6QowJrX
Vb8MYyvQ18kGVIe7FM/4/iQyA/vGtX1UzVx1u1+tZj8+39zT8npqz/ceNpxz/bBq99Pcw0LeV9Av
P7T18h84tBSGKnx1iA7zWdJftwoDvPnCo6jCnGHyyJyTr+XOJsXRVaa8SxtpQEXFn/7paviRo1Ws
KEnc1HtZ9b7yepV5jLos23jrKOIWvtm0lepeyoWqP2SVjq3nGcCx2hlFIR5p/eqoeB3i3R50WaBD
jZCPyq6o/lcfi/1bpeUpjqoVn3TlBavb6fdKcx32RovGIFW2yqQ/S8mPirbTMYU3q48+MDTtfxz7
CHscp0IPUyeb/Q3qTS0mecYdC2qpfhrS0qFYlRa9Npd0XqsrRdSkPQnsXMy8PyO9EKMdNvnoLEk3
ofoFiBSyKAN4dEgFf4DBDqUCuGp5g6tuQofpyzGwkP0Jg4Gfk35AtjKTK5GKE2r9j7awTKtmZads
14tB26VJDtqAdyk98bEv+Z5iTt4QON/FfpglKmxdxg4kNbFgql5nGW6wGPGurYzX1hVzlLjAoiLM
Sx9UY9H5vehwloAwNMGYAnBZkX9z6i/bgYyJHJGUbpJiF3K68lZ+hW6lnUY4UtR6/0XjCXPx86ie
0dvrYyLJxowIwgoKmo1tGObKr9CI6bJod0QOj55xdJsSGT4NB1cujDyy9k3dHgbbsn2qtjM9rQ6I
hDx3/ZFrF/oT5PPsOsWn4rCste0ZEhFrZMfraQ1suJ5rrFv2hG3+68e1OWgTsicO9dMKku8UW7Wd
s+KPrzcHu1VnXJonaI0gz5c+80z0LQ6llireHGUmaiSo5YI75UYTB6wcRYYtjYFJh2VdV/6ELZTc
5xFaNfn3Qq7XYsZQqUVdT/+Du+iiauT6jCnZSs1fU62MBE04UopDd0FqzKKczGkQkR9Z0IZ8LFP9
HGNSEKSngSUInB3ybWTxwghCbZoPVG7+bhO/Q0JCx8MrUm6aexFmNdo8/KRXCOOUu+nz1U4YTlBy
MRH8EU/vS8dSqMPQ1txmBch3EbtG370Lhpi6TTg33cEvOjVDMNow1DdQ4miccMYGumygXE4E30+K
J1So+iJluDBZnCWD8FjeB5SDiz3kQAV9utKU4dfBr/LKrLks8/l/cLcSr4HgAfdSoZAMW5wfIxsF
6qIHgaR8PfGO3vHuwp4e2FnxGFIC00oObJ+b3Y3pv9fYMi7e4rh2wHyeF8QRd4QtBA7IZFoaOceX
WjyFyY5dV79bCm4SO/sFVu6ma6haReSJrTjqi8VViTz1EbESU/+ew8CT73/wCs/l0kiuvD3KwcDQ
i7l7J/5gnOViOuUK1YxG2+LH1Dg9dFTZ8vA8/2bnyzR/0UmT1P67Jgzn34aXNCQw0wl1kukl4ip5
j25lmpqkx4oWcF12revL6aojr0CHzvD30tZdHXGm0UH6mjSoKqdYDWYR2znwHSFbY2lXZa7aCxOK
S+b691cXqtYLaNCfbSeWdm2ehU1lAvkR5Qd7/uN1A/5vYj/tRB+iAzs/rn+DUmhT6oQg7w81Vb8W
79g+6+uv24SpG9Lfeup9IvFnZAKSI0RaIVg0L1udDA6ghbCBmCK4MiQKbY+SHoNIuNDjao3jeK3m
5MWA3vAhtVcEUEkuyvRhtHmdOSKGfD9nXrzSoNMVYMa7axFt4p+E7ju+PbIw2DVrC6TEXV/HAbOS
8VbkKl5rLM7mY+nF5j/TAaT5TbmgSUK0xui/wJeN2vf11pj7Mgb6yZND7JDpsdyiNoIBwyE4Js8r
gGaNDXs+Gq265bwc1GYZ6HOzHp7rPD22AoRx5S7HCbVAXsqrcMVLXX5lkwnyArotb/WkBfuxMPbi
+DnIGijVW8SCW++leEXde9bHYGK1osUi8z2PiPmLJKFfmF22ZTtFda76u9QCb4tpS73OiU/eA63E
bIrq0Y8mEc5F9vuijo4cWpM3PYIcSk0IYpKIo7ci2svuxJIbEBOraD6M7VnX7BPnTEsUnfbYf+5V
Bo7XDG8nXQNvstcZ6QtqTQhANBV7dxLam02XzVRwsbmeWh6MaBlGFLYok9LS+Ko5oIJjIdH++YDu
wnVG17/4a0N6650lnS1gk7OnaXXMV4VOmk6d/G1Ffk7Y00DJpBlJNJOwPQrwAmVoXUNt5jiZZv43
n9HY1W1vJgbRLYtUZs+oMkMd5TMsm5jdn8d8tha1dlUkyFmCGfk3ACi+b088AxzNf63JD+W7Ul3O
0PZIKQr2PLU3TCMNg8lva5GpaQaajeaQMlwGu0i31g7e91t2n2cY32PnatBua+ooa72ZNEHBf/BP
KBd2ZQRjIImKi9BC4KGsMpfWUmyTAlUXCOIhzgfHw7pejtLDYFROq6ICTf+rpFwqPNYKDni4JAc1
nT2CZ+4BoNLHBF7KdNysvwWIgIGR7lA6A0daghXX3FWbO0WsGwIJoQj85C18c+s3D+vIqnFtl04Q
G/UBOWJH9iWBLxicyUh7tKhkaA6rjvOZYsxpLPwPPoBT7E614XbA54vDXmBZLI9O+fWCN2PTZSRL
+pReAth59sJvlfzBTZ7DuEbx75SWj22lK0fFUgH+u7bvBcfgGFuDRHqc30q/Y3jeMefE5YpmCZLQ
qfGeyULlji4dwdo0Zke9dYdHtkYIMCUqEblPjNKDoHZ2VTorkeK4SAw0YslaBmChWjelD4ANIgzO
k4eyzY0PBEobjR0M/ETNurvpLUB93VbeS7rBmdMtayl8Sk3fwS33ReALH3REIVBGV6ZP35QW9/SP
aCxPVbwm3SSZdmrdAXOljBMhXozbn7SFlsX6Cv9lEPIpgoqhNmQO/vJMWhNWz1GHUiVTequL4Ub3
T+d6X01JV8V3fsz03bR63slELMiGCrd2J2yyjISc/GNRYgITvtqmoNjBmNFk23Dn0acw1XUwSGbA
pcPryl11VzYN5U8sMSsDJHxQms1gKA/yEH9NKh8JZxI2n/t53nPsIAfGip21qV+DOeirim+zuXCm
2qOOhKAfIXcLdoynE/WhrUPT5xvzsPVvJvK1qlqsyvvcm4CmaWuitGZra9sv0FAReI/t7OKqs9Os
aZYb8okzwr3RH/ocOhxRTfylBRKZk73irzzCMvAJHAh+Y9GbLxZEZmL4K5kIFiKAW0Q7TztZ4ymJ
ynigYC2CeJyNTYjc+yi5PB4DguoKCOTgLk/YyIakxHhr1UMlOEMbsLgQVurl3zprkgMnJ8x57Yoi
sdXroMJ7URSDDuN37wjoa3ybvETXWEjMCqgIyxNQV2Q6VR0WEnW42KTwdXIGCdwFyBMrlBI97aBo
ZbGePG6PxHLlY2flAGT9GMYfYRf5w38FehXIjdv444zIJmmKLRy5ACruIVxqmYceg7XQ2p7PtS8/
7HWLgdtJTH/uJR4NdrG2CoISWN1ikigRbyB45rtdlTO0iMMvlVKVzUh5XXM8kGMbVUGS3aJ1JRZ8
DcaOww/fkFqh/uWMr4I/DwkhtAlmOn+j/U3CkNCU4bF0ILF5rAm0+lP1ia8BssQghzUbyzAEFrZ0
o9C7lYXz7gjjiqKyEbQXb6nqfM//2RKrRBQ2/BxprNUfU4PmjubtJMJKE875e5LiEZf663/6rNKz
IE/oP9Tfjt7W8IUC8fPbSIeDprxUFryXrFYNVPxhoQ1Yx/HBnW8hNj+h357+nEPyZDy+PHmaSDkF
fnB7mYYlQCQ+Gny265DssaMnTvGOMoH1wjapuUueHVvquAFPu+dfpZXEa+n8umcAQx1zRfZLSMhF
kaLiclQ7QB5fu2D0Sj/OdQgIWTCpdM+wxQsb7NMy8n4Ew6VmkhjgxL35pFtMQ5wA0GmcIxhLnbP/
wipztMLPck2iLFLyD8/13uSRW1/BD42Rt36ohx1mTmRthYmhrDKpNWPEoqC3OnbZM/ltXq0Hk7/V
ISyabIO6cl211S9hRj7+7MWWDmkikkL1WhkRrdAJNhWDd7ZgwlN/HIcL39jvQbsPlAPjF7PGVu1M
03LAP28QsEebiIT5GJ87Ksp0Zj8FU5x63kngIPGbdsrfL/4nYvhcNSR3+gGg19ZbRVZde96Z4Lnn
5BGN3A1jh1QCwcURJMeDbpG8Ks/8VcxoljaD68ra2i7lcGFOdrbd6Yu/wNiqt+sJGckiWc4tEv70
wGkvzN79s9ezyouHlcr7rEijT8TIo3Gzm4EG3rFSXYR3qUdfB5dtlKLVEnhf/CrgSL/m76sLjg/W
79ZqqyyNJYrT4vljRYaG6NAAe7Xu5FhSXN/lYlXgH2c/AeGb1Y6NJUf2gQz2XzZxOd/20a0EsImN
5K0Pr5grbecuEGswMzeoZ20u40VCHAWsKVS4WkvbwKuQH4UUVV6y6H5uGIhXbBcM7OoPfqD1pFF+
yeWVQKUOg7V0thwJ2zMyCbiRfbmpSrddqwuHdSkzSqwBHDNzOluc8O9S/Htsi34O3wl6cQJ5a4Xn
sTgLq+EsJSGTmmLFhp8phpnB198oRQo297S8NYaWAC5Oh5lQHCnKorsvQhiK/SjCLF63/tMcuQTr
TCg26SEGpGUvyP36Nrs92WgqqHlSXNxCPpbHAMNPAo3l+L6ehl5VzEhqbkHwsBrTpbLjSGMkT5g8
YbCqx3f9gNvghRNAmtTijqgpAigJYiPZcrM6saCacMWEOjzDwKiwypUqnBmYIeewo6/KYLXDIbL9
qmqemRdN+YTxvh6D361Q72bco6k3nmOtElg8uMRQQV4nTQfGNcN+sl4+7IHsHWGXbX4fcfVg27NX
c5xKVMCnf+uk7GNWLRJmiXlxk0/LKKUeT7XdStI5REHqOkag5/RYn7qMBRj9YrhZfSkh2d4zgAig
Q2ZXtAOImrTKei4gqa8RwBXB1/i1hUxo6xMjc+IYi3WlroRD7Bf69z9fZWIzXDD6aSfkDDH/SY16
muGdL5MUY5pWut0w4Ao3cq+zkViZxtwhPTJc329kvUBpEOakFq7U2O64F7CfWKeW7XmdVF/ppz1G
tdaoWxWH7XdFNZdoRxN3i5zAhNVAzKZYJjRmJD8Qx3H3KrnL2w81egTtMucYBNuBjwKI6oRupgok
pscplkvAl3Rp7Bk0wLfBsRwTxfaWE6tYEQHN6e+CjJF45FNqEsDAi+cm8yZDkqlpj8Qutxn8CpqV
grXbwMMz6RleohEp0MvBUbqXcCR9kCR+f8qVTa87Q3m87HxPYh8DmPS1baFB8fskt5IGhkw6H+bi
PJoM46YuPPbxhuUjejJXdk3l2w/9NPl/enauG5fXHEG0hEyr+Kk1m/WDmD2ijlz+2/VJEq9svG1n
w2xu4N8Cs0WR360NGY+QZmK1EOX8hyQ7dqYlBewaqgFCTj6wCOLgyB4/3QwvUa//v2dypQgT/4Ax
7xHnBhqDVXmmuGlaVGL7Ju6DWV5QLSx2ArmdV9fRufXTEbPiFlIHsULb+Rubjb1sYMNhMSLHWYnX
ki/UqY6y7DxSQnKjemQ/a6FafBxxN9hMCFmc/laHaOdoLGuCZnDe/kkNueWLVP/yM89HNePwi+Y0
ia9fnk5SLvA28g4rrPxSIVOR6bY10fqWKeBp1Uih6j8fVbAIQNCHevBI9CX3RlnWy5ClbvVJqVU5
ed/kaSGnYC0Lt1NPdAe3HaYqxO4oeyALN48yeaWJwlG0UdFnyY99GITDhPmH+nXVA9nhxcKNXOUW
PaAlks8hBllPTt2pczN1pXDElxWmd6GFCTK3bqDoE+yBJ72zQEaf11wThb/QrnWob21wM90W7erl
xNs8bzLbvl0bjsF59zi3RRgLN0a4kvyPHNHLTNKpen1rbqe3nceJX0QEmEfUtdog+rnM1Aq1fW4C
NvaOKXBiR+mHPlhX9eNCHEzTtKPmdgmjx2dTM1na1rVhL8MRCGsBoUrwBqbmNRMAyKKiYx2R1TTI
LRiF6HEIeQFnsxIIHRZHJef8bTZhHZd3SP6WFmgycgO/w2nP+uW9I4idGIbWPRxHQnVHIQTZknQi
wm0L8K0UBf0aDtVWGCxzUt7PdwrCxKPd5T4Elmgq+ieYxzhlX8X77WqbNVNo6saIT6mZ6dfHRRXO
cSO3xj6TJff6jggdCfN7PIkXXSCczBJhhLpS+AYcj1sqQuNgVRhH1WsEdoNIIeDyNHUiM/5GPlmr
rszUT1Y/w+JtYh90AGSPAMPXa+xdo4/xuuviAaVqSxocqivItZQhss+ajoadOCcEhxv6bSPfUc1l
MHtVQ8N9c+d2p7THUaaD60fppk0Ln2jZ7tz/mPkM27/waQkQGl5bXRVFzWmgd4vktYQc10JvJB14
JIdKm9xPtHAEeovGFX7yUmBfFJLYwCyotnW/wGV974/BjFbj9z/UloRQ9Za4Uc07uKIR6E30npCO
nk7js0X/xhWIZSytj3WNhcSPQ/KFQA8oG2r7xmVXNsCKjp8P6yjkZlqfxbSSgHfVC5s6pStdnEB7
McHM16U0124P6RsD5NvS+F8xiBrGrFS3/rgdzSmRCG1g6/IL0E72TMOJ7DGYqy0kCbKfGRMQXqTI
kMTAtZl1r+Y5HRQRNW5FhICr1nJqajOsDOkQj3vbGC3W11KsuH3soc86okqd9BXtm2yIvZJDwcPV
jr4UJwUiO+Qj/dkgvdJzIq2KMkQPi2jhWaGT7MLv3ZENqhVoobAZelsVgYj6YadOLVZeXDSNTt6j
zzGVPLJ6o5kYJZKIKdFgM5ilDUfXYnSeK6HWx4LxQpwmrRmQ+KZcODVuerEHZO9DNBYJ2sBhC6hN
kW1+84Fu+3XXWF7c4NpmKV3xerUY4CzbqGxlh8pSUy1G5PuwU0TeLeKq2f1Uel9mNJeFn1S0C1zX
kcubLU3J/GLr7IiB6M7lvFgd6T+MJwze74RRRq0D0IMvJMOyfozPYh9vhi+zQ4DyyDa8hrwlNvZv
ZtBNWM3gvG9B1XDXKHZYp7kYWqWgyfa6m0Rc+gytWAjGtyE8/nfvs+aILyY62BatJeh7rNKZ6+Dl
paB9h0S1WLG/NWoierkr5RMTAQqTmnX3EJu0PbWcSISfupBUbKkhH6uEQVX7jjbhmZhpRSoX7yWf
l/Levc6sZQpM21Jt5QoNn+Wsi4ffAs4X83uKkNGLjgSai9V0kmbicfMXelgaL99K1+fMf4QdhyFj
gYtQwW5zSGoGhOTHznRpiteaXAfSXYI/Ui6/DbakfcvvWTxCIWru+hSmgT0lknb3zmnVXBI5GMKJ
k7GUSGVMYWGdwnhBbxmPq9i+72/lTksSnHhKnjF3MQULgMg5Ad5gk2FhIz1boj5IAc51wmAnOd4v
mEpF68LCiPOrpiT0LBpjUCGV5wSGjzSLHta5lpoZ+VUGt2n+loKywoXp6z532lS85FhKGo7xClOh
QCqjoy8lY0S4NybilDYcIBkzJ9qITcabCeAC3+zaFWFhOVFom5epHCy34/sJlqqU7IPYnNdd/+Q0
F3kQGSIvIz6eGAH8xcUUn66Oe0Liw3N1ql+aYMKNNtVlVVNniiaLIOiUKifeFU8HXvaaugdT4Ila
oTxuom6bxxv9hA3S4O1OsUlGzqokqIpB9UjJqzBdNmDOoeM2K8FzjmFdjDyyXlrxJ8GPUzbQwVG0
AaCOIz/2S+mGj+1pz1T4YYHRm/JIDD0Xso1+DOMQlXD0zLTzbIerKqRYgi9jcSIH1xyeg1dlgppP
6gimop4iBMBOfu9j/LD5EFb9Q4+4UXOoXHscoQnsx0qLSmfsjv0EPgZZ6wgYiPPSyQ1vL6H/uwcf
NpZ6JDvwt1I6zz3Wy4T9l6aparxRVZ2BsAoXKjnD9DN7bSKw9SKWYH4kMHVUpdNTdvxoeGjFANv9
zng/VE5+uDT60HALg4h0Wwr8zsiiUNWiMWQTHB3K1rN+HL/+qDKZKst4GoOYCOsynAEICdw1mn0c
Y+TDLCaqVE1ruQGWd9cCY+Yd/FUvHUZ4TneOm50dtwSQeh7ATI3zODQyGmwCidGpbvB0TKOgBY3f
pGU9i/K/yJXGwFeSysB4nd7i1gMKp9cQNndu5UKXN908imDfwUEIHynq/v5yBmzi3ry8HcNf1UGm
9uJCU6KpWeIYL8wdg9JMcF1xSOU/avNp3cid8Y5Ktgji5O+IBzhqYtPLIKig9O30BfCpStrlgUB9
g5FP9n6+K4HvBAQrdDkdjpkPb3QmhghGwGT9o6WSOAadhlrQzlTy+otZedhHuoHuzIUsUIZj8DwX
dDuYXfte6S+DbRgG57sm647IoOqNUhLrSr+zvO3uieZrk4MKhE+A135bUy96JNTdwD7phJRdRQb+
Efi4rQ1r7rVaUqO5NFKLfZa49cS02KASWphWO22dEkXOuwH8u+4viGcowWzkIaVLzYs+8ub99+J+
LfS9ERv4NtW6HZezZzlPDeYnXLx9FaxRvLg38okJbXxm/iUmA6cMVE2IV9U40wIdqqVYNFH7T2iN
e4HNZKffuZoypc6pWSfQF7cJFKisjMjcGKVCrL8LaOWlvipEh1VWlQqK1vGcf96ylwhxYl4aCAxW
6M52tZoTz3rMrZpUBCmbbUgswkS8UvXLeIfVeRCU/eXMTc3LwQJqQZf8ve9lpknMytk3e21ZHgF5
E9NuvvT+D7YZc3L6S0XAZk3qaVlUcmgRxL73ghgIa/U0bfgt9PPTjqws63hUPzrP2O9da3mqdqYs
aA==
`protect end_protected
