../../../../../RTL/axi_controllers.vhd