../../../../../RTL/mult_add_sub.vhd