`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
IMfOuVszrCgH0ngu1ouJoowV6ohQv4V3V1+Gazj1q7/NtU/bt/5hbSkxOIH8UY6CuIrvK1LP8d5G
dzqe6i5Yqg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Rj3sIfrl5jIc8ouK+xGH9+Vmb8iAA598D71SREywIYt2xeXfaqopcekSzKblJJjcwJfZdPL0dLXy
9kZiO2mtmVgdOmBXAe2YtOT2bcKuxpS6fqwlM2G3v1wW7Q3PIYgy1mQXWjyO2jsud8mSIcZlHuWR
5DtyHA6yt3lm38DHV3k=

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
qpkKci/TPEjLiZ9i9notBn0cPPd5yWYioHamDNIDovefkaHtyEsXG9ctqMlttCIlQwTB1rgpsB3N
uxFWsNGrYh2VAwhBSMzkaSEKPC/4zWWRCf23uU1Dm/QCnGSkybfVmlLVd80F0xn8GQCkhGdubqgl
PRwJQoCgttQUmYoIEE0=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
G/QIk8ccKB0XtXQ6fGfHb+EPAkk6gZMzkFTIZflabNi8KZ9oooI4ZgzE6HKi5upjaTOx0Mr9nkQZ
+d2ytByhIiJagHZ07OuS9gpp/bpbXa+8v4rKXSXdl+9wCflZZHkHW3xrVc1RTLpqjqtfZm75tm/5
/TJx36ynWxQO+h9kctxaZd6wweRE+UOPu/xNRSG+6s6N3yb4PAUCs4uRzDlhCRoWcEMXWYU6KnsT
oa8KPuXh2LGaD/U1MQFRYl2Iw05SWdpwmFWX+XalxTIPOVfTyDSb4m9WYtIgNW31H/oLWD4gOQPn
dy3k8qJ2TkA5fgwhFEmkmycIMmFOaUse+mNywQ==

`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
jZ26NORpmZKspxhxy8E3nuWInS2v8SVmkJW7YbNM5w6seYC6djix60+PuZfxYZ7kYFJ/52hCpUm0
nlkFRVUhh5lOsAXwHOUilGtX6crbX95LdjWJpcaakSXkSao64l///V1aogbquQjrFFMwDZae/Itp
GGStYfEAvZZF8v2cuoV7CDCyqdbNflaLJmv8cNY5vmP6WyNlo+r7+YPm1Z/TCSJwjnIdepeTPWy1
kQm3+Xyp30gQq4l15O2XxlnvMSx9hM2Hnkxw3sufl+8Nif2AMcfY+pyhU1SsIVi/GEXBguzhdTXz
FC6SYAJGYxKQf0WBT8hclumJaE4zNictG3XzUw==

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qcEeIzaptklUrXjzLRqVvKspVtzhkAnZvVXPm+n5SiD2fptgVEbzwyjbN0JRRJVziK3Fx6wqypeb
ueCQWnOKML/tC+M1ajDJ22dLNEunTuCLt0abx9vGEyxsoifzV8Dy79WEc6gj5QBZvCssFHNviiJw
pJ35EblO+QKdVSQblS1KBaiPQSTQkiyaxz+/Qd3UeWb3mlDNdNal5m8ORG6qevEbY1xRDWMR5LRC
7pIj8KyBHZoF9fJvBpVW0kgh26pl4BE+Ys5l71OADSKmQsPX5UNqg2O8G3/obQR4JfiUUmRME1ze
wTI84KKJNC46jimrrZOpzLXBHkFeFpiZnfhkJA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 52272)
`protect data_block
Q1YHzuFrv/Sszj+j6NP2B5VGLlt4nUQdevnEehFjO1U+2/dnADZbDOowqDypv9U0cu87laQTUF40
M4v0HKBwwQW3/OaggNERqBpwLYb+tTS4NAWkFBvgNXePc9k5sSKTc/q+5iDDTnEbsh1qUhzaQEdh
5QBOyxNdc9pAnjXlxG2Kl7bnYHIcVwlOfH9ymRkBHjVn5NyZz8rP9h5DBof6Wdis+T7rgD3BrN16
NqcfMuZ0Q69taRvNbCxRsY1mlHL/sI6QjT8KC4fX680mg1WQO+UrmRqvBOhcs5rQeiajliwsPORV
zRnpO3SC0qUZwAT93fbVx5pzXZeGmIXfFgOR/ZmvQWuB1PjfW2Q8KRkgd57tYbDXFGVshVBSVh22
bEm3NM9pBy1fsgBs0sCtpm0ei4wcEP0FsB+KYTTWGrSBmJHvDef4zbp7zqSaGluLwT3h+5d6y6NY
+hRHyoF6s+XF/+an7CO5SI7UgByYWLI9vtWWZb7WHm5YwMxUSCLOyQPq+iBXLIMoEDMkijYLt77D
n9Oqh78bsyp0obbVS+UqxDGubDdfRCgtTQwAjRnNcunrIlttdL817u/fbEwbtsUU7ml6Kg8/rkhJ
+DnB3r7GDEX+NmWjr7A6PPmp9Ibb7BC4hITVZaggdKw4Tw9BVC8b3yqdeQLChLAcFSxjMZXSehKC
LgPONnEuryigf5hvs2rAyUZv9Zctf8ZQe+ShCxWfeWyh34BOIuAOXI1zsN9mqMrXzwbCQCbJdn7V
+o20Kyt7xLkP01AJ6FpEki/NVjXOjqyMS2Lzr6UEvB0r6OzIJ4KIsNi89RKttgGNvUDjMLxU8fKr
KjMK9QrDbk6YjQwmRiVOSYedd+wnbA9sEAyj9QXhf/qVcAH2z703llL5mpci+C3NaU5TQuHDbJwi
fN9XaJy1GeLN/hvJheueqCVT96DFayDwtVfWeFTw7ehrbCzxKfzds7PtTcYiUneTdwr6NN6CiwrB
OOtUvy8wKAxcfe58+3/ML5YPmPuKzZ6el51MWnAhjh7z6XrLr95ghqS+j5MriASXvT2eJg8UyH/n
nFCE0ZBnMNq+neE62nztSlZgajoPj95TnZDr1mPzOsnYW/NLxMYQ2T1rms3ZKvQVKiKB8/U+icBL
9CAM1jDRv8NPM6XGM+dkzsSC/7719bTm/JeC6gpB0SLfCpqVKhMBNGLiJay/vK0saqWGvF+q1Ozj
Brh/HO0Q2f0+XiPmav3bC8B1ex8+Jlh+Bq4Dy+u5xaDZWqlhtHZi4BNjd64ZgUamUky/MWPjpCnZ
4JvB2kBMdfIdKeJ37DI/v1M4bFQB5Jsd0mhLmHGbGIOtyy+hIaR6wCmk4sV4XufH6Z88MyORH7Ux
x8XptLx4fk5yQvBnLcn6eXviwVZJNuhKg2UQNrVqiT7X5Gv23lQe4cC5aXS49fIJ+DLG1L2L4IJB
n1jCIhBKSFT2ThT4Cvk/j8EFV6UWYgHi9WUv3zY5vktxlZNK0j8ltjo+aGmjXsL6dvairVvJg+AJ
wZF4hl4yGF8Al/Avufo0B0iZvuV1JnscTUGuOZ2ygy3PPut0zL7VS+4CYvSyNdDlW0vW/diY7sUN
iAz6IdcE431OMh6cWoxIlSXpI0GNchPHCwq5j0KZeUK8AFLJy3zpOafMaJPJuTlPeXEY+Fn+j5/D
yV2I3zCHl5suK2OHBKsmlHnyjmCiSagD4WbIY48KY00Q++Ze1VH5Li3k6LRs/dmdQQJUvlvkCwEF
w/FJE5g2YNTVRwDl0yReVmwufDNS9YdrkFyqkh1q9mnjqJgRWju+Vrm8HoOSZ37eUNd3jvrKQ7CK
n17NQzfazkOck22untlalvriq/sqXQL38G9LBjRgVCYbiDB7Bv6CKH58T6KVfunGAJEEdQj6uEri
iyFYEAUAasaACIcwOiBCduEAaucniBT9k9ZpU3U/X5EFxtzPlQWv/UC9V7SwXoPKxvQXTZ2WcHsd
+X1UPHH3Zb6certPtqElDhkG0t050HKPCeKoW7ZuS6n0XPMYw37IzRGpl3izmrL+NaPrPI/3uqLy
tzKL5YbritxqSz+Kz8RcsUbf9kF6p56fVnkV1FsAgqRYhRqz6onWBgfT9IvrHlSursHP0faY5JwV
Da9V9CYRnum8zLoP37ac/+3Z9P/+/I4ba/RHCW62EDZTOk14Tv92n63CShVZ3tZ/HPIK7N03O/u5
hDVUyEoDyuprIIQM2N8JopJcG7/4n0Lr4WmnmHddOuhLCLSqnklFSIkwV1xT6yWiDB2tP4vYxTUv
IRTbZaWANz6O5Wpp6iuOkHo1tA1MHaE2EBL64xS2arXfy0sDO2ttoNqMJocXop4sm6v8iWd4XVg1
yb+GGjDrp1NNe9aCHLcOW2RDT6EFxUI/D7vhu7P0XQt6ZfBzDGY0caVOD35y06AkTTePEH1ltryw
OEwlDR+L7HGppA5BuXs1Alch3C0wZs9bL1qDIGS7IsPPGX5zjkH0sxuUa5Pt847TKrNp6NtPGOVq
PHFy59BuWvNRjo4KNGEwWxVBXvZ4B2IQ+gFGL+o3+XRmmqCkZHNACDyNh0b5XFahmUYSuGlJPoyH
MCoKrHXivUZ4uMHrNq5/Nw5EV5lDkiFJhC6U1UWUfeAZYLndIf3SiMnfV4gXyST7Khj3han+/lTU
lIJxLC2Vt1vVKTDTcoHU4E3nocnsfirX5bAjFMPPBBTQaP6qkfg3jQDneelbTi/DUBxS1DdFpbD7
//2MRZl0k+k6tuaW60dDYWzN0eXdSfsFFeREbasapV9woYdzo+CiRVrxv6drFuIuOOWz4sXQUEXY
sLea3MHcWTBBjtTpxBVTijyv7ESxvA0Uk5C70A3bgHmeNnhzsNwx+epgUWQxqLqv+lOzHw2RTg1k
Ws1qYEHGIYdPecZg96cNb6F+UX7wq0tiDeDi+LLC37yTA/BTVbfZ9DkkJNNsAbndHsu5kmGWEIr9
+iljNjm9Ofj8WYYi3mqYeihoHPcqXxb5eVwDKd2KKPcn5+YKv6kEn4ld6d/6nwzD4+IaVBVUTfsr
rtth7MASRtG0OFeoMpkvB6AUKpDpu4DwxAKaFWu2piM0RZqaj7xeRlSucj9gG8LRLs1UCR2Lk1HV
kSmScbRcUQWJ332b2jx1R8wVUij9JlPUJaPn1VMcBQ3NTYHxJbDiPcOkm/TmBaCPQdILIIg7PJo0
i/dv53L2IAo9UodvV9dVDrMOchmBm2Y6Ep3UoscOXPoUkfb2OCWFLHCMlsoyjCxbfuRIwe8If5fR
xHWaM1u1BvPM2INlpDHKe7azTYOAEngBJXxJ/hWhK37/I2hO10EqEszu4DYGx1ABhwyfip4wDmPp
p7x//b+kmWlfltU6rSxu0ucGoKpljNxl8yrWJfOA8YCNU5Lqhz1TU3O0PbfcD03nH2sB08GfmQyE
nXf2rZO+tykc90TmW41tzMR9ZCktlK/mW5JVO0Xk04E11owv7R61CNYJPfVRjC/hWPWEHabdVeO7
DtLypVmoYG6iwAXshgg8eiICPaUc5zJ0KJeka1Afm/qgTDe5VteIsY6ZMiYG5jbKzcjqcrIjzmsd
+CliNmg937SHLGEIoJv35cDb8n79bswpt9aSHVVQAlFJKWGmNG7aHlsHoj84dYomyzHKyX7ojD7L
E08XLhWF/B5PvWsPRbHaeDm7uRia6Y5y+0oy17MaEKZgYORwpITYMa+6rJCE7/NlSsl6rEv/+r0F
QlXCCAv/czgJ/mjibT1LmVQOJ6+J+xh9SVJ+I+tiju7C8XrNxfEd10KdFtSZUqtWCl67jQJ0D/K/
N9d0W8nl/D31CloBphvKMEFkzz3K9Na7100GhFjgieGshj9aqqNhdvymWMhcDhI20EPr5l49owig
Fu4Hf/+K8GS+vhGbboy4un1ARdNCHIPT7JqwSlpR9cAxwJ0PHAMZ9NUDTp36pvvDEGNiy17eWrMa
9w+aa34nIlA0uAti0aYFk2OnLWZVQzXad5e2gOXLPV8E7Uh6K3J0hQZAeagZ2sPt36kuPYXuNuLE
Lc0/j34gJf0e7BI0m70VwaQI1taQN50Y8yTIoXH7CP0eqJBAd9xEPZ8dA5nekIKPWZQYdoX4159V
GyPkSkjrYbawTk37AqALbTzNEUSdQ/Cs3O3ofU0s/R0RoutzH4u+JT8AhrYhcgGkmXrOU6HEQe6r
mWAIGLjNlwtCLTp+zqfjEwBg8pEf7mXP+HMbOVKxGo0WCDurfVYpiJKSN4EAoKyDulhZtZeIS/tV
7QHkekjkArQV+V73w9nX6DDLHYRK/oHnnF9SRViYqSEpdSKhqcbZYXZBiSBfRkLARnpnGEOq7Ie6
n58iZTmlk7flcv93VYmQi6bGylftHhObgHJCXk8d36K7aHXZAZM3U8PWQYR+v8mcftaTh3VCwy6H
6C96AiHK6DdINMqc0PphZuyeoNEXGryhvC6B2OyD7yPYfl/UWEv/cU2No9WspwZb5rfN0bC6pb8f
TdqHM1jRLEE0NRBfhX94uTWpDFnTHrmAp5azd5zs7OGeWnelETPObzlDu+tLg/IIrCbOZ/5QFJrV
Rrz8nRIup36o909IiYRJl4suOzftJ3y2Xb/8EnX5hBGM9WSAMVbpwpjqrWnXtUFsvIYffiqcHDNd
38e0EIKTR2s91VIIHYzzeGWskB94PTomWeaTM12jg+4Po2t+NUwqpWz9ebd3kzoGoOyqTKMANn5C
820HztonGdRjBrjb97IbyFalGf446XrNZL2wVNCAqL5x22gXEatPRc0C6wGSHGMVA1DnRN24S+fY
r1ZjLWn7aSXx0qZbQFl+1gn2/5+SSr9DYtiNs9C3ESAVYGlu1ctUQWCul/fb/mfVLlxAtTXhsGIH
zoKGvbPqMHHa+oRnCfVFD7UNZlEYeFecQgkRqs+cqjm4FL4h0uKRMuKqr5w7a+sECln3Vj+ctXzl
C97Cn01nY1k2jexfghBhVQ+c5t2a8kysxn7ABOM4SRF9VG7/C0cvp+N/oVgcuU3uZT+lEUiJhYqk
92gcifKY6RDTP8GhL107aIgScX+4mD9oBQuK5LV2p2n3uFDiRhdn/1ELgQfo8IPiaZzt+A0T4shI
jpddJHXDu34Jo2/vNt1JNlgCXD26PA1zl3KX5ZuuG7U2e0cvhY1m5I8JF/53kKOzblx8GxmluIiP
0umIKZObXsyY9Ru5UC2HwBWfscc4eOzcQeQO+cEO8n5NbdVtWWd754dkIrKHUQmlMHcirw+uM9Cr
6xv36lMDFhzSiejGAz4RmMKq1ARNnwjKd3gSScHk6V+vCiddnvz+d9Nv9b+b2URv2gJjJRWUvYBg
Lo2UEHm3lWIvz1ybpe98Nr4n8FZ1cDMUxx4LX5HmfCzsmkEFJuBeCjCgqibSYRHYSvHWo5CvRSVy
/zqMYRGakiXGtRsG8qYJMYOmpcAorjSRkK9Cu8+RVtLU+mVZcylBeDPXPCKh+CImJXWycddHP9Io
BfHShwfdvjbGU/O4Q5fUdpnxYixO+rzwyY1XJDObnTU4JjgonjOxP1RK6WKFZL2WTDf0AZ3LmlLG
VVBTkqMFIl1qOWz9sAti9LpItLglt/H9BnUKpe13yQqb2grB2fTHQWgLAsMZc5j68kLvIsb9NuiF
PTGZ4dgkA6SCwYnZQFGpursdwcIKqogiR5+XUeKYw5uDM3V2l7hJ2ETxAz91j/TndNWOjA+FRE7n
KNWyGbwmVy4zadkrTuxvhlqmwcLcKRx4BrU7iHvwz00zpWX4G/bI0k27ffUliFF3bcVMOyKbmgwe
aYWdvugII/j27INl+z92FS63U3YVMYwfNpJJUOXZvFcU6zUwa41Qdhdc00hvsmP1Q0dmzTYgeUbM
3/ehFcJm2rkaMKBajx+AvCS2FW4nbnyzZOBLken4Fia7Wk45iwuLBI7EyVBXOM6v/4tCHK+SWasn
9G+DFEJohOrOp1kjFBrVoJCjfMVKHfbglAfIToN8kPOFRufh9aEZ4iksqAEB9OaKB63JfBt9iBBu
QHCGaFImkHveIdgw27tme4uUf0y+7/NpiQ07gjKP0SE5EOyNiOpg768uMekl+la0n3Ew46GDoKl0
SCciyUka7++IMBJF0XqGOFLkIgRks93f0pz7ZGqN3OO4OzrGt+v3OlB1BHo1/UdxvT8LTpxb82Dh
wKRx3W0aWfx3QyQI6txQQ7oYSkX+AJEAt4xnmkylL4nIYz6+yTNSpJXUvb6H0+uTk1MOQYEGLtCi
FZHP/SJNXsa3Zwl9IlqDjY92thVe92/aiSlXEUJ/Dq0oa0mrn/WNER+WF/jfU4qNo74ET3HZqDbH
/jgUNrzGr/3M7qwIVa6sExCnkxn3ke4v5Sr7155G8UiiFeSxOb/8erPT1Po94NHNa16UmkkjVJ24
TRjj+mYzw7jjMkTO9WI55LG5VaDV61E90My+JO1WxafBX3IEOP0u+yOvBUejf+Bbw/XkNXWHrAN2
Be15RtJDk00Q2KQ39WpIAv0NR60MurusG1kR2+A07cB+liXm7OtWfsCiXzrHFKrMJ8IqpuZ+BRTc
SnKOtB7Np7lEo9Jevp1byfsiuf0+lIUa5iqRTb812Scyvqm8Cd6Su/0LH2tFgY3GV0oHr3P1+bx0
7ZTaR/ok2PpP1UOLBRqElwNw8rf6NJGJeffd/k44HUFqEGjf2RjggknlloivbxiwUHMpxsxhDIfK
ix2uhFcRU15QjG20jmFolVrCgszwvDlfzKUaczoi2lnPPd5u0jsBRrbtpJGwyAgyOWD/fi8OwkH5
3KMrWnezaOmTkw3MYYHjLncKjIv0qvSBqKsieG6Qz+ZoZujkK+/Skyan8LhQuot5XJuyiDR4gtW9
UhRGidojhCEeFOIX3TNDObXXnLc8MuQJXLZh4OiW2mqsVDiSYweSRxvLAhEQHWX6iRJIkC9ubY/2
ywASechjLDVROk8cx8LW1UgNX1pyATxLbAZOOlO7Nt4Rp5x/B0s1Dvg3Xm9QzLDd6px3iMKd3r8U
3g9BTRpSE+GDePD0X2LGi9nXyTXvdAZaPw+8nF1XWf/XDfN4kmB/HCUDwS/MqjVLAmhhWzjzgmjy
zgWpcuKQga4bKWc+xzthbIB9epLG/g8T9haWTiHeHn/dkLTYQkjjMEyEiGk8edKE+FHDksFfzAus
PqeXjj3DK4HhDPDUlIq/5H6tOS4bx0PCpc47N+C2smELOb3JLY10bZeYT0zSmEW8f7U441c4dAmm
zxRbLHo8/4bMYzcOQ9EOXumXrH65XEISMg8Dj03oUe0txJ0nYScxemebgECJJaIR4Qny29rhdnNM
uxipu/nW/FHVKeIC2J2zOgeYwUhlbvnjcXhp7y/rJDvhqowDCqYXCd7RkbPCG8XZUgs+KxXHQSxr
joVl/7mEL5p1ijkpPBPzT57c3kbjBr7SR0G423gx7PltGtbEXMC/Vgr8rpzvBN751iZDj2UmsVWG
6A6W+tvOLtJyBfJuMg1uKiFkwMUWhoOEvEHcXCiw8tcjQ9lrhmcuj6GAeaEUbQgYIKxkjyvTmVOU
73b7g+rVYa2MCg/KKRVP4YyNliQFx2BfcqSr6xO5GNJD18xBoAqIIBJxk8RyUnny4pQ/B56TIL2t
NxHm6OpSTl1MCjPAzT3rW8IDBN2/6S/o/e/SjRCK53GmQUjfP4cHyBNOIJtrJAZdX1HJCXY/HRQM
Rfxjl/cI3IgtlEX/1RUwdyCbOtOY+stjSwo5NjpOjHbAoes7Fsbvh8v8Bz4J1iWSEJLT6QZwFuWc
6E8G20V48Gq0h+u8j6dilNzpyAWJtWO1LdKWcXMI0eMQJCkC8NGm81YsXK4xpymbthaaHR93VAaL
nsF3D6z8EY7W0ihhIkkrVlhiMt3DouBd3bBJuXDcdORmdleyKhKtkYyQh8SG9fz6vGouDC9aoL49
wYzLydC6yt6tRq0mvJwdn5q7gFV1qr4KM/JIzSsH9JbEytLPw639dkSW0vrmt5ILKDo1ZU3nAlE+
59+oHiVO8cEcvmRlzqZDy97PnI83A0Dg4aMMQE5Pl5kwtE1ZvROKUcZsKlot+Hx028mfH7VkSdnR
A1m0lck02kQhHi9BpOJNts38kqVXaSfvS3FLFrHkSnJrv/x5zRcjGMKV4w3/aBif3CivLURwaY3M
GL7MEGBtiqR38KT4DM+xRdt4NOeshG8czKcqU3XukemO60c7pUJywV3/EPbsAY5S7/RGDkLAaYHB
h4HCPu56pmaeBY6JjIGq1+lhos05kTS1jmtMyXGGXsE+C4F1ZdnnkzSpiIO5e8sugQCJRr7Ud9P2
W7iLIzMvqH0w7QsrmN/7hCEvk2NU8gE4ZdOjh6quEVhB+ojRLp9444G++JnSuDe+gzlvXRBWp2zm
iPo/eZos46Brw6xi2bWaNxQe4acz66eIk6/y4gr4/Ef/98buVMVpL+N6AaRudXc4Ul0A8JtKCb6D
xJ0tsCvQ3D0NjKD2BHc9inC6d8FdPwXEGZnvekRXeYyciqv3Wg/KtBDGosYbF6gx1gajGlJuQvf2
yZpHxf0yxLY8ZjCXzuOziQYNEkHTS36PAraS5/aR4Gjroj+TCJeh3PkQdeUv8DJbX4sivOt9Up50
pHQH5CRMZQzeXxTta2MIv38UoTGgg+dGT5cv8ubnFekvBiaEf2O7gqkHA8Bkb8FSHoKiCqrDeJkC
WMIgE74c0mO5ijlm5X5WwzWvmSalepF07s7CJZ1iKwnV59Q0P114mubeZuEELxONjuvfigwTsvsR
WTlVPeARKuhKzFBmtiuofW99Qo+Y6XI6y5wpY8Arrt+/DVe/JoFOFhmENI7c1Pqu3FcBVWK+G7iy
aQ3QzwsBMNsHX6EtesY9B6dTixbL+6oJQTHBmCAlkRzKNJZDtrTCBNpw6OYB1MK2kStyS4IjDbeC
cy73q5SeyNlVluXnzeK3gNkfFLcDHbefMO4hCTOr5lPRxGy+dxcRWItgsDC/D16+z7F3oZ/P/otA
NEPCzM/mF0AP3nzgkg4jIVwSKhRx+sOqSYmXG5PRUHfW4R9MocjowA59Q44sJ1pjX1wAJxtcTQtT
BUyGF1g/QyX8tRGtgfaTOyAKiY7PfHbrJMwhbfCyxpvoFZk865ZJhIQ42wUEm4bt4vfN8KUVAQmQ
aXwXhr+vi78rrvG3xKXToGb/JB3vVJkCr+ToZzoAo0xtHoBY4z4NzYg9I+SJAkYvsXt5PAUtTDBt
BYE+GXB9aRD9JcvWALrVrECjQUn+wLJU1XFAGSKUWVhtAUgHg4o1IfW52xI0Mhi/XdcojbFzunuK
PU41ss72O7WKYCmylYJ3272ynjfwlt60O0Ha5Ab3lj+VYtsPHyucgPOWjeOxVn6purKHvL1WRXNR
cKqXtgt2g4/jaVZH9BlIB/SGXXhs9kw44QpBbmTvQgJuwjy+e7J1W2j3TF0eHQgpSTeX6Li2Jon2
sbgFxBI1P6pApAcI+h7co5JpJ4UDfnsgk7pT662jzxuTJNHqQ1CIhf0Np71MNpg+NAR3H44S6MkZ
NvpPjGYiqd+h3rzt7mY7r2I0gRKueH4k1LRHmSErl5kOATz92gpI8yDKpobA0gnAG3TuYk8s11oO
fDDIbpfcSyTpwbsa3NnLX2ifGA+1uzBKh9CS1wmV05RfsTV4c7pNZJD0QXpbp+QT2jF+TI3vJSBy
zpWiuCscTaHgNm1xhIuK699Hs6lr9U1QIy6VuN0FjVOqqpNomU80EDuIrfi/n8Q89Uisfhaph9Yh
bMJGVd6ezB0YBr3H71VLoVlRL1DiT2G0ieM5AwSGgtrqCafWn098nwbjD4gl+YLBg2lUzpmftKru
AQ7ja7273m/Y7g+CEzRlUTlf/8Yh4okuN974bVkA3l7/HjLKYYu8e/W2evmOhkIKFx/LwoDZ0im+
N1/Qs44RyiQ1cJPrwWJ1GTiVe/SDz/WJhKPDSreoM0A8PG8Yff3eim/7A46wz9clujr33u7ljmzA
jHyDAhaBl/RQB/I5dZ/OxytPmTm/OEB0CGJ3FShd0fcNFkDZvgWO8QDCc0s5Zrp9bGLfP3Xkp8pd
4k1aAkBQqjwbtieG7BJB1+SMLbWfGF5/K2BX7tqtP2n9G5HFXxXPG+cPnk8o6RJ3x6TOTqk1EPwz
ofogou2eVCYwr888unYZMYBDxaHvvFQizHmTEkq2t8RWTBHdNVbHgCtad+WVm6cjkyTjEKwkxsvd
gfeKNtO2bPRWPJBlrtul20NGskeLHPdufuXfNlTGCG9P9NnGWWvfnZW/EhnCqfZNV+eoggrh1biY
/Mi2r1CEqGnZ4r+RkoMJk9M/3soOUjcxR0mqOKWDQGZrN7WDLTacuDsBjKKAEpqTFWbsD2Bwa2YE
7asLKKAIqXU7NlxOeNsbR/OYYm9lFTpoefWT0sgh4+3SDhE1JX1c9wZ/+hm5/6LIyC130CpQAhXk
6fLiFJFdOjMZe5ctYr/u8yAFS8M/zRWOk9gO+pPe1OCIjIFKNsas1u0Q1RF38eQh8fQUWmPbRHjU
jUj1osOAid8m9Xmgbv7mpwlTgnusu65c6zLP2Tej12nyghTLm/ZNz6H1a645xUMWJ9dNF8ySiLFW
8Bs6sjl8QMQpuJGvAp6r0ejqJktBlmDKVhZXtPyZ35INHsrvgBuCIiqFnrE3CyOAbtD3vbdcD/A8
breQnfHP0xYG2QcsKQ1WAzOPpLGPwM/WykMy1zjtXy8tRmTR6KeqrkvuhLEckXIs0u9rVDVS1vXn
hXv23BpVxCJs53DM8jj6voaKzxeHnr53IjKsf1LhjAmpV7/oQf2TPZeXwxloafWFJNiKwkbrv5Ro
klXV0ySgQOZqptrQycwJBdCmDd7sSi5prlzAftQDLU98QNa7mEuNWETAibVZ8v+8PYBqyfDyRg3T
/0q/85NlBUVH+bu6tCEAsqAmXp1PUCRi8Yt6AeyDEOoLDtUWLFkUJ+gTWeQw47dF5WkkjNEyWQpL
4Qm9CMGcCSAp6JPvb8rRse8C7AzCzpe6rUNYz4J0Qe7yrxNZCfSB44tjm/3SSHL7iYwMnEb6oGbp
BxNsZ7StydJYJXQ/syCgQ6QMbEuy7f+TpvYcTHxQ7uMTMRtWhmrq5mUvpG0ouoxSZs7kg/k2xQ6q
vGcXAd11Onkkb/VnSh/QDYW47F2mqrzFZ0iCLGEDpQ8k33JBa5zHzdpAc0v7ZUc4Kn49u00XH6iR
JjqSfb2lfHypk3ykoaU8xGfL5E824XThGODDkxtfY3CC40tY/sFj/hL5kArMJruXKx8UfebH9L3x
25kMfKzh+YOlkos7e2Zmfky7YqXhP1qphtTOv0tAauNJMM/iuhGActynDAz0uq4hTNeKkEzWyHoo
IL9X5DlTWRArGqKutxPXM5N9SNjGcZlenFnUoHng85RmeCyiOqonlP/GxKuINFmYvZDG83/UzHPq
b77NrUu+MJbv+VExVxGxVrLStz1mzOd41K/DBoyjUA29destVM7eTQIEyFirBSXFQ8uF6vhlEXEJ
4V+nNIqba6BT6bdT0qm2Bj29eQDCWsg17TwsODqywEs9Tf4vuTFKGRcwZxOCkBj8jnwvHOnf3SwW
kDVC1jMrcLN7sCFjL7rLQAysRQCfj5cVz5Ck8HGsTTjaGgQo/vXdqUkWaTgy/WGXD1e+/UvVpFzS
RN9f0hguz85Ijy/sOqk+1O4wkMaIsJyO6BTtl3K7ZKcsdE/LhgeCEWPCTYm2exAIW2s1Q44JLbfu
S8QB6C8kAxB9kh4D641N02nU7ibHsfshTFHAeE93e6FTXcTaMGBAQgNca8q4FLBLm24MizmwCJ2r
9/OxiGymeXjz5agHS4liPS2Zr+rbu/N/zQ3yoeBXF38fnCWEpNI+Hl/9px1TvtyouFHA4x290b0k
tIs/POU/fJNVUF6V/dW5kf8QvjW+pDLvmn82sOKFDsRtnIPb/Swjbjn6AEvFaHXs8+H4ztZeXFI8
QWrO9MixdSz9qEl1KTvEgrBtcPJbt1bbYhfCZeNa+RxMvLXG2Abh0mR3MoA8SSm7TKYB2fbdmae4
gGeMc7Sc1F4997YEAfmqvdvf1k5OFnouL46+U0EjHW8s3e3ds3OQK8Vhnh3ZL9cYLzxq/OPqXoWA
EXuvrRv8s/Jq2SHu+ZZHKYzAP4AYVAbVg/xqygMq95SgA3nHnS8DZRi7l3Hs24h896zq37gkrC4R
Pxk/i4gvh9w8K2R4vKLcp4j+Ids51q4IaYQmwWhxuz6CyHZmsDcDN3QjrnHknm6WjKiJTHBLbtQQ
CFARtWrN/Fvs011BOQ0oQBe/VwLYkG8ZigrKUg8S4ON2Mkxuw2iUJtt442RJ30tFGQfpEPOC06kn
pTJAY/Vmi0uvORtfa2At/vCax8nQV6rz2yU5uUUdzc/CrTG/VJnqzcZX/fmJYwZm2IBkyCXFFy2h
1ln7jxinVtFiNfaI1u+uYFVfPCyhatxjZqPQq0XZ0tVQ1AT7OoDKrxbC1p1VDR6QqbMe+OkAUZJZ
alQEuqUEHc9RryVl23GSW+CZ4qZ1b8uTybOyUs2eidM4qo4xatcNiWlxGFUgjTRYPXRAfK1AA3Rx
tBIvjJqXh8vDJ0bXyahImGHEkYgpM9rRvrPj2iragXTc58sMs5G0Zc+D6SEkZ0t7tJzNf8EuN6wU
w2YXceUdYmcSf0oMAFELBrldjSBaS8F0nUNTFQA7KPfcBVA1nr+POL7CEuG5+z6m0908JW5o6Bfe
OsXUsv/OzKpJFi7T0zFoc8ZsmBBeclFzYTOX+ml4ZQyd3cR0gWszwo9om2XydmsHN1hPEOEIGhMw
g8yY4OZvXNGtX7vDiO/qz/pVIVWuWR2GqKacisJI6c1e+ntpyUUufx/m13Lw/HELl5wknq2Wb8wu
ZSqInvWWQtElNeGxPYnWGNOjCpvPtkVcmPSr9NZj89o/gBDXeClMjKI5YAv6QUIFsz34B7/Xobon
2x1/XikaVZnTdSDiZkS/XjwsfQDE52PS/UeG7nrXCklPQWxsTH//yIN4ex1VyIbzbeDT6gQHjIHR
tiQFv1gQH0REEOABbBLq8HkQSx5GAYIvYac8EnXpqL9BSJ2PEsWLk+NCqcfrbu6sMTOp/AAz36C2
e1E4lNjASP1iLgHoGz+fkE8x7buUxWAMPTOY7a2lb4A8O6gqLWF4scRuqcSjR0P93/Ks9IqG7Dzb
40IVLVQXLI2osjyv5sXGdyY+mFsc3kh750x4H9gkk/+41ONOko2OVunmxs1GMpYWjDDT9kNfqGZs
8cVEBgioBIT/UO6c4zZQZXf9Je6GHyTbKvL/ZLaulh8geFti4xv+MGTi3+Fy1nXqXl5Nk3Rh0LLo
Jgi4RSOzH6o1O4D3Wt7WHdINJpBnU9vCoXvB8NlB5u33SOJjDgq5TY9NBfrCN+M0R4fSuKbDRIW0
pBXWy0FBM6ePj7W/tkKApZHfkSclB1wFAOeMFrywqeA3jRNPlap+EGfTUnhXUgwfvB+ZWfAfBgqO
JLk5iPxi7HE0U1Krcge+1rYiOs5g52hYC09UuEtXd+YZQkqqkJGwTz+Lz3eBRQ4rwaH6EmkGuWi8
Z/FFn6se2S8BjBNLBudZAouRXbBVSODt9KIBIqAZyu0AmyzL6oJeH5jatUnudUMuV6jOT2rnjj74
HV2+RAovri5BrYQAZf9yXOB1cq0CnzJ7anVRnNHDC/SzxlOvN2SPa0vbL2cj/eJZN49AB7K1+ZQb
5Eh4++ffZvXgmpuXd6jHyjF0Slc8w2rKn2xkHvlvWFQT6lcbYPIZ5ag03jAXLIPECbfv0kGACBCn
MZgS4IQMB/uQeSAi101qBRoq7v+NeMVz23LfYU7c8xIwDFni79L+VZq4F5//yR8PtKWTHLHNbjWV
KLK3XuZcm+sksntpIueafS+Bpd9mcbSZK9dKURk6bdewuP+Hs0nRzpJCyVLTh/5A/Cq+lHOMk4up
3BJruZNG4DKTyK5pnxSSP3vRtSsKlJvKuoeIuk+sj+RsrMKzi/iUB9aRVA/3T2spgx9n4559+OYa
ePUMZHBB1ASOX+QqfqJbQrxnQH9oi6gQ6kBRTzOjAB534JZcYZ/hELq9xqFBYh6SWPY1QW5ipC5R
ur8ulS39FppdpahvI6yYU2ln/i3pZFUbZvCDId+JXDA/kf5ydxgGltKZbHupqkukyKsVH8Q7TmtT
ffanAEfZ22gAL2uZr9w0hvNdc7l+UbEKL7wQPrfSzeLG8Yz8sSyExH95nSZD357wjz/13562RHGZ
ya026w6GYZmGsU5Rz4Z27I2QJ6JAk6qss9uqJzbHvy3uGWhqDgSDR3HvE4qDblb2lfmdYfN917eb
FmEylPqjYG7Aw5416uEtxHHu/SDBy3b+g5sXYUO6/ddVkm6tFBfNnvzUJoWRCrsM/8BCyZ5KsH+O
CsoYg9icpjWdRzNnI1Xz2FaGhrZWB5Llv7AurcAQIqAALpW6m1EzTnshEIyjR8Yc9mQjH72L/Arc
jcUNxaAWGiENdyusRwdOPZaRz14RNllBw6qGrDL6Ckirr2zrb0P7HmQ44aK53EzOCe1DeYv8JERd
UiM51mIFbQl7hPP4HQADXO1T1W5oZ46HSPm6kEn9gg/QzbErPwl0OJzDQb1SI7hkqu4FT37l91pD
+hokBM7hQkSAF85Ev8hn+s+/nxvoKl7OER8csiVn97EBTNC6OJqtk4NNXqhKmR9eypPuHG4F8BZn
bQAlOLBDEbALdFn/DD5oAapCByHlmSMIxb1gMW4MF8DYWjm3AAjHEbD8uymTSv59CNq6sGp+C/pV
kb9hnw5xpXBvPcCv2b6dAwTh2RojWetfU0hjnQ5/NaKXxFQy5vRHEkWrni4XwHk6qGA5Bq+nruyd
W7Lz0S2PAvB7HrB8ZrJsNAdzlCt86p7aOurXW6uyjrlfXumB+Kp37py9/s50vLcIwYIFQpwzS3aU
fvKJ8On/fvYbF8Ysax3DtjsKSiWbEfQiPSn7Soro5QFU7Cv0gaEbVj8AbwFdWdYEsHYZkKzIdsVu
VcToWtswXQyZ8IO15y7AdhFRe+1x9gulzgb4I4QFVBzbvX0RbgbUl/jeIr/IVkpO4LtLdix1w30u
g7NFScO8ZpdjvxFab+tliZvSLbupbJMQ1B2RNIlKIr02R3uFK4EsVmzeeUZc3gNCP/aCT+bU63ks
rl4Q3BZgPamn6A8oiLLW24wmU1fuD45DinRcfXKf5u7Ks63BKeQA2ZjD4qqb+WCSZrYYoeQrlAm6
l54WfMbgLzIEm4FR17iizH6Lf+lIvj6aD8tjBBV90Bh1HzOSBybXNydYpUrmB/0EQPzaNQFn6jOK
+hfX2yQ2Hq2eh+h29fIJ3CeqghkZ1btfsVHIXGA2kqTRPaSTthwB3B6V3FKaGy1iAOx0OhOkRN81
6oYbKAghVcR6sX1pKf/0oSe22HNi4ux50B3TXrmrcUpkeVnIzP53tX0euz800Y/qSzNjOgy1VWs7
So/VEGXeTy1jp4YwL/W01o+BVScwzqNw6zYaLzwiyuhhMlUjZJVRpLkt1DiLCStr9jNK1ate/NqT
BcNV/N9qP0/WVAA8lvNNUCpUuZAJ28ZuueT7l0ax8twStg8s310QlyihalsdlY34SxRKO1kyq8Pj
AKU799Dbqy7ITA9jBzBbD10ESuxwzPNFX5ufqn736VJNf2tQ0oe1/eFjAHblIGQR7lT4soC+VGY1
7WhVvJKEiKdPgVIA/rMC8dPV/3jB3tru8IFGx/8ZqzD2PO9aZD89NtjdDrNUgQnqjNslIc9wxxOY
RUPcaw+Li9/0wmfezGi0lrJzQ4wDZ9Uph56sR+3zGia2Z1EtDsqtcfglvA9Q8ImXKVXF/yvoslFv
L5yPaiOPrHdQrMrYz8oMAGXBNwl835gyewoxhgd+KIo8xIAAvrodWpwmeIRPwhWQDO5IL2tNfG3x
3vK+53k5dZWScLgx1QtDZ4mNk9MeYqDGILVIGpftFRl0aucMBpnaCWNSdf+8cTXs+RjR0IY4wNjy
bdVEv730OuPRgprY4k8PAT6wicfMWKopg1KRcxwg4K09G96GjxCab8tNc/StB6mQUb3gbdBJwT5y
KSD9lYthDjvGtDGYRY8uukEC0FJOs7K22Onc9+r8L4kceBkh1FkoeQMLoRBtAq7WeiRzdmmZ44Ly
KCrUQ/B0KlFkxT1xXh7o7fOti94vRvHuy2UyU8/NE+a5nHiziSnCsufC1k1dzsdZNKCJgDL8nU9f
MA1NuLBo2UydrNgRny3VWC4k1Hi2Emz5Ju2AKvEGH6uQpwHp6zoORhvNSwiXPs4WILXQErBD9JMR
i7Meex1ekmLrrjBJKe891p9sZMHU+3SHFbEseKzsbNjUvmlFkGk97w4j6KiCiw2o19QobRRKlNRv
TOWrwCR9krpuIyaPvt7yJpFQFLY47mOjkmupZXYMZ+QAQbLQtjwD5HvrAXd6OBHnLyyivJhN8ey9
y2AzmreiPY+0wUw1/X8S3AHFlFZoyoOYLwPjNDuemQcF53Nx1NneTm40rW7miy1gFOc3bfcgOgJ4
0j8mBKhwxRchZLFQfoezlD8nPscZrnxdWd1AzHANxOfsHCKjJOMtiClwDA03+owI3Oxc9ojtmLVJ
rE2uTyrT25HJ8f93FhT0Ulxx1jVtZY5Fe8tmUF3FNejSEgbTaE068wo8l8oDM450SdgAkmV2hs3w
H05JylGQsVK/w+IeNRatOugd278xMrqO0DNXZ6cE1+YZRpAGj6tCFeYJdI1vUZ/PuezLMjstM5X5
6AOIXeqwC2YVOJtUi038ndJ6pcjW+HDYad+ioLl7wqQ5i1DiiCxd4HZMgCIItnohfBLu9hBqazga
hM3yJrinxgqJeyZyc6jarnL5V3hFiHt/f+lnBp3x2l+ZscD/xMEAF/CNRmlQ2HBixKTX/pD9gOZC
x2Zwbw4azQYyhp/72zX7JZ2x8ql4cm5KmZVfvB40BSfRWExETogJdYtRle++OYvw1SblpOTzBFmc
koh/kJrGplc5ppSbRlCfydBttXfQSWnKTYhGGk1OBKY+pfGpszEhoqLV3ersA+49RmIxC3pcATC3
grJBHngGvsaoEvCXxEUsYbhxH3xKnn/UR6eowRA5bIOKMbminLOfrevbCGa9Xa0sC3JzV6Y5p6u8
uCcedOfU2gqqsXdHksfkuRqeVattXUV5F4LA/xVJm6XuJsAdMTcPh+ui03y6K1jEFE9vsfKSTn1s
t5DoP7n9NHo+0BRZ+/5rtKDdiroLCiP4ECeZ7SIbKxHWKCxCy6KXg/QhiQTyGftVeHSkaGfc6Mnn
ODmfpak6LO2vFzzz/94CPnU4TvmJdUi3zQPV9ra5Bf9x5oxErCvEVzdJ1vj8R9autUvLlc64Z9kp
QUpQ4VK5eLDjKhy45BVf0fcv5L4V4f+S9jccSwGF2vlHJMz/y8qRTHezkqWygrr/u6jn57kIf5Kh
0XHOLkw8DcRTxfIsxFuujhNkTZp1HAEq2mc5LW/RJx7RvKXjM+ObjcGcMYPvcqLf1nZxtEw+Y4tu
tpXSFVC0r8Hp9QnKO2tuDOkzdKLHlpat771AGdeF4jXynOXlWK4rFxwNuE6T6+rH/od7Xz2H1pT9
dsWMERc7Uvld8hZsvH21SHpdvS7q1ZzJ/ETPVtT1ll1Fc3smdyP26Zw79FMbCFoAboqwoe7o7fBs
lDHF4s2wVXYpbHsc0aYJcWK9Zd+Bj+ZSZajhKCqqT6/5WS3IcWiEJTHEABpLYSWnzvJ8ihMMBNpt
nxAkly4mqs0ovQjPxd9uX+yxDGuRUMWXNdOcu9dA1gnx7E90GExEP0Gp5J+wp+rZWHhpe9IIvbVE
6kr0eTZQMDad0tvYOuOIbqx5viy8he++kFnpPumz+7HBtaFYbNJZUeyzOuSrHjQDBtHyN8ys8OjW
PLxJKBNaYAaWCbUe4N9xt6k/sbtlPM9aJv8BckUeHVGmy8jcsSyaYNLO4E+8Orbq25BDlpl/Wu9H
FSfFOWBnbaTop3NOD2cZo0a+hmRFzGBtc3gsR/FlP5Qpng9g5A5mDqXf/aDfcRqWVC7kFL6cabyS
doYv4DH7Fl5W/6yCX7NWR52/rzEUn6J65hmOamjBeG5C7HM/1EiFJlI27L1nyZJKCp64Mb2G3bVf
nmUcR0GDSky69sVqwNvqgf78LB/aVCE79SwsHydYM5qlUyTploQI8IOfliFciLUfe71bN6Mm3c3D
Osl9zNPgyg3o+EUvxTeAtIWf+Ikp5gbrR0Xi73eLlxG/8zwVbVsBKzWjm+BflS+oBhQ7/O1So8Qw
+62m5ZkvLkKC17TH7tY5ZdxthlS2gCuNTYtnMDJYy34tww25Uis9HqlilALjH9idX2xdtu39+a+m
j7cETD0ucth/HmF0xij1s0xbaLrLGSkDRzB65cZIonzjqhJmFtlZpWOJCcrn1yzuQUyihBoKgTcT
QHD4JK7NjhuzdE9QdnTqCOjep/w8sAj529/nokbD3vpwGEKaCZ357TCa2idxAyWCuhNN0cydblNl
N6QyBGIsH8cDdBLU13f+LCm7vmV4eayBtGGXFDxybjJ4suW3s4cJL3GKsz951UrLU7p1FNSklL1c
OJh2QN2E0mqn830ZvT7Sx+jW1DLXdyH0LDmC+vWS4npCOibGIzYRO0eypUJ2byHBojOrg7E1M0h7
v8A1oLC5E9Z5fUsgBVBvGYDSnlclNJRdaDGYPjTaPXs+QcMbFKqlrxuZ1pR3TAqL5AvqDHLvDYbG
sME/pkoNOVazd8CjJhN8WACvpv++OO/inD+YJCdXfpCPwnPhbCGCusyvw5P7ePfPsalBJQVWg1XE
l57qLZSV+ZhZ0Lz3f5wz39xTsPhzW+bcFpaUSMHJ6PM2IhDEz1x1Kh2pqTnDyiwZ3IzdKGksFtlg
lJmkN/plzrb/74fPIHeNmrjFs/bdonY5H/84NaG93LmdBNdCU8Fqf5sAMdSnbfE8Lv2oVeh8zkEH
2qrevMtiODf+xxIkhRXh2kOXLHld1i+uP2oXMoFomHHk88H95wYzEJJgU/YJocsAMn4b8rW8KsWm
dfucgPdcEVb47ZYTBvlm7JZh02aaotMr63xPp9+mdyUaZQIPieQvIudJTxt3GlSstAqzQw34JFNS
trUws3VAtwsX+j7nxjhRcT3y+faEcWjnkE6iqnNrEn80hZyxTirwVwFj8Zy2q5HWhKBIAL8QGJev
DzDl5rrSi1agxcE1D213lxHE1JN+TeBiKL7HbW5oi5T6KLtBkdXyvXg8KapnoMmrD8l5lxUvtACu
ndK1iA/kN52SEeI7XRh52LXSy0EI5K9HN625X724VRTgWPhjpSkCO6XdSkWzJ9cqVT2njAhM02AA
NrlXrL+ywzhBZDomBFiowwL0lGSyCRZF+grraBxUvm/+//nEsD5/k6HeVhmOeiaUnBVg9xVWXETp
293x5VBD5PteAR+ImEKf4bRc6GBe0LPg9r2r4Jm3pBTH9eWFYGVK4tqtlyZ6RZZI2JEXEnX+Nz2V
XjueKyMaDFUVC1ve4UgWSCDtoXF7urTM4UIT+GwRej/+m5JZ+8Jwv1EYewpdv07JBEWyudi46/fl
oUWXgiYOcizWjGAbEdowmZZO1M03fKqsypaMQpE/KgpQrmxNVeoom878qYkOYC5LQ6IffNPc0r+u
wgG44pNcGXScHg4kGAdguXWOZBrQgCA9WRYusCQNb/jcxioLfDiuo4P9mLHGci6iMUnoNO1j8ATj
JTrC7+DW53pVuoD3N5YGARwIGSCbQCQH7OPyPIrkWzima4N44una62f9uMDg2ZxjJ5ydrMGoRQTq
Jj0QO0DZH0ksAfNIHtHsKzdee+IOVUMf8egIWvMzaPiC5LX5z7sTt29C+8QU8vrLITjzOK3mL7g+
NQwTY3WbO1gN8tICh8hSmXTxoJkAtvtskBM17+NFf91Vc/lph6E5VszwEHFsfppXD/5T7TV5IdYq
lf4dIDg7gsRsvMnknDABgszcqYsJieZC/BbTdozRTVgRYdwpvko+K9W1gEeW2mXN4/m1eszcG7U6
lEVPmTR2BPySYQa0WmHC5J6e7jeiFyBwOESIniE3SBxXGgiu+nSgxP006cwN6dtT2pXwfTQX6PmL
6AggetFDv7lorQyLALuncgkxhuQ0MxmNZiONM5Ec8P75Fb40qQvl8RL9rRo0P8aprd6KKkJrohUF
HZm8ZndEGqo6ZEoSnk2diL7t5dn/HvZB+SxGeGzOAuwqgeH+PcgfVwR0xNEiworFtGRVp48Tq6q/
jcOXgjWtw6FDALqVpLjwA1HVAwIeLYIoQgAfsRbSpDJp2rZOl+8LB4biCws5Xu0J8MpJU4tpsvQc
NHwM+c3MJoiVruLs45oVcyUm7g4D1+65+/+jW2xOi2lFk9AOAnTdTm6LhEZNrBKcF0x71S5eD71U
rd6KngEmWn03ICHxCtDpeKOtqYy8/JKPoi1jiQV2PWXYF0hH391ITLqYKUCkv4lSDCuLau4nLUCb
Lg+iZJ5XE7F8sG9xlqFEEttFJqUpC+5m/QbS29tjtLOoI9Jsu0Y1xrZuL37kDFXbB2c8gOAVNMUG
x6j4CWFlnn41ZivB2ZAYDbb+3sTE+HhVUJhhRMY9r4Eo5jgIhO5ft+w35veyJpP30X/0Zk9hctTO
GlgKOCrLohA2T8b9I2xIbNeOZXoEUOfJfoQ+Ob7LjxJzZdHXHa/S4dAacem+CTPlUf2Mxu4Aectr
beDrVhmaExrFkDXsSZi+gIE3BXjkUy4mjAtt89DNRDejUgNjcoHwNm4IHtuaH/VhjJalrGl1eO/T
mECHC8/P0M2bMOqw0nua76ids60M+EkO/l57jjHlAGsGlSyuUx/IXufsR2kd3KlLleWLDcmBYlOU
IjEemdwx2RnrRPv3JE1whrHULRqjbUHOk9aD526lSD+zwbO39HjZ51TdCf9k7Ik3atvLU88K0bqs
o/2SOntFuAuwt7mnpLlfzEWyCSoRfZN9ddNm8lURSSK/ddcPFUn6lNLuL+FUtkv3FOreGloWg4aG
kSfiYd8tDS2qPgq6VQrLvjvr4mCupAvfMkDizPkqgrOrk/n86eGCybi6DjCCZAOBHP0t1TlWnwgo
+MzVolaXYZM7tXDl3AkijgWcfCPv4nBo7fszVC/P+ECufXjHq0WaYCAmIhq+uRWWum5v6QociVx9
SbId1Z6aHurni892Bm+XJ5WK6x9JzJ76szGnyM49mzBupmHKtYgM/zlh0Jo4rlIXHhRwUWZQD1F1
BwrIigQeREzOGrLhJuJWymwe5oQu1vSkH0goEXI06cB+y0B6rudPBnJ2bRLfiozs2jS4rkyL7RZB
ZZwdZITsN7xZJjKDq3ByjClI/nbb9aM+I2ozRxdf04Bw8b0EFceL1yQRKpav2G5jLmXOS+lqOdQj
liBd5RK9iwwOkMrcO5ekK4d81kCcshV/KEUhmMQ1WYkQrGXKN47gKMRSSoH9rPBQ9hz/B0f7Y3Db
c6/UerYtx/Izn28GeRJObzCcBpB6IkBHnKC+gz4mADD+jK8OWtnV9XVJ+5a8YGGOMTH3cvbH6n4b
OT4cERXpN3dnPF6QQmqy796aQWjJgKY9DBsu0mCuhTI17j6BObuQztBPiXjr4mom2q4Ts6KWMrvu
q2IqHwm1PfHkXC6KGKkJ1HAu2emzL93MzScemIXUS4bcNhCXpfvLv1Dxlst3Hyptg8YGL+E21abv
QauqHE5PkdDoUPImLk5VKslovLQVkg6LYHzkC7ICwFvWDi2k3USb1nuzR0iGwM62RkflXTxoW1xu
p5vGibHdM+GkPOQrV6tm5AnScwqnjULT+cufZsHYr+cXb+qy5PHDhTi5YGqr/YwtdUVyf11Rqsg5
a1/eJcc3F1ovfEovKUFGYW2hkqyS0oZryTGGiEoLUIB1uyFsTv+fb77fg0SdkmeU8EBfMVfD+AUR
OzeuavWrIywvgYy1GKiEMFt5IqarcoF2EgRPNxIrDidcNNG0nusOLhFRSzUngek3FVnHopSe7ejU
MxX2CIST/E/wGTqotug6qCxy6SOdNDuiwdJy9xJsdG8L7wv0h+veJouiPwBsZznDBI0QWPZBqcBI
INeVjLdRTK7S7UaDsQ3XBGm1s0r7riSEQdBM8kvfp6qhAhAZ221daOhkLMayy4aiZRjyiB1Wzfzy
R5XZquzkrwJTustpA2+E2aAyTyNMP2hE8s7QSbW7f6yNwQFYTKH/CuD+ngGR0M8DyDyfv1Z+ttBU
FX8JQUM8tlhbwBcDKYc7YEeG9SDtDidmIdUNksrAM+2LAEa7+87BX2LVHsW6luiYuGMi6tlkb9lH
KQCh8Wzqe1AYR9H7TEvXqUIBDe3dJ5jdnx/UFYYnpPrfMWjWgRfSL0LYmtSKsu5ZFU4k5uIHid9x
7J3Ya5GZes0dXAJUX9zvxYuG4fKc1ZASCWiwgW/6QtTXaq7asXMVViPs+LBTCqQk0Tn5Cc2D/7n0
nP+yZQZuIm7AOiLd4xXSGrJHLeNX2O/dcqjtnGw+soWP4ockJf+/d81Y06Mb4TyPcEVeSHyXVdPk
AHff3X8GGXutT81LvtLFD5kMI9c5Gmpu1j5RgsGfVbZWbH0s1OU6YkP+naWl1OGOi42sBymve1BR
BVXfyf+2uP5apUoRpSiowln1L+uvCAbSF6JJfXKJ+7jdBHeHZtT4Y+v6lG4jdMHi7H0zWqVaCppI
UkgOUf7UuXRQkGNmNPh4mTOxZ9QYI9HcMJY2MtRRzoR4PS/cwkrvEYVwvM/j/NdJ4aX4uuTlWenm
0DkLPaWyHTwthbmTTBy/fUB7gufUlfIrP2CahRS9G2+qVYeaDTVma4g1RSP9RzOUJ0ZaOopSQXDT
3rfzLRIsRxEoBSd6yebgxcVb6orTYXrz+JS91H6dKnCjLbPNq7SYOWU35tTZz5xERMW9F6OaGjUy
uFKXpzIkW0cBtialYh2dYWknmmMVXChRiKrxTW3he9zqs+B+oXc0tlhwyhni+RgJVHth5Pg1cogX
+hd/8RONe1Od9DXzeHV0HWG13FavL0nuMACH/th/1GDN3oWuNh+zdcPGOLt68KPscgMnhebuBWx9
xYZu+dUQykTsBFNSSyGWRCMpRCxYLdOxTdkN7irdmtXX2J4hVxAToFSO2Jqh1y+J6EWTklavj3w7
dEsbL5rOohgwHQgZ9SEoSLmgrVdIpudYt5KIn9zhB+DQ2a5MVakr1kbaeqGgPtW7j7il6HXHYnit
mcU9plbmGRTny9ERXOfydfaFHlrjeM3pbRbvwLqq1jsiE5Kmx2zVzPnexsLIeaj01NMZ3gHb7Dwe
m7T+lYsdsfkk2CiqO9i0RQqZH260SdNvTb4ObL2+5lvP73LlsqxSW6uFzmYgCujKgv88W9SPa4qx
J5TneyeHoW5t3mnzTWFCursfSrjviKKmWZDQ5RET7EvKjsahGPAGWc+0GAwzBh+XEh0ExxGQXQBr
2i1J3jDeFGEX2G7tRCzZ8dgs1rglVVpvljq1VMMqLzEKWtxLLL/nJIgtUkyB7QbtNS9IyLJ3UJzB
sbcL4OctDFmL9BkFidB2Pwr58g6NBv7sHsGyug2P7CC3a2DOqxRA3wWpTPU9jgJvxLJerCz84Oiw
/QeNYXR/mvKoT6Eb6/2AN0zHctZXk0QO29GpA1JIXFZZBVvbkrIRhr+zOTeMQnhvEU/Uu+BMbCzL
MpZCtK5gqdWQ9bbUrpOy1v/NEib+IuKKhC80SH3qdRNtO6k/RIMoVdR3ABwV0DsPwvmSkOMy6q8A
nIIwq8yhCHSP5r+n8TOzET3quacsrZcXrPkgu6h2kmrTqS1MidVgEXu5bwrBn7acuI2HWv1BZDSN
Zp6SRdhN3mshMXPI09djtxZ4+1GTYJNMludbH/kpVkeqIULdGG7GGiRoVsDGMVf/wWJvR7WNY/K5
ekGlLa7HjBN2LpPQelMLuRcWthRXATZwNfvQHpxgJMpN2KgMxXxc+qLuxHc7PFROMm5k4T2zVWWD
bcR0i2ieM+7Kb3p/7taidr4x3zWHflQgicdwXiDDMSduU/N0vnGoG40v8L7WfdWcQ5lQ1qR+gniF
7Z9/V4AE++70v0bLK/PxfU94vdbDrxpvt27nOWeBxR5tzyenmoyaUcWNkDuYpye82Qvu7QEj/tSL
m4f8ekoEDpjjgL7ucZCv+++ZbTtsX2fTMuQAvpGBwsMIZY2hRfiGo0iRUmdIA8ZcntxWim2fkzXK
83R/l24dByi25pRsB1P9NpkpFn0jEemJmg5V2kagdPWHtdV3dKfcrpo+fGQohsZ70K5mmrWJsnyZ
wOweX1RfDhPySVz243emuIONd93UxT0nvzQoNM4BRu0X0GNoT1o0cAp+t0IDBPcTEe5A9iiiO7oP
/k/kCse1hOLxZf/s4bXpL8IhHmhdSwY8/3O6pWGgF6b5ExMKe0oZxD48N0B22aIw2IQmtyIx4ZQW
iwks2FgI5Rllg5NZAH7dYovAg6yoXDwTKGNsiH6MrOL+Y9ukfoDw/saPF64U7PKfpkDTxuYwnHC/
d98MJLDVWbufcSktnmVgB2RjUudZkzYi7qP8hK/zoK5fO1A7Snf+mW4uAkO7LFWp4N2i2H7nGfsu
LBW8ccnKYF4ohCcviymuPEWL8daL9YWWsCtiVEK6AVFxq0IgZOqmQNiHU7Ci+DUMSioYOH9Wy+dp
lEjlhT4dp68AMBS6qM2Lx92fyjv15NYA6tdFjIaIuanEbo61wEZ+IvvXB+KyO7xiMMitO+lmNAaV
fv6RahLAJUu9xWWF6B78zf7SOW1iHS2HDYtXFaooVhY/SjA4fPiaNOcYJBn0ZmZySTI8K+JieGMS
BK11CQTfsQGhGL3qPZgeqhMq3OJ1Smzser0VlKCMohGoetmlJ/Vw8hFjuFTUeNhZ+AdvgsNcsQ7u
lNToTzFN7BaCbKwnqXZ6PdKpqd8fEeyCfVSNtuRevoKD+QmvCCzjZaFukzJP9w4ObEE5WVgKGYYa
f6RAHOdaWj6/vBNEbB1ohYLZf6W6c9hlF+Q43RwCyOSCaiMKFakkyxbceGpEsE2s2TR8rTUEpvGW
HtRrQ/9EeAVVzCgK00cNFAuuTDbO6HIij3mJez1uG0lAksqQNjAgcrT1iEqosC/m3AvEBBjfXzuI
bY6eWsCNFkZ+XlbOpwjT64ioyVQUfjE3MQMc8IvXCq6NnfGbOLiZC6HXZmm7pXmHAGj4wbEHLPvm
h8zDRMmbHBl3ISPDkimDdwoOYuvwEKTKvOCxqRx9FlCEoHuzM67Mg6YknW8WnU491QH/L7mEHyGx
nop+xpEZ/O/Sj6aCIeZuOTE2j/83KrqtlguP+QFwGWN6K7jDepspkiKoVX83oSJj8bVbh1BRNnn8
Ul9MTMxQiy3M6IEQMSR7c2DrOTpX8fFTot22T8kh4YVr8qAnzjcRnNQ1M4L4BrbxFw8Z/9wBMwPZ
jX2M3pLb517H0DKEPiNZET71bDnuqTdBBJ43zhfTC0fCp7OnIVgBnJeFm0CpTEiRTuw63HhCONbz
alZz5NImxRxKGuKv4SFba0w7zI0uuw9LMjBRJOUakrUbJFxACaHzx7bIIf03I5gStjnP/AG/vfBp
PdfyjDwcbskKab81vI6C3TS+RaIzN6+HrEsodHPF8fBLyYQX6xFLu9qDmUMHxSdL9YBEJBbOPB4N
meAkC13lS77dkoh4y+p+XCkPY8stpfvWj7O6XZwfXKsKx4GQgw98OkR8b+lxv2JKTGFgpxvwFEU8
FwvtTXDrdHfiOut3dohYOcqL8VjI+KiNUt1yP2v/ZLaBXWV0IV7pBKNI+jjb6HQ7WgqDuFfSydpI
fZLVPwNeVlD30NuNcHt2VVbvyP32PWFNQ6vpEF72/GpYZJjpEKrte3WVGpcxQTRm32U4pNL7SnLp
EPgBW8TI5+jd021TFVH1QwX2gjk1sW1b0+tVA5049KAwcSQyhfWe3Z2NFhYQ9L9YVT/QI9I2pz3d
SMkUFWwu4FZ/VG8QWgD3Df2bmUyK52g/dgZWXNBOiuPovx6rY10s31TR9Q8zkCAcMqc/S7p9O4dJ
POkiYwbVq0mtr3UmSRZr79q8hSjWx/reephKDahpr1ttIXF1zi8ydH6rfOHQYD9luTOzdQr70gIK
qtXOkfjqp0q77Oe8v12gvoNP/2F4Rr0pXeOT3i8M8MwwgIbCcL3CDaMBfbV5kt8CDsDlew2HLnIK
PayFiud+lq9xM/oljkp6rm5KHUVb6+D6+Brt47DqEj0zm+dbrxCdsv7nSETddXTVV0Ws9W6nucZb
Nrj26vkCAcqQEjMmYW25hz13Yoo2PbkdoCwWIWDMIH7j0WWgurXqcIvOe6ZlDEkz/KoFqp2Ogqo6
TdUDTArGfxU6xG8BwzpK86KqoGrKR0VG++JqLY5JC0KgfJUt1FYoHxZpBlidJvl8ZXl1SjIT0Osw
TD0gR2xXXnPSBMgZvrgLwlIzz9C52Fr2R950F7ILualD66hHxibIeVn6W9D2t9CgBRjakHFI6PKL
ZGylK4OD3IkGm1cM6BEfEnv2kY6DJdGvg47Kg8VvS0SeRMGFW4NamVeFoHGUGHDS6EowC9AR8pa8
sxJPGpFAr5pCLzQL4yaZ1J5TssDH01smPHK15x9MvORxPlkAtye4XX7ZEbfrryrg16QgWFchXtS/
H10j8JhcEu9x6MEsdZ9PNul91R67Mgn8a25O5kHXIMtfSvIapGJjT3W6dHWRYSti1l2fAL4OeMqA
CfDrcB9VkkV2ZvGb/62NOgH+qS6hCED2yxmyk9l8FSfNoLzWEYpEqQN7a/se+s91XmXgYFsRN3T3
nuB2OnuJP2yzzmzb+Gew0rLGxPcHxdPxxEi8ShOWnKRKoP8FZnGdSyUGru8jVSVv//CqE7/xYxYy
fjm9UHbDHLpovIBr5IBllIDRrxUvqabj6GZo4tdGB6TrU/myECL2Zn2BTG/8iYGTMy//bIJPniKV
lYEiRKsbM5CXVoXEeb8uCNn0s5qEexy/0SVzre98lNyDSBOm6vHp5dZ8o5Eu+SyKllJ8iCP0YETE
5nMgx6C0s7jh6EcO1pywT0QnmLEJVbKS3UEf4YNFJZVnHFaLR34qyqYOYlCD20ca0UyjNfprPwR0
Xd7/9WH4PqYxccGjuscjMuFq/LXUv/3XJ5i/goliKmRDFWR5oDbn85nI9TV5d29idlGabZL57gmQ
jc62S3onYBmZbfzt8V5aUSy9UoapbIgVNtDdLlnHncaueUbAKKHFuwGfTdfUKQaYa/tPpDNowevq
Gs9ahcGNcU2o45ZY6+e5csE3eRWde+MSX2j07w/cbapTphPZebUgeaRMspClpdzJOJA7E/UBpTP9
94+ftW4kEiNnzBlNzQggRzHNfp5TB7JoxxFiSACqD8dtURrpJSSWRxR644hkZ0tCy/kSwSByGb53
762iX/Vo8AqmAN99yDc/CAXf3Tu7h1yMFkdkR+jtwzMBiOcWTsW/EhBX1KlzTcLOnCJzVipKXSzj
NwNWdaHdSz+TCxYlRE0+CtCmacgMsW2ZZiG3AGpcZ++HyvdrDEotHgvOelneNWIW1WRVMCAStSeD
A8MU1sp1XuOnJQshl+oBJozlaPRtOCWWzXqUDtRtxlN6QxatyJo75wOwiRVyOPL6M1zenSQIHQtw
5yiE95podq+fvD0hDz1QO7+Mx475UOvsgM1Z2JuB8d0Vi9PCtCLxkoKelqyoYBPdgWDNHCoFocqM
I/6rC58hsshIIs37ffWnZu+nM4MSR75KVdQHzlfRKE/GkUad8056vfM3wceoIyEqZ0S2ArSK3ldD
ney2swl1fNSod31GWV+FmiULnzP7ktAHWhjqYiNRUFnblWLRHvUasFMmxToMzYcKo0td/qEyigDa
YON0WaGUVfPiC0EqZLqQcoT0pUUHmCk5NaW2O9Ec3KWUUrbBP9VWRdY48YY5y/J89JsnWpr1vRVV
uaSSSeU4vnk/zGcapp6uxalF5X3akLO24KtKDvGJKRRP/zCumCE4Oc4XwNJM+hX+U5ch7mfaIhgq
vvo8GpaGx1nkdDTnDwgzkzecT/ndw74LczsoEBHE8jgyErjOMpC5UYcZFJoOe1yw61w+J7WI/kyZ
U0OHtQBsybk9E/PmuOP7c4WD67q8zCbHwoW5nYuL2cZunr8b19ooyfdx6NmOFOHVNDwbXbNmNkCk
wHq8JjZKMuqgWgW3O4DBELNBjn7YlYunQjsOOGKwpZ9edzmNYqCNXwcb/JU6ZLKUcdsuXlUo1fuU
YI+hnLO62MmAjrPJFmWLqakpUBurdjPnJmoFi8bjDlIX5LcN25sIfcVnkOOZmeYSuCPmW4V8ShZ3
Zh3oLY4afyza7Z9+JCFmE5nhttEGXxwUNF+P2MclbyinL5ENdRlDLgBodHfDyk6W76CaFjV7DzFR
9SXBpaAQ8c+ijeHzrw1oNW0X6XXUibV5Ifr2yFS/gJNw2p9bYLIkYlwjjUM/TlTSX24lm2UVls2m
m5SsiC8sqMdcpiLvJoMEQxLz4u0XAsVLZmnoFjHD5jjMtepfhbdilT9ydKvjzMZf6FlLAGYRZUTu
vnEisEZz2oLkWfbByasgi3DTysiju9JzjZ/DaIuBjTbELv0HkETH1q9gkIuFO9cNev7L0M7orI48
d2BFwGuhOMm4CMadfbPSkublNxexQNSSS8utnuCzIQe1S4Dh0LEyVIN70xtRCSvXinoYEakTkdRn
3ImjRXUdvPs242Bq4jDaanUBgdN9/G3RG13yJrSgF07nlgFhQnK/SS0laxskElwakDgFrkbWXRNN
/jOWl9WMm4AB4+B2JPCO5X5CdmcwSGN+IpSYBV44ePEifiF5SVvENDxhAhmmARHjV3BQDZpn40fG
AWREGh2qbTMXZFYCLzhERUQJi6xGu+4L8jnQ88Fxa9pAieSjHaWSlh2PnpK/TnnIPsxAobzDmVvy
ALur89kHo3AScMuH7htsq4eunzXdW3Jq3FalZHTDPyWjQf1ICwYrZ9FdI7paxXI77n/HDAX1aRvF
9a8KyqEMPvPjRCfrgxUfA6MYcjPZElu2KCqojr0kwZ58Bh1UqDIdLtMtBtUIC5nnquY/7284hUCD
YkUBeF7r0Ve97Co+eQwMNd3BlCnYj3sRVQLx1GLRAwrEqnr179VTKhAGCtsbBx76Zy6EMaNAy5Bd
POp3cHqY2EatQ7rw/gdYfADl2aLauifg0JQ9Mtk5OFKJtHaxYFFsmcsB7g9T+CIyy5gEmkHbHZCy
dnLPccA7TycnM+CnwJ7U5ig242KkCh7IU5tjk7Tolm1tcv1qsmsQoY8/PDn7M0KUOtGk1bcAtsIT
OmgICJgDqpFvYZTOuuEbHki8LRlovA3e7BmeiXDxiNPvB7M40ARKST+VauT4Y0Kecadt+dmOXDiY
nnsqfDCaVOnAnzNgUYHi+iHDfQtwzTE5S38E/ifG53t83XWTdKsxAcwpJiWCR44V0oQtUGuEJff7
ZVUUhBxPuAR7WyNaBfjfruQisp53xa0Q3oTfiofxCWidkPo248VEuD6/d2mnkb1HXg7slowzfeMN
dQu1b3n35hxbZDuXQwGby7f5MkxrqQ513pxntAyNOThVL8doKLPEXChX/vkfvX9ynpztSAyImYSu
lEniqbvpLMdgej1dVDFlOHUM73biED7LryESTNimSvFtwLZA+ADHTU5OBl05PA5b67ZoQElenpHB
9CFzUiW5TM+UEjF9ko/xPyG6KswnvJihcjz9DRTe92/fnAAkg8wVN8jADS136HZfeoUiS/WnPnJP
E5HQ+LfyGwrxuH+xZ3aj5JF33fIlEnyqzMqSpjAdYplQS6ivun5IVRcWnSoVx5E9kI7+7OgDJ7XC
LekwgoGhBntdoM4er8zMXxk8DtTDFOjC8/C2/uc9HPWvfxwXEz+yp69GxmBQHmX3kFA+ZT8t519q
kvC3WRht3vHu8+TgGJ1Men+oxw1N8C/VVRXTYUhqsHa5tqc+SBGrppKRoW0Uc6T8aVnn+k0a7PHj
Ch345hSvBl/NmiVLEVsu19FJoPpzSEOf7H8popQKpa0KgHH9GksCtxmad0m4ZSrciQe7ClZcacZo
6FrKWCpOMQbkFSoBDml7IlcbFhddRZZzvmjLs/FUHcdaPzLrLGJX7bW2cAzx3C9Q0x7deAeXVO33
Qqn1vTZpt8Ka+Med9/jxGa4vF71hasGenyyPZeeFmLE/qu4PuksNJ4CYafbWRgv1k4z1zh2j9esq
GV0dvsjYGPBb6WtxtDUcqirl76KGPv6Z1xER4hm+InIRdedCxIuFaMfeJ6uxibLLWBz7mvZ3fQ6i
PeRNzi/e2BFWzB9pSRRXGrJYzOXEbZITVDBtZrRHLfjq/sc4c51xB7qENyXLQjhCeyZybF9eTaww
vVA6ubR8IM7HJPBv3TbUj/IDLXKCynef+WqpfkeqiUTBJ8MmfrlStwq/uolBfpbHuGord39s0aGR
HYL5gb7VwvUV/Rwz7TuZaFbjtoD+0TnGTWIsitSNv9tRDPc0F7+xOOijpt5/ySq0vtKEf+MlG907
hBiK4i1Zrlo9iYqJKvtV68BznsLpKQOp3A5Hcd1HsGSaHlu9eDAugw78HnK5Y9NVXaR1WYoNdTH3
AMvmZGt4ixovP2JLPZZoXgOLPEc/CPw1N/DSgYzVBaXLZxFKviIUSgQXkSMxa33c8uitNT7F/Cnj
gkJuld3nBQTSRcXvHg3upSd5UCwLkuGDCqwF05hYmNsqWDrYDJ5lYbWK9ZmLTrQNWBtDV9+DoXOA
HETauP1xOzjEhfrNhIQdBtDlYT29vzZJRrkzSP/lFeDnZMo0b0NkJtYAUgMWIymI4GcCXIBGatsr
jEKDAeUAx+HbKaAfcENS4ZS2p6YshebLrPK27oqZb9HsEEQZBJYMlkceHRq0LWe3xq87/BlMR13f
ILOc2xJ69ZLZL2BGv0KGU3ILu0ecczNTEak/2ISxsy28po3ZeZ42z08tPxlbf+OEJnX4LCLmUVSa
BfhgEfnNL4jwdBBcx4lou/zbNqm5UfdLNaVEPqmEE9Rfd1JoQjR3hpQDnUg5EadrDFW+VZf7a74X
7z8zMdZ5kTs24EcFd1uwunrrxrz5fpUd4vnNXn83/e6Xtc2x19QDYH7ir7stZO2pj7JmI/0RokdR
sSj7UMkfr7WyrovCE/X4kq9K2XLQVSixJ4P7wehEPQbs8SM0hF4Nsu+2Ak9XBiwJA2vdjitakCz/
RJM5PSq7W29E+9/6uL17AdNV3Dby163e59PSKStlfF0ngIGT5F5OoDH3HAH2MpWzqqPqoz+CaDsC
kK3VGI0vpvSWwp+spCJcYfvaixvoKCASyh0wO0b7I6As60NrqPNO3gpilr07nHvdr9njtyFwhUAO
CCxsqs+kUh5BfRqHHx6wrxqeKiI3GRzuadmOkEe4x3DCtgC37hWGYeMMwPokLh9FcxKciLzeChNJ
1Ng9yN8HUfWnMFCT59oZFof0SaqlAwa25UgYsN0SLgZYfftocY22vUYMvSy7sa0RndQXb0onor/U
/KGOL0x+hZx6XlKF7U1h2P/+2FK4qswMZ8URPbPxTWCiDVbcQQnpvzEMb412pvnlJBjhmdURyV7k
x987dkwA1puvVu0062v0e//rZbjv8EQOBKL9L6O9BNM1rQSYiW2siqTPx3URoS8yGtW5kGRwhtTe
VeC/tyughJi4AfueJ9v9JEezyB6QD1eeDFW7YFNGz9QQD+/BdqQ1efjwfmOpA2uJ1pFBVmPV8hqq
oikWhiXr52kgD+XbONsrpIYdg3t9ZU568S2EzDMLItuexKOAPizQ7XF8HlsVfqX351T57mSyG68r
nUaL55fRjd1RR+ym6qyu30DU/BayVpIl2j9M1lsn2TujpbfKM+xkjP3ZJIcSEFv9j1+Jw2sMrmiH
9EGrA5zL1gra7qUZXObXRsVWvfBEuX+h2WR15OLt4almBkvLvKvv7sTAIs1BXWeOOWeXEaVO8Hsc
/2ATZCdntQlIVSlcawtFy835hL7M+f6jfd4TkIxH790R6dTwd6ACXO0pgrC3kL39JTreB41+En11
CoKPgIAsn3YMiyTD6A//SSUhpPPc1LlvqadTbMhyXf7T2p9O+E4o2VN2XYN6GL9FdwvRyWjN8o0l
Jg1E5g2M1Xvy4xdXbkPLnkHOPGZSNm+wvIaQOKyTecOw+C2FTJtmDGyvjhkpIW2pqhlUN1KqhxgI
rc6b7KEdy/2aVDNso1MrIsPoAE2Eee/JqkPc4jkViZjivLBvBnAwP0TWei4fSnd8qPcYrynOBI/9
h0VqyJQ2T3FmtCdbVd8A2QZPjDh9siOsX81qyaK8YvcJ8WoohwYxXNVYhb8Nn6VujTeTxYDrlR9o
6ZHpWWCwFeb4R4sqWIXHcdbdb/hgsxKxD6mLIaw5BMeN9xOF36ZC3fOSZg4rJiYhLZdQZMK9TNJQ
GgPtFrZ8WNx2MUnpPYH5qjPlM0xeZBxCcVeP+Vqva6o5LjzE3Laz6Re/fNbjhIuvazKOgaJFBHd3
xsPUY5xayDXck6JTmvsNd9zTE9Rt60u848JcNmrLuum/YCIKqH3lCgXgQ3wzp5nMe5I9ohJNBOCr
yL/jhK2PUwZJtuzZ+oPupZsgpA9cUvyt0Cw2xBAZ4fvUkUbM2iB/9b3NSvcHJ2qQT4ooiwAlG1BA
OaRD3U0cF5aFhheyzfpJqfH9wTBOrn7+tUE/sBQi0rPsf7nmdebrNBTS+N56EYQ5ViCOneT73E0y
zn0SCJRZK8Di0dyuJ0uKJhIxREY86RUenvs1sK2uPbUfkVw2QE0JBXBG7QqKcY7RjtD3EezMNiBc
weRMEiEO3zSutltd2Y9rIFqXVaeSdnY2B+sQw+fLmvby0NQ1hIanNMCg+U2B7Lizc8eOq/MF9hWk
5nEF0pIjT2q0XRQFc4PQtxLGdiDMgEFHwOXNV9QJ/6DgUYuCz4PMc8z4XYTFtOB081akPime6NOm
w0R90ogFV9vUVeEoAq+JpKnBRQ9OFi0IaQF+6GiLg8ss/5GcJbURAp5CgbQHJV+HOrKSeKWpldIV
da3VEAVNAvLgD8oPJ345OfF2V1PcP+LcyhXcPSNo8/+GxAdlp2uzmgII1iYlPidVHYGuon3SdBYC
Y1jec3b+ZWM8pbZAksiVQLWJmPfcNdaaY2Lq+NERcvQtEZqVxquiH0Jbv59wVEeRu9sw1pUX3+fk
b4WV6OP5g11mUsR1D8AE2fD+KYzzCGJJWwD37oE9V3a+8fSEZp/24Oew1kWuUDbYlqSVYdxo5NYR
Brvt7evrrih1MSCsj5qQ+nSMn/zQp85T3wXNQN0g3ueXIEqWDbsI2psEndoSCPJ1C2zq6m5hbeXL
26b0YHdSHGQShTfXA3MLoOfikQFCEplNb1utBDRqEoW7/f22QIJHqEb3DnzDI5BI+m80aNqjVCxm
GkQ3VkRAiQKHBYRYp0BWg+JWYxDBnaZTHvMHSzccceGNvq1BuwUeIfI4z16p0xxVgLIKB5p9XD3s
gaustd4Rl2wiVQExg6QeAs9DdutmTucYo6FqVHIFbK/8D9B+FJ9yaeP6mgCsZsBemV2lFj9eXGC2
W3bnwcs5cHOFaVGATftDHLdmn16li65d34imz9l9zo9BMW0W+4qDx5Pt/J6BbauIVJhfxgc+JZLR
A67enGyJ4BFVecQmLT/0YU09hrsHFlloPcaFKOI9QzUleYknNz+Wo8ukkTvbXopfAfZsyZi8ihNd
A0SzzB1KiinUu08oYijl/WBGm/RuLod/SabShebs6xsBpT+KzP0wJppIzqBp8Gxx3HTy1jzBaKrt
veFM1IzrAE+dJNxgSvxdIhf0wzW7Mv666+I4aTtJ8dKKuzYJbYlwpZmAqGlbyal0Ht5pXTYiUB3e
2gGRXIrxR8VX+ezjwfRBqCtbTJ3M+ADGpw+lE8Z7QZsK0GJbncd2jeztvlx77sALixaT4G6LRn1b
av1S7UqLjojI0+tehYG8rSEofgCo7eOBDbiBYn8O5/ucevKGtdSuA9YOHraAPJDFEe6lZxZ8fY4l
jkbSKZHX52vPnfXKeseSaHszX7Mn/eStPBvE8Oy/il38KRQvoxygV/yF8UH/pHrASd/aXEKqx86M
8q+PYjw/iFS4B1KKmU2y3VrJ+D7etALeb4i26NskCayorYPYX2d2XgWosqyFUulkyAAawN3tzddF
065j9EzcFNCmJv7s5r6Y/zgulGBQTIal1vud55Qv0zFtVZhU9OlegZ6L4aeGZXAh4xwDuZ/wfi+6
iAmGXDTviffJJqOoLIC6vly9ySkjhAGqxJ2OERGVYsk3q0Ud5zmhHq8thgMspwI1/Zr5nenUW+LC
NrUPA713okeQe08sJRjO4tLs276yuvya04tQ4bzbaqtJc0JvMSzjnkqDNvx1R4fXxpCUBt1g3r0k
ZNu48219MGLHNQsLXx4Dp+PllcWfxq/myHoOrAHVt7pqJgZH55VXtbA5x6WwDu3svwlUBQgWH31d
EoABZP1PnYL7lZOi1jCp+0S1MiPGW6gqcC3Uo3NyjumA9031ibi1OzjExj0gb/SiIRJrPbVMVL6x
/e23WbkWXiN1N+eOc+F57mZ/XzyCg4oxCQe2expkCK0y2BZckJe60BVirsbMDVf8k/sYXOH45ZIV
hVBTJ70RJZHuHmDwcXQLY1NQb/aKFINUCt5SxkgAcCrCHh1EphLAtcAVdNzSLIJQMGoKi8WL7gFn
62QAdQQJ2Ixh0CULpPr9DHKH0lZlo3vG0v5Sn71CDAiOzGuPSKVFTtQ8KAi/v4XKoVwgqRe2Hlbh
5Nj3JOnzPvA3fk6JjfM5N1+iQG3iEpdrsl9zzhLcbAzNZ6svPkyT73Muxa6eGHiE0kfX8xRRziRA
nMLgtzXpWH3xeCW3SfTqtY/0qv535gGn4k9gztQv93lzbCjiu1YHVTvGea5d3Adb2YVcd/J849bQ
DjaVhXmB/KVOL2Q2uj8KO09N2rEFL5KlV7WuriCXS5YduK+bV0KezH9T4oIMz41m4UOB783Jg0WC
TeWb8H0xJCBJb8BajVo6f2TcaIpf5M9rdLmXXGO/aZmDG5h5+doS0zpE6D2tMLQB7QgU1GDDSKqh
RP4pCiiSBqx0wUGpSj1dCCu4nCd0LPosS5a+1VV+HD+uP19AJH4gb3M7+Jkl2fYBiIlA1fLxFW4T
z5V+DHtyvQm3qSNwoidahSgcY9pWvdaH4YuNeAgY3knzLkb415ZKWEkqaVk1dYUIfITJfQ4NhDA3
1zbXaQl06hTfCcCvQk/f62eqNiBvz/zHGG6PXrVDfSYbJhgdvpTh8twnqNLfZjiePgFPXBt991k4
vGvKM1if3H9QHUjhmvjyFs4M3TiHtHqj5IQKSztfJeHThBC99juU1fTkRcpKj76dY2Dzgo2x+rSX
XiNr8di38aDb+iJL0bpRUE0dcnbWZzXLxR7gIRRQIaB5hDvSOPGhcpxt3htG+gifPKdJuW3oCrDH
G3EJkF4UBLpjqpqPmKxsJI6/x/I9iykMRKzZcJvpnA652GnuQmtMU/SGWKwPGBreYL4ALKMWF/7K
KkNtnF6LJgXalh34toO4aeBxfm2FoUM1oZyyDb8LRUN5crOaRLTTsR6HC700VYJAASNdfHCZuRH0
9esF+IN1tjrjzW5b/MKPW9Jh7K9U32clVtvvnTtnZv+xTM5C5bmPzdWpC6b2MKssDWoWVql3TmpO
Ocb1RYn6nq7iDJBY9/U+S+nchoNlWgczw5XTXAXzYQQIJQcZs97Gi7tEvUxAbjKd1BE23PcINcvu
Y2oS1Cp3ceQgW4kBlXpwbD0GV7oXV3THrJQ9YUaaZlEVK0X5QFOLvfcB5EIuzWGI2H6vVFfCeC9z
4C/roDjllqF7B5GVkRE9ebK8CxBfhFHJ3TFsVJuU1L93kCvEhNgvr7iV5+4mh6JFtETm7yfJqOTm
+8tdERqmL8xpeNzaGak8xIzTLoPGDMDcUSg5mZHaKsJm2xsztJq+lMqWF05kzYsSWgfJhhf1bS6F
HUbA7RMiTpePTpU0nMaFY/7iselvnnjrkdJPAPp0kdcv7MOLhUPrkDKPCYbTZW3IryZ1LfV9+XgA
x+pdVhUFjdqWMmkxzxUA6BEXV6dgWv+/1RQ/NYOKbKfYvG6eakKt01CHQ+I7oInhJ1Wla0Dgrd8c
d9y5+grL4pRaVq21qBtftzkDmUmVFLZC22uCkCnvmLTQTBNZMPNm/tmDDrbL8Nu25e8KImrcXTsR
UQWatK7VsrMxYFjSMINMlrui6Zei0UiInsJiuChJfC+6Q2H7pgUIYOqsg1SD2klJZ4kv1QrIASyD
3b6ABvQmiDBU0iMYLJbOxxoAAEz8lbvRS4HN/Ue8ixLwbuLveHY5TpvAd1hfMEdzlC8YPWe4jjuF
u3DTpQqcCX/TPE33x+mHV9aCt1apKrA4rEKv8c+WDB5HgynBZmTrVjN3SsVAVgLLgNDY0pMNJ01d
GlysT2ru2nTklUHsZfCmI13DieJ7k4jgkS9ZI73Gl781xe4u/yf89nIAYWrUDxgQAIVJikOxdEJW
1ZBAUXzxcZkS1oz82LIKt8/ZpigPyUyjMm3jNL8skj10MjyCni0ettR+o91uCslPzkSEE3U6Y0E9
fAzyKHgLnxEIgCOXlmTXs+IrJagAyodUCf1fpgFZE0U1M7RiRMObeA4GjjdTviW3a1KH3+7mxE66
QLVi/WW3VaA2QjjK441VnPhnRfYoyBa+k87NzmUAKy5zrEY7jMhLVuN6IEf2R1VSXbHQFF9kcZXe
hKunwR5pBIjxx9OaKX4lscHPOxC+n8JrTf0/Y12/XHYv7hMiPCb2dYd98+zzmtEZn1oxXpSF4Oli
9ScsF8fZ13jbBMo5z+uQ99l3dXlEiVK/nxjuZBG2Ljzm6BZD+Qbw3r1nrtiggVLX5KSCbl/NYmJX
GmkG4HuCk6r9mxc60fEI4hYlCt9CDokiPTRKx9v7XUrRh9kiSqg2psru4KUhNlyyL0NMc9Ul9Umd
D9Q2pAFcfvpeaKHM5BpLHocH5z9QVoM6e+OJE5l8fr0W3rSBBx1lgVvLt+Fzjyl3cNxlSvzZB0iW
7gh+vU3dK+FEZXTc4nUrPQ0EMPX6NCk/yHgVNREy7Jfw4xjAnKfh5UQdaOG+N4o7ZFRSqfYYMUik
WEBpFMXoEYMcaYzJo3bWkPMTh3PDRJ6F0Yx6N0ggkGKpqSQt4w3A2Ps7umO6iwGANxfkP/IOne6M
Uvqx57CFHvFOJL0vSMJ2eSz/IqH845fsbzGm+PkVD7y9PyGvdI+XDe8OWNYnPRP1EQYXyDbRfKv7
SoohKnMSqhm0jb5tR3+09DnH36WnZp266RC7Gvkv99Gpl8RtybPRDjuC1rsaSWoxUdDc7PL2PHx6
sQzZfmG2Ck1zUK4oLyZuiNwTS9uwTJ4lXrVxK9n6i/7p32ex8nAjOlk2QfxMIaxWi4ZSyrZCJ4Ys
kIrXimub1JCMwwxRpKNEe05ylVZHdNpR7YlUuI/vXMrDJrXg9xWCJ98XqXrC50otBk+hUM81wAJt
W+/NJQJX4uvHr8rWj+uKzlsDUzB2Zi0c8M3sMCd7EKdKr/WL4Lm7I1mmUeFzkbTX2tv0C3DQN6ke
Y1y4lDlQR6fRhgI89K6wqFHsuXSDH/DfxBy2ECeQvI+q6U0l+I1Lg7Kjnz7Ga0yWEcDfMNMztsOM
ze7bG9sXhMnJWx1TUNib7ufaPzEBXy8PuQV8mtlMsGc4GgGeMBgW5S4rDMruNBmIILC/+hgeoBki
L9cJ0mdB4gHQiP+rM/uNaNNAUwEZnBcC1UzKtFOzQaL7eML2s/5XP8+c7ZgzhJTs8Qk0OgesN0I8
CoW4nfXhGS/8A2/XCszw9Z7W4ZSUwHDD6jvKzb1QUzIHwKgINiQqWJ8skhGxVRIfO5PgIT+8h8VS
qE+BRJKbUwZPmxB+Jq2Tf1pssLT781Womx0xXj8nX1ygNyKoCinl+wxxeziwNz1QMW7sGT3rmxsw
zAbOhQJ4jZrMjUAVLRd77ldjOw3YaVE1s5z1PffarY9ce1ELS2oyGGuhCMq8CkTl7bSWJe/GEqRz
M7kzCNDzp7WRfDsEJfYwYhk2gMO6E4LseB10Mcf8Wm5SoDspJtl8/98OSZ8pV/tz4RU+uTV/yz1b
HMdvFeM4ioo2sklxwbLNlIO2DYwQ72eZStYKFZ5fSholCi4hmsmm9Typw4a/LIOXRLlvEzjeH0bA
9NFdOdk0ep7fae74QjHcX8JDFbAnZioOHTQjdk8Ow/IeU/uFyY9GLZl3+ZPYD9x2jDyCpFLNPNca
O9UQFAqMSM9dx3Kgsx/jD4tCKUQF02Zt6krxMf2aoPkbDyK27C6elBMHxExeJEQLLj/aN0QY8l3e
k8Pe3RToTFSLjekQvno0voN5bC99iBbfKEADKWswcnVwRGZoC5CDizdCnV0VrxrRBWE5I6outaro
oCIQHzpRJ+wNljxFTJSkY8E0XMQt0wfOrWylZtGTRt1Z9A18HdN+DKYcTH6+UgIx6uCElRfU8jcf
jXu0p0U6lEFO6u58GILshX1jPB60hlpP54HIY3aXmPeDB4/MKzaxCqCeNgsplLMl+ijtKoyegmCY
ojCIwB6ESXg7e1kA/tC9kDAEBjgKmnATI20NtoohIKNqfwpLUsbj55OHEBicCluKm7Sl8L1krFz5
dPnoyvKEmWNU2Q5L/ZwnJhm8aNSYwtrUDWzdFvTbvoKtcc4DNs+LSNfVvmfCIshiawUyoUD/ekHb
r/WKDIzrCeOWa7FSclNVYzzq8DvEkJrEjv9XfpYLX+Fc18UDHkndu71OF+tXRPadxYFlJmkRaR8D
YdyjpF1akzRIINSyFisTvemoWAIsAJmV4rnUkttmVODnUnc0PVc8UpIW8h6fwIju+u+qdDSASADU
+u8F1UXbp9ZWgdoODIkneHZgP48kKxxsG05zTjgh2UFy+j5AGnExRJdxpM7+NOEN2NGnkK9ec1jF
ftUmsxxxPmseeZne0Tk/Ss8+N0183eJ22kvpcksYtREvM4fwj73VogbiiOisWqXPvfQnL9H8AEh/
okj3v0Ll4m4zDoS8YRrur9HiR0C8cETBu+fr3HUuwastTLzZEaegv4/NONybpJVxs31obIxgiIFD
rFfs0jFrE3hezk2jyz7DJJmXkRuKPJw1lad7KbITHPj4DvtvQqZuPx7laC0bccdBYU6azRR17CMp
EVYZcs5ToeoesK6MtYKP9X/SZ5qvbMWmHvCFU99MMnQSDlw/lt+x8qUDeKypdMqfq6NSVB1vX+4o
SvuiB757BnOGeNVl+C91qfkaLlLslNpYk4/sUwJiAyBTgXyu+DgAs469SwdS/j7w3j9CXIP7XdnE
yTQhtytvSEFZo7wykoJx4TCB42xxdVq/zaPdOgcmu1uvvWJe2dVlOsazz1xuKVX6dJDlvmWJ194z
vT3jisRuslBkrxRT1kWBogNTsB9DiEVrNRCMI1txoWYHnRFlbA8ndL3yo5hRiOvU2wE47gIXdLNJ
tE9aTTHTpLFMJTD1nX3JOuLwlOSJwDxtp8YhcveKm/U8F/XjOt1s4WVrkiIQhem7EKYRupxvU6lB
Sp0cZo2FhsE7lAX6yIlAv9HHPFEOG8ukV357k3jyNaS8ilqxCGDCbS43McA6R/WpRqcL9HVWjAWo
vlctIzliHqdlouNmnoUSFN3/dsnzpUfnSbHFxd2fE/eWS1Hr9QNiqkJG0gOtUvHYV7MRRtGzZQV+
ZVJsWHKUEthMJdNAZLVZF1OJlGO8zJos203gtjUHOSg2036MsQWIISrqtMQVkSVvv4gtqWg/4UzX
EGVXWwTWni5v0E5+KiEIUQxWse1kLox76o/35c/b6d+jA7hCRSfLjaiUD1vPFArJxZjwpQoVp0gV
5saytmIZXeMs0grf06/hGV4NtP+stCPRQ51l9aGXzOVyddW9xsFrzb+DV7QXD6iyvOnFeDNqvJAc
J9FrpVPjgTzreTXL+PLrninNOjEQplzGC+2d584hgak2NYSaStuk1twpTE43S1O5I7k6vZSTkKUV
UzgDG3Eino8DUvkS4gb0/lUB90b7WzaNHSlfcRBjYKRNYbn4y4H+SmAoBNny3uQQ8/zXfJpjQ8a8
eR66FjrKwP7QlHCXfjz6AuBgBCNB8Eagr58T4FlX5tckHYX8u9e0rs7Lh7eHSC3plkv3YP6dUhV6
HCeDtPF3RNim0fq+pT0pSrejxpPvY1X8ClPaRX2VkUTiIAL603WdTDDpqxJB3e+stO2s7sFqbtrd
Ei0t7kLm52v47DXR27FUrmEFkzRucs7B9yY9U8G8Cnyapohu30cFs2opw4D9aKDhMRsf6uHTkHju
6YLCQG5cBl6eTMwbsKG5PgFGhsnfph6BUZgnuKnaXZrqtQefOxIwZEuiYueTDfuw64EOl+dFANKi
bbZC3KwuXoREgNQao6WI97iMwfsy+3yR+Do1CcYSK1FeGMhvzcX5zkNnHPHUUZW3yWR1xbAMP+C8
Fsz8Q67Oak8q1KUsTuc8D652Xgigz0Xf36wUIhaAbQlpVab7tnNHEYhYH76A0d7Cu8d+jRg7A7zm
cJjsFpZ0SmpPGbUPLlN/LBK6xP/cmcVKByIIqSQawSr1S7C8EYp5u67JSVF+QiiJwHNH+O6K9RBW
AJTRdK251cx7zPx6Z74KrLN6Ww04H680xdQrKjOEHpYX/0fG7dwaXcG9uy/dD03BgOiwf2+Hg4+x
XDOUK/+5YRGoU7cwupd3ePMsIhGvLJtehoj59vhDb3ac/nXfgLLqsOfOQDc2OGMqpmqp9H7BMJRY
+kZ3CISxhm9yiFWcxRZBHjpTq5ZSQ6DMkQyxGA/fyYKtawMBgqrJAH8mB1gP7zg1LCjC1PQ1QN2O
VsheKsp+h+l8+514J6tsXRcCWa5Tsz2IqJDncvhHvdr/kzBXhgY4kZj6kCRkTaJGbzgpIJ9nOlLp
iNUHHAs/zFNWrVnLAfkWkhkL3Fr8ZTAC+X37zbT6ommsqEo3k+73Q4+ts6GoNk1QFTAEtjrMMK+Z
pQzep3V4Y++eRS1/6bwyXkAmqgXKjvVDUXLRMNjmE0MY2IlhwHYv+A4z9fsp299GKgErcEfysS+i
LcvN8b77XIp5+mEdDFAqre6zsOlrUp4omDXX7F0sBrMPBc+1sDkpbbgaFSkyiBg417M/vjcFnrSR
MTD8GKYolpZJOXHh148q/wQXGZlkVLbefh73uYgm+rvnVhqmYfFZloivtKOqzRdAz2bI3zGJfUq/
MVDgspr92UtkZKXaVcR9T6s7Vak4H/IC+UorIT8c7Grl8rkG2ZLVOSn3fzp9S6cXrjFpaV5w5zwl
dU04jEbE7RrpcfsmjwVD7hq/nSLbByWhpVgrPuuF91vi/x57DYgTLtl0A1GiAHwau2siny1/Qw9d
jEru3JtU2KgKn4XQ9/0hLguM7EII+IGj3eIL7pT6j4TwSQCPvrLWQEv8UNqSQA8a8HOdvKHMAe6i
9wQgGzqk9Mb+8Zt2iJJospo8Pi147VGzkeHRFidkuueSIO+qZvoAKqzCJSEG8dbDymrJYcKK/nDM
5X4JFqWFf32I97q1lws72MB0s4iqDd6gvBzR623CvAhVdYytmqA87n0aa2HHIs5K1HUtxjXQY3M9
k7osIg/sHTXoqpyT2GqFi6iB6XFlIL0r2IFJJPq+DeksAt3MiE8CprWVpszw0lP+8zjvkw41PnG0
RXsb2CKSOqjJYZps9Z6rYxXW230Sc2vhlGZ+zXg8yueUwJzs3r2lMrvCVWu2c4sJ8ShvDCWdAlJK
nVHgRKswS0k2aLOhWeo1NA1iFK+NoPk5ca6stRGs5HFEOrNMHNCH5txgVoBr/EnRYmT18c6G8/04
RmQIqMOUkEwHXG1OC2rPK7LJXnhrmx/NVBa9skpFYef+HjNFS/rwngzoNR7uGlA9KqbmTQCOROPv
27G40PQ2RfXH9FwTt0Pq010Sr5wUHd8xN25b7Dd9sYhsccpChwJSLQlDAM1HnQSkVeleHR3xh56d
XrT1pJInx2uCWJDVsp0Fnigdc5H9+HlOTpPglFglG5/Rp3Rvd1IRs5flJmTgvsIPzlYwBUjHEpVV
VtWGDVAFYN0UHoVKCx2dd5O90bIHaZ1lpEdovl8cnUgNTBJigH4rvF2ku6aDAIFb4B6LSROyy8Ks
SqUWR4mDWTXLGpapYsop6CL1imXCNhH7yj1YMfOHmOhQICKm6GF2bs6XOXeyYPVu3a4t/kNyztpZ
TD7JDf8UJvFjX3uY1vmPihEWpAkIs172DmRPF9xGGiTsiVmVZ0edHXxSZqbYkR/c7/lSg4jGNxOH
C0KJSbVUQqLsRM8BjwD1cmo/re2pa+uymmtNv3oxW2is8Qe7sYQV7rQh5rg7Qg6/4pO8on0UKa6+
YeLYeH3IURSOaPD4e9dk5Gd6r9cEObeQ8NxI/bnimjnWurv4M9CPiIauuhhAGg1CjoJfuj3gS7Pv
NpuaDx19mEIxzSIOiT2m0sAX//usgADxYkNvjj8V4EpwmFqhQr6JSkgs+h17FfvoyOVp3gGsAzwe
VR2fEkLYCMMxxs7PCXvgF9yctu6YPUsnIKfbygjVo2J6ZZWm0hlytfVbTwpL0iPV6XWsplC8Vuix
TXVmofvlGp+5LfZ/+Y4Lz+9BPkisw4Nqfk7vzU6pw1aN9fWOQ8I6wp4xWQP4RJqj9slfmzDyAFyl
pXOCYJtcfRKwSoUq9qKfI4FcRDVdb/ExLLaVC4hckjMmaq8xio0JcM7cDCg5kfUAaCszmLFqxxjQ
gkioyPEfqKf7iH5+QcOYBxHp6g0MMZAJ8CZaoBPtFw89S8p2FK4nK3kv/Gonj3XMUUqUmYh9X6ju
gKBZIpVRJ0YMnch2HEvybNCwgaZaLWgG03ToT9mHTOFxoAmX7qCOnRSP/1ogb9uWKylbvTUsU1wZ
LF4Tu0u+CX38llvzZpjL+WAzUQfDHStRcz5ItHsbAN2llwdBc0+6V/okJuObx5e/DF8jt5XsFqOM
Tn9aGrsB/EndrPC0chcs39oCsgrXeUE4Ls1CH0Mq0LvNcX/A3vWa12ruz8jpi4AAU61EFoTtBlw6
iGlDqLq4E7mgiStR13hi26JMKlKoq0ecK/3w5FRos12XLUxMGsUuTwcTuRXi5YIK5zwGU7oP6uNk
+5N6UyU7ylfThdfQaEmsWlpyeCyoWs24YyQsCwJx3Xy6BLsFVpr+4bQxmqlf3M20cpeSyFyB0s0Z
A8zI1qp2VNk5CRnuj7L441ubehDwgoFN01AJw9md7dcHHQNlVk2VRicwGOPV5gD/fDE6hv1u9Hm3
ujH9E4tPWW9fnvTGcLC5850B+b8zf2sl48lO8f5cTD8317K/z0RzefWGNBKrP1J+CMLySiooBA0f
vijrSuH2gSrx8rvxduoPS2Nes4dRStdT5HZJ1O6FCEFwCXJLYhLLMmaXl2tvWoG2dF4nZLTKwUel
HLbAxAH8H+RzyrRfJB3JTuc6V4+S510AmXhdI/3WKIz8FbFFJvxs9cp3MMklw4ZmxJo3K5rNoToX
2LbfaTt0ozlECahejBdjF1+cS7UYEZplRBSZx0mqhGUWOrs3O2LXC/vDwI8iYAryHrw9GD4BLwWX
1UYqAyT8Sg1wuNq1PrWtzLKpNlC9ZSZ14FWXuDg7P3PtL1Bnr7FtxpYDIL9HF8HGRv0b2VLS2rE1
Krhqe52GTwEwnJQc5oXugP5FdAKCDWU7q7Dof7Y9LFp1aZvOnKdEs2NVhGUARYyzMKmkRpvAsj+C
/E16/O0JbmxVIp3iPLtpAHc2fnpDmv2jn6+EJFCtsXX/k1Yj50qTrOBBZ6YcgiYe/lwnMSCr0GoM
dt4W/ffnsTnKuXbYobSxZ9rNJpIpn/aEcZYdmicps5BJW3rXuVYlAKigJ4XXjKj6qIW8myliTl0p
IgJJb3YG62FMoTwhvNKzztKHqbB042xHMU7boLOYJUuWgldWzmAt5/nUgg7hGOLddKsZuVEEtCja
oye+CSb06C8kD/Mauk36xjUTKDdHQeDlu23LPQecw0+zCcuh0803XiTxOrBIXDmqtxX6fZ2vz4y0
pZ4q+p1GdHFPYVd71aGoTnEcECx6c34HHKh2uXsTDGeI+PaSP5xzbGSl/6nj/8WwaXS1KT3OOGun
GvzOuHo9FX7o60ZotKQm+jUWw3vWSjBxsUvaZs7gWH9QHgZzvs2F5bUrkRG5Uy5HED5mKVMwoo2d
3WTHHuDNolCrfPT+XNK2p8v2Mden0MdCUgOgACccQ0e5Q7QVhz0MEjO3m45CYmaS38B7yb6HK9HJ
sjdq6clwdkzgBjFy5uAUihZkvy3TcSTsIKTM+Wzn+wcRSEeuUTNTXp1IdPj/YlEeeqZUdUhZaDaJ
UgMXNl4MM4P/CK44IYFmW4yY7Mjjp44YZm6sx7aPmxRZODRfplcAHLHy94dkqJkOT9wSnCEltQ/6
yaxVlS7rf1EYvzLf/TOBVJokPlaAzyMv43e96bXq+u0kn8anlSQ0g38/EAG9FN3QfO2c48HLp3gI
KUTXDLPst1fjjmJoSvtvzNlT8WZM35k1yWZ7CSxwTcFPmBG78YuIL5q17cIsdcssPuLAiCqWEr05
PgrZnUFfKEa1LDzFbu/emQ0dRMi+FljoizqWhOprILhxTsLnc87Gpe3iusRp/Tos3O2ws3tG8aVP
7/0kL50qU0ol1jCXWzJIXo0wad6uatknnXMLcwP/q/0mU3sh9H58j9Af2Olfocjq0sHseM548Lsi
aWfRq1arAt6C2DD1nwTDfnat1hBIdoZyTr09DdvOLFnYKg8fZhVwvxtRPyEBV+nAnlqYWHu0E0x2
QKh79o5gsKza/Om5HKxXhegGcGwceXWF9cy6QdTGm8xPENzqz8FlD344zdpVmEA1be1gL0pUIOoA
mbV7QgvielcirpaYWdmkbMUs/0WPlmq08bOUb6pL73XZUHaVAzADo6ijxA7aRvR3+nefc0WR9Xa9
OKO9FQAXaESYWlXxLdF6pkLqXt0xfe/OW8ZnuZc6ieTX9/pQhD481eqKE4GVuVqG1BZhxbqOpkPB
E4CzVPsu+/BPucHE+2ntY+ER5w/x3p9Ic/yLbHN7r7nkx31h8q0d8PzLQihjYg7qENYof13aYs+G
wKc1xax70ADWbkkOdQIvivTAiXVWJJOJZH/zK5S3ajgaCsMuBfYn4guqL+h+tsG1/WdG5Y/PeTsX
JujcjVgGR+Wk1ZbaUCF5eXibfZ654OcDuh2WKFvnCVJ4o8Qyo4ZliXX4vzvsfnxFF7ePRzsABgAX
RqBE9FumpQDQIYwg2EcRCEphEykmsc0wcfVCTr+EY8k+niqCRSmerlfsfC+417gB0/3VqOQo8Gsp
FZR/6Te+FXWsrBTDqdHWgxXbN/zysSnvPdEitKtkfcSyijTpQ1EsGB5VW46vm6CGMJE6jpefxwEb
CZh/AWcy1BXeuePjwHXWVWx2YIUJkNaowuH8b61NjVaPYccf1DPY2z7U3tSKuLq6anuZBrl4xv2H
S1FXVbleKHeSklgYzNJu0IxvFEXPKFyXK4BYy4UD4JC/A66kFeCvVkQ8AtBQli1JABmrBJppBWbd
A0g+GOWeu18WdGUKK70dOoQ/+7wkK9RalL753C9NIeaYT5VAm+Up3fJQnyNhQQa1cNEt77VRn0/n
fqCot8SjXKFN8KKlG9ngx/Q+4OU+TT2enLuh0trV3tD3H0vt3ux/1RPSvB84xA0OVgBXr9LFfQwI
hA+1AI3Tgs7zYfl+vMwnnQnYwoLUSq0mUcn5Alp+L3nDi3TQdCcz2p5eYlKzI5bmoZKk5MThJjEZ
pXEtUz7hWvXhR0n1EGQNQGkkwZMFsjT8bvvIBi9Rjqg/ANx9zuL1ST6oPcPoh+OUaWmP08Kr1mlg
6sW7lPCgrH3AJfqbGaod66z2yN14FzS2QFc+Kv1tT8A/HuRQanHMAHR0zC7aiBl+oyOh6yKc844k
y2ezalOwOpw7fLdRDl3lcs13DYKVq1TTuHr26I8c/Z/M1DWW15Cqw72RCbhekc54dPC+jt9RPwQO
44F5s/p/4aPlZYuoLgw0yg1gjplQ6dnvrOtoAz1ZSoEziBVxQbZK4hfKd5LxIliINbZLCze+U2iR
LBGPaSrKWYxnH1xwemNZAu/Edxm0M+oTzy38dVQhgdIy4gdtzCkpyVyCN63EzYVD4iJp1AmFiYly
s9PPa4y0HHXXtCqtThFOh1ktjAqmEg0agbjsQYsZAasxAhrKexuKEu9krcNt9oKL40Ne5I5wsbrR
HiNt+Zz3U2e0trliP28bDBviC658hR5ptF4lr/7YPkdNTE4McA4r1uFDYYoYY4k1WpIRUJ3J9uvJ
8be4xKXptpuB2mKaoXV6wPzm8pWN1fOUVf1rqQKEN6qeTGs2VXaDM+U38p4kcVQM0qbWzYq0qHSE
100w3QVEApia4eNXP2PogjhyJ41tgklbHhk0qwiS49MjOu0jseVh3tG31l5jxdsdrM/pSRDsxTIR
Nia8/WDr9MkdHbtRvvxMHNCIRfpb7+s3wA8U7c3JtgsXcyxFnMXqNNpeOQRl6UjJKIy0HPEKtwtO
1bKNX61FrR+r2VQzlqIZb0IHdPWRNk0Kmur4FkiHWsQU92xoPSApofVfVS4RAxNmzb4qBJemcbFc
kFW1ZTcfz2ltlQbQo9soRzSQegbkIf7TBZ4UqJzozA5jLh5PRYMD8bfBxd/13LTr+gi5N9MdLjd/
vvz+fQQDe7bfZJUo1xoWl8dWZcBCSKJrsG7GCbJbX/e0LT2SlBImdn7fTCWCWRLdeYlS51ye1JEL
4u0nLJVh5Y9XVtBVgEIxRF+p5vpxAlX6EpAvZ+m3UyN3L3ZmMNmbQoNU+wjn0+DOMe5yro1LZ2sm
sSdLysj5qZrXNxU84ixxmv7cIGARgzdg0Fa6wI3PKWAUq8eo9lf6rtpkd0oGdGxzpH8g2D9PQEsd
CfL+CZkEBcCw8djACqIoZ7+tEdRCfFyL5ujOmdS5vPXGdQTDIBJD3TOetq2WUJTxpLPlarzRjBD7
rG1Am/PeiD+i+y9/WevE6z7CtTtkrK5mzLUpd3PgKsSppTWBnxKJpr9Z3GcV5+eWIBaCToDJa6HB
DGqdQo+JMwjOji4D+iJzKs8CJm8OA/VjJ/Z1HjB1Dirk9bT0yDg8LQStSYlRc2UvdwL9m1JH5IUi
C5un2Rjj/+K9PD1CZaDOVw6AeztcRsvqeW/rUUCA1ottnZ827SU8Y7H4gypxVlUb6Vwd9fyIINE9
R/RBLvPrJ+TtF88MUdlZZKbJE2wipzX3sau6wdzkxpQ5QgYVMGhTecLuZnQRo5hAnqDTFvWhkGN2
Q5HqAKntau9sHnevyP4g2JIn062JqsXM4w6RU+L/2uR4Qs8ldjS9vdtVqEtLR3fnoukUEts6e4es
LzL+IXpD8suyzdPm7z0rP2ABJHTyNZukBKztMXEF5vG5d16eTyiEixv54Pv6pLyFtJbwIHWzoM41
fdEttarNPaXETsU4bFtt9QzzCDnlQmU5N8tSvmOE5o4HdKihn1K3DwuoHZnH1RF5tY6IlE249Q4W
6lpUzOKx4SWxThOF41c3nC9o7Rf7EqZ924F0v4Xm3WOc4fwRCyV1JhM+k1C9ifSO/nb0ELaPeNNj
fzm6fsQf4OWIzCWj2e5IAgEWrxp6aGtGVxhzOwUslgaYwE9bj9iyJFAaSvFgCvLWatmERne5tL5d
BhRzgpz4ZJbydw5Nn5OHzR1yfH0NOd9s4WrUj5dr0MwXSUlNeZdN1Qbtmd/B8lEYxr1qOKRUlybN
R+ilIMpZakoy62i57qahPN4VGfyt5KrBfdUMc7dRpeqT4x8bPNFYQN2WYgDXvj4c+q8q5Tp7Xpmz
FpBuDBd+ljCaDn1/MrVmumU9IjHkbJBRJvjyExyXV2d7ncOGbSfRX93mw5gd1em4w/Lw3ZzOaFVM
qlafEVOvx7+t72whef0BTkYxWGWEZBCtPmXgOnOglcQ+ZoS46SuT9hfxJGBoZi1IARk90t4+rsfC
FsmjQWLimZrhtxFyghsPLi2fJ+2fNa8LvAZ/Yl2qYwu3myYXu1UNknmKn0JM5w9T6r5tqf+xW6ss
cDPI9QcQLLD4YxvrjmVvNyRiuK3cadSl+etsAk1mhESH7L11aTYcyD+pIHVh8vK/No5liFRmuA4G
78Z9EOm97GKawMokGExjQJRCg1DhDzbhq0lSLPEzvcfNTa8XlbB7gj35rOFxXoMs9JNqAlKMl/JA
Y2GjCe1uzXjjFYKR5KaekrJDA+i+A0tqRId41qUAmSYM50loDTGd+ADZ+OdsMxOwSWOvde9A+dWu
nkM3sVQ8PJ2JKBNRZbdbKeVjIK6Z4i3BdGPCgwKwSoCRdhiCJE4n0oPg6rei1XAhk86pO8OL0s33
8KRIzSx2xq9c3ikqLZEuGTs2wf7tXRSHuhFuRr5v+mTz4aSeCRzuGH8M4cmaCVwlwyI6IfkeJ9Lm
ew5JX/mUP2oZtQszxxV9f0JeI2VakBGY2LrzSKYQlPtsgmf88bLIi1VighmGl136FD+u61+LCOjY
/3N91vchLf9+m05F489Nl3gBZNgWSDKgjgO7UJ2K6DNnn9wwlxKYDspZx9BSWayiOrCLSKVu3n57
CX/TIpgyQo6mTG1J4slG1i0lZP50EfBEiMZQznGEaSEEAkyXzuf8z7S6KmVDAvE95W3+lFYrA9no
9apaPn7dvCLeGcMHaNXQnAs2bdV32n88xoW+alia7DfjFQGHuPzVS7ua8DT03HLuFNRW4xErBPqv
Ye//sULrl77LWlpZSqaYD8WgzhsK6jMsI5CnS9UZP6ZfVNmM+uIQYQ/d3tmdokOmZTWAme25rybH
GDiu9LVavyo8tABaP2/AZkX/3PmjG3kQr3bHtQpPwUJxW4mtb8LHVBQGggY7cETCY84NCtDrxNzP
Y0NpoaxYGWZeuopMzcqSU+wb+9UOjXF8gLPpKNTOzZEe7WDzmVNnzOo79nEsvJgxhKsD4EKDT4U+
llaHKV8XxdIn0467Uj7JgJ3foLPWa+5PQqgSM98kyoJwg1OKacHNaMYyHnZj8n1lwLEgql3a/FG0
4TD8XKZWzEvLoemRdnfvp0TNcHA0vR6dq4qh4LRlHs4A7ZZ5kuK9MCM6hpTflAZC8oRuqLj6iU0b
tI20aeVxAleGYwt9Vc5OmjzOWHt3JTRE8lzyrjRb4nZ/6gfnT19ZD/cOFH7dRFk6V+Jr6hLyARXZ
JOBsN/AK5r0IdOp0FV6B0ke8gcqzaU87W70ml0/eR9n7rjWZBwuCv/p1Ivlg7gsJyXE2Iod5CQLL
9D+rHXMkCAgMYw4CpWDe9tlFb8PFbxsofjiqWOwoxXIH5DZM+W5JGxtid7ZBSjcNMXJqilJSzEcd
CeZrGWZqIn1r2aT81zxydH68+0Pm+x9sVfDd4DGK2gFkG4xVq21Tm9haGQ3rrVs2A+5v1M42Ac++
h8TutEWJawGhgsNG2upxwRrMCVDqvTnXYg7K00vIAXioucc6yBemZA02LAsjOiykTKd/L+xfOvsF
Us0yKM3Qsn2xhuXG6OtqvpoIJoiw9JWYwVKliNhhoHLcz56MRMLx+2LG/P5pFvStiSetvqRjkgjX
xgZFY61x061zPzMduvaSZfODIgSj1qocBr1I16DvRbXV7LpJ+pJf4oqm89TG8n24r04bSlitaa1O
FdKl85tfAtbY1QomAAC4pbLap8DNLY43/lbOK8igixqrE2yTe763dgpWAX22+zOsVDAL4P4ssrnI
ctZ0X5TFTnU7zdwqKu6on1xt2LzvI0SGmjQC1CIOjkLS045bhFeOxXmmWMjLptpZ0hjXOP6j3BVo
JJpCNambGfoIF/GTb8zA+aokG0rwB+wnqYrkW0eqWmn65GHS7mPAVVvXK65GELGzaPhgGJ+db60E
iwuXRD0SG+DM2C17nV93Qyv7ajNQ+D7AOqHwHkWMrz/Uj0zQLjesKIF3wae8cdZJC2MSQsPDbtdz
EGyqCPlMqwJb7wyPz49Yc8q8cMx5XZYkAYYcJRGmEDU9wZ5jP2tVxxC1TyobhsiU6j+8COhewcHH
SqOq8g28aPx+7CAM7Tvw+8xxP2ClX1fY8ZPFRQydqWB+MuKdRF/k6jpyRfTiZ+84nzrO8CD4PVgh
ihbtgP9n0vGVyITvzh3DsbO4Y79m3GGQ9PxkNYwPoRZGVkCxYxw4VwGClphxcwhT/e8ImcjmjHYn
Cqi5X2E3q7K9B1cfomv+6XXpfs8rOiDaCzw+a9Qa57iK2rZyA8a4a91sBka5IOLQTD9x9eZKtqAd
poFAU7rG7zFgTzTwBRC4praq70iOSpNQ76W7z5XHA/u/V0y8x6nAPRzRYh2qiQ18ruY0gUF1ZtYX
CpxpNI/w1O1b1m2SxfLIfLsyV07jlOO5c98SZsM36T8mt8GRgI5nHUjGgEdww/5/op/RfLf7+yAA
yvLKxNjKYMuHSrskNJjSfetOFDPl232mwhbPzoODNHxeNmWB1/thyP9YtxR7ydBM21hZKrTdb7HU
sKqUOwx3CGrR9BYcZCqO+WED3AtjYk3j0vkq1RTywVEDhd9vtr+b6VaSxFthOemaTkvfYcf4Wkmf
nVnF0FZL1X3gc8k5I32Kh6YRVm5to9s3AOiOolYJrNW7B06vQh5OdshB4wnxl+G505pimPtjgsgc
H3If9Cvy24qLqjn8ZxeY3gi6+kBgos1bxqdWNugjeOZEO5LQ/7W/43oMTspeGHd7CesqC2V+Sc7J
iHXkHBWS2QgBjeRh6jogSAm3FSrOFqMkN8lT5SAfmAhBNBHhfU4UQu25b5sib2kIQFtizAue9zUO
Vmh2gKJbyfRK5nGk2CVny5lYoqnsDgOvfIeixM0PTZgLPkVwvPeeE7aT/FnF8N8UBk1UjPcbIRfA
LtLOYZR/eNo20nke50NlxlJRkQwkx/a8uqpmAU34Ci3PevSO2y9w8EOTfVIdVxD11HE3Cy5VFy9Y
KoxbtuHk0U3+CjBPcpR1ecLard2eOjZF3PWgGT3nRhY0cZOv6DNZ2F0wbL3XiuM4L6ox4cV/cLFk
A6R7pkZzPDolX7YTtq/46x5l2x7chXmwOMPntvCvooyI1t6MSl7A3DfSe8E69jn/UaB7Yzx0UfgU
RRrdyvrrGAlZ/iiSR2+J1W+BYb1v48Wb0NcN4m00N9pApPob6t2JD+pGlgqUYLyE02tl+ewqinm9
REFhsH5oqssoGOepP7GS42zgzEi68H9emulHopZHHyBvptqwllgFOZhlBSxyCUblcXqB3n8AKqz5
/ATprTgUqqeAWM8CJ/RkLEw1OOnJtNa/RvFMKabJ4M+ucdz+CTws4Qpwr63P0iYR522g9knAmMHA
rKbzMZLAttDF6o9NeHPq46GHZtzayYmCoiOk15HNQmZzwL7B2PsmUXBZdtwGV8awHuyt6bGv4OWq
JYFCQWfVkev3RfvNPTfkQv5Trs40c7Pfmfo0B0jIHJXr3tML9RTAGAEHtYALk2CYieYlT3uyFZbD
QciFz6ypIbEtbQJXKmj1BP+SmtvgfTLNarqXZJncn668X4nTj16Jcnjvm3cW9r7KL7bS9NL99EYc
FsnLn7c7PxzOPZIdixpWaz3I2/zg6xmc3CziFEk1Ejvln9Ct1A6XUS1dSotoYEpbFVV0gkvJGFtW
kSa3EDD/2Eb/tXnv2CCV7o0NpaIiXQ8mICQsh7eILmCVuQw0lMCpcGXx4dX2YOltBS3u0IpEc/Wo
uUAtSp9UOIKCbQk3sshjN7YE++tQFl+ntNofeu/8EEswSO00NDvSmNTkai3Vp2+Y2NGTBNtmkfqM
tIttXJd+F8x55k6WPUMY3YVzoqn7jD3IPxesSkv0gY9wRcx1ldrQBSRibJl+FGPrQtid02vkgSUT
fm1aHdARjmEFcW0Q7CNTxnUqn4PGwxsXqu8j+vUgVDSHPN8Fy/CNMlYHjpvRhvYkOcRZR0pQr/PY
/0THvXn8RT+VQvX2jkHzesJp/AvuC+wR9wS9P/NK/H1U5EVhWWGx5jdb0Sh180ceLy/ZS5DCJWqO
CyIL7P/oI4bHRtZNEmGwQLqJk90XAW/Lj4S8iCg8cJNizOpWRbSx90Cbvinnef2R/2/3oC9ii9pK
u9iSozvDODkLyPQBBtOUa1cerOY56jqKCB/95Zk2+IboxxVgv8AWxmsT+IRy03cOyrMSDMTzI3TF
xznsYq4Sbx6TgLVgJcizenkrlEVl25GQWeYfYFii1xElWXP47Llu4JAWj8L4xqjHKv6iCKVhFrpM
XKPDYkcfBsHCwlYZbfr95o/JfRAtC0Nd4vLJiCMbPvqqXlQRT2RRfLoJkBh76d9qOmJHqz4p2T+D
KcDRAS/8SlpIERXyBwrsFPUyxjPkwIMmpT2qrVg0DsV0v1aNCd10OnTW8Neq2TaiG/bsKuIUs98p
Fryc9SrPM43lK2o6t3U2iz6NT9co0FDcJz/DclJP/8hX+LoGOgS4BVg0S12dMO7E/dLJ7F5CPHrn
cd4CljwSHuAzdvcbAo0A0l0dTyF3Bc2lCcgqzPFHzq30A0DnllSiBSHH46mghszn1R26yzLM4nMv
fhz+PtC5sYNSe2cZfYj0jMxLdIsgl2pMTrQ6zN7yxRLsnYIGDGR3zjvvpQkp41K+yD08qJp5ZtwO
/Mc5JNdn4SjHf7JgLjRkr0HOxjbGfqrqpl09x8+w2rf17dnygaa6DRgxlhJlkYd0Te49auhGp/bz
++EmzlCCzUqUcIN64DWYzmH6bxGAQahktDnvyyIYHE+QDfbyhhAr4l60ln4lmq4JImPUSygmd7MP
+WcFCFjwzwxonAZLSgfmJSBQj+//bjCH+MCEc5ivtFQTo7nPepaDfvj+hzmPOZB/Ia8pK+T0wX4M
vif0VYSTh1vW7RxCpdzkqhAWrPvnxTJxa8g0DICLgGbrCAWMPmoaPqPAmB6+2SUhYML9Cmv9o3+4
S76pEVLo6YfZKlXcnOwkbJFwt0mkWVAGvCRGjDjFyTWj5BxEeqSJPmohE9HWlTDNn4kabhHw+2QX
lSUk1TgCl48cD6pimizNu7vIbcfD84ruf50u8ZiXNcdaEl1cPSgKTRZkbx/7301RgM/k6d7kHFvr
zcAZc+bS8uKC3LEkIiX+k5jGgrRbpcGfH8ym3JvtzCMqHOTPg39zaA3HiYAB4ADPDOPcHLxAUJgH
ZwPocKABM+VhXZkkr9lrZrvGOr0cZgW/TjJABNafg9NjZ0W8LoM+tSCXrYkpZB+vzF04Lb1NnPOI
RZcJ4shOYS8XPMh4R6GK5/hrM0YGLmPFcoNIggJmpKOfG4t6xzPuKmPg5L07hTOOTxjQmQ2t8zWH
ti0v6eTb4+f7ndYzqt3tfjKz1f5qRY/SkBTWniBhXzQJtGIwaWmgxvPQxjFSNyscRR/sq1/YAWy8
5pRdWeCSDeaUvSSmlqmspM1gdmpHdvaXM+/emWOc2bDKUmDU2GN47rwKn5Gad8QLfDqc2LRvAxcV
sRsF6z3+GBNwMbxrOoUj9o3wbvD5hJu62+M7IVVuQFOEzXtvoWoBgdSmea0juGkdPKWcrdPqnzPZ
+w6fqYIVQ5pMrng6ShTu9P0vaxRGeUVN9froBaHGOYahQus8DGc0SgVpm6tYd6EP6fp/YMKcMNl3
wW+OMUybEWrQepNYgvpo5kvtRw2qn8ngLoAXkslUglRFHpwraiG5hontjyaEi+h6JAc9v6M1gti3
eIFMe47I0Cjg24buKK8zAYdSEashS5or6cUMwqW6TQHWtMnhAOoXAjHgLFGT1K1G7Eo6bm4j3Bd6
mivNvg7CNsQvrOmXyqHKRu82dFM8R4wTGNYhM73KS593TQYt+OY3AyZsDj4+LqaZptHjwrpAJtRJ
FMWDQjbVgg29HMiX8OfA/EOUkOiqPHTgjSder9tdD+kC3AiiYHIxeJ+V6ZqiGCmwyLjvwcit6iPN
uL7NrsGfMdxAqvnkagNR9OBCW1jokgDRfACxN0qJ3I5bnxD4J/ifNv9Q2DRqmsznlXAqV079nVJd
G8klghjFMGgz4q9HcEt8UMMpldCcPt5Edt4tCaGi6C4qbSyRFkC/+KfYb/teV3g0ScBaNoIMcUv+
R4kJy+k8TaMO7xfHSVYJEnyoMB0Ddf6MAbj7/ymZi6vElmLMdQDFYNyJ3GNwiKeLkdoWL2iNW2nf
cxkno8tJv7Glt23AfGMWmgHkrFIREDHgvUIbJ5vYoxbQY5vxGyZVEMlioPa0lYVUkI0nfFACgkrD
XyOPHyOTX3ClnNyyhwFE640scJO9HIlzWJtIaNGm500LwSUavwBGSa8ebI8nUYKr/jGt7QPPhElr
BqEfWcMkFKyxMrbqWkcqIGkSv2UICXuR4l+jr0b+AHGVZd+Z9m/uwF7AFmABzmey5pyMTgdubbex
IPgSTWRlSco2mJ57JOhSxg2rswgeX7eetg9kJdZ1pfBCBOgcFxNHCrFo9EUmE2UwBHedHRBJF8V6
iQZJOz8171e7MtR3cuPDNy2cARqtv7sgltez52I2p3JtDFADn6TYrzJXWq41winy9w3m838Aanwk
3C0CQvOP7rqoxhdSEJ1BCNiDfAbuRlS7q0NnPG/CTCPJcdcYn7PAlne+zdXuyD1yic4AQDkShbpz
9eCH6IsYAvKag8+ST9Ty3ueLSCoURLJT0J61cY1tKvLZP1GLcM1oU3e4fgopmxjZWNZujYsEpZ4x
/nYk+Z/rgeoxwShIWIlo2J3+vCOD2L8VYVvh378dKT7nb/eV1jOyQmmcR7WKl5U6lleB3S5GnL/F
ch4WTwrlo0I8lW7Fj2HZsLjOyMnu/4snX2/pYd1ugLfplsEzl4fo1O9ao7Pvpo7bpJ6XyxiQy5jB
JqiAjokUnak9Cn1s4nEkPRTM+nWf0r66vdO7FmgVZO6CLAFPWma43a2MSFWON2bIq30O0TV2MTIT
Wihrrb2cbZqOS8z9bO1OxkhiG2VIMYmiyoDx+OUafzAuTkS/1PeWXORi9IEKW0CyC9o/FOh/33Ss
N2pTpsEvszSLzBQXEPdu1VP9LnuyGkP3yHhuKKCx1ZYWXG2HgObabihyYROEUUw9hp/0OGi595xR
HpwCJp1WkrBH8s7ByoFDzgo6AOdsjFbbI9q7+CY/Rb/7fBq2MAmpENXNQUduRxrzrV9yU2Ga76r4
SqrjVreFc7v+Rc921L0KXTTFYDOhLXgD/0HemvVMuU/OosFbKBgmMN3zy3N6S6eoAa/JAmLCOaQ9
g788hk7WcQQvzDY5ystDBpuiICW2/qXvCYqlYGXUu0r0AjNA6epWn9MJxYUnk+01xzpkFIm1gDAq
wj4hqqn4LONMKZJkeEyQf8rOoYYC6eEJzBiayZjXnehBzCpeRRSXnmNP3w7RmumQ+E43oH1uzCTM
PbCz/+FgTMpJLzU0Sng8oj5KjLdMIn+f9MaVUmDnswaJlKkcq+Ql3j77SUtM9Iv9nDe9aCAZj3sc
WCYyS+YjOmw5SkR9uSGOGP2ZFhhK6UL35Skr++/hT0c+FjjPZDPBfXU6GudU9InPiDwt7SwY/XE4
RbfXFVse+gGM8LyUfydKWVr/F4FsewfMhT5PwCgsFGz+inlfnr4rItvmZuuf75uAMZ4/bNo5T7dY
fX98Pl2ytRVtt4HeeakjBfTcYLe7O/NNLA2I/WnLB1qQ9USrpRZTYKvajVYoTKgmfpe73xiH72Xx
PjPf/OdC3qOPEAce7aTB/UIhYNeLvHDc20tP+m10hgUBTzem/R7qTJTypXG1khGLSV2kDZS1wUd5
4wDaKdBk0wLuzsyGifJeB8aWKhOlmv0FCTUQsnVEc2JYtLxqQdVxg9Mpe14PCXP7sQZ4TVDxaUm9
HMhHFjiFNfnC+bznvoPxdL01Tj6HCrhTvcvz9xJCWmMhy9CMt1LI91+W30U9tHJTvJUkOeSDdv23
1mGFk507vqg6bo9sk3Zv757zDky24VQmkei4NE5BWqYGvQ8GvP+O467/qn8xywxwTpjA6vsRVAph
qbG0x2n5RtLdEvPxfbc3nlrIIRG8ERA8jBJfD3Tf/ODwTeH/mW1WS95yUh+SulzSQagMlH+3KUK/
CALfH7ygloYTEeErkGEx4Wtm6GDz9LrFJS9n+Q0KGmXYG2viM5CL6pSUAs4Uxd5SnruGlBpBfCc7
gEVQWWB4XSslPHeKT35tJpdyn1kRo13RKjfuM7N6gyEcZ3tNaZle+fm79WFW+hvzaHdhWPyoN1Lf
cJI2631LEuX2H7n6So8r4Ym6SSMr9VThy5oHAkI70iNU9l3QQswgzXcatsGhKLWiWCf/j5qh6FLn
BjsqfoOZ9SvlvA1/mjrDorX/Z2bMFYbtnqZ7KbG7j64J682lJFRJDAvPBfLx8A4p0z6kD334h07R
ETiOAOA3sdeZTfS+w0WziY64HAMmzKEiSdOrY2wsRkBrI2LyghnamjQecTe6RLtItQFyn7JjpHpe
jkIcorZu32Q4P2ptybl7mL2lXhOpcstUuN+PN6BYu/t4lBOxszqCXadDhZUUO+R4khX2YFPpO9lj
r+dheImm6Yvom6tXyvCVLBfneetnYy8faKzHdA2+GzBk6KfZ383R5ZfiNlMdCmQDgZvBDu+uzM+s
XK/7O+4scVcC5+rwMXtMV+0kgc1s2LTlk39R9Uh2XYhipacNfytSanEsYShwzSAprp6aWBqyjsBl
65EbdaJvpRsw0hUSN1W5I8n6QKOcmZSCzbSXS1rGz01WXWO4pbIRheFNz5mIh2UtGYZTONBBdDH3
hXoZaU+s+C1sFtNb/aCZpEHxEeH7YMWmAIboR8bIh3oW7D0vGi/C2lbJ0fLQ+q4k2l9eiFhJQ83p
0zkpagrTaU/RLL/CjSfKLG9JOHuDtJX6tCJUN0xawPUMSHTwjYYGIzrsjwzDgK+g6fj18ySUVrBd
Ih2n/h+MCyByCOKQIlEjEAL33SwmBfqbvrOVzU0NMKlX8YQcGJfz+UQbGIAc6jrw19qsREtFr75l
zxs9EkD+LlmjnxE9UdZanPRP+nR4kdFmxDG6Q6kv1JiBFOxvujOuBclytB6D6svbaW3YBoVkBTNN
lCfvHoYrzbAu0zSmVzUL8dW4x4ZOAQPVApNoIYnYiUxqPeC6GtU3TsP/w1+3dLfTbITmJNEI9Do5
skdeMewwybphFT8zqHkrrddlWhuVcQwFWqoE26b3CMoAAiJlA/sOTEVJ5DKFrLc6Zd9RN1ODP7Lx
CM2w1TkgbDmtXqR3GwdWlJzxaA4n9f3zOd3n3N9vxYTtcI7j2EhtYzsn3Lz9sbApPJN1Y2QDFB8w
Lrg766TgJjtNEdZFA2PpAy6RC1U/JXGOLd/SEfJSPHPCMwy5tByYsySQkAJGK0fRFv/9OTSaLMXz
EpyYtG8fI+BjMIspaYlmZOMG/s3eZdNfEdzZhEe0cfqeKQuQEGonFZp4ciYxPdnt3LKyr7gm7zDo
oVcoppBp6v6SQUJqDYx/DLL//PSW1nwM7ZK97htq2ISBO7UhO5dgfsihP7lTYU+OrEO6o7/O6pYC
2T/g5s6Vykl3EbnBY7KzLblPh8aAfRE3EXzy0rB/i64eU1eiUsrz3DhTQGqWju3fWcBStC/D1uyu
ZEjgJhxoX9iS/SjeWyaNr04HbagSV5O8IjSBbUsZAq3YB64sgkraANxXf//0cxyaqLkcBRht2tjz
lNrYuaBW/+tbyQohBUxesoZyY0/Rxuu+ekqADcnxxAKc1WBiRWBz7QcZouIPdfBtt8S/cj7LtpoT
oflHU4r9BThkeEExKwrPlWJbPD2GTWiDW/NoUf6kFo3hOH92kA2nMnpsvMBcfP/XFqQlrieXqhdw
jEhOuRcBs2NAcr9SQs7FDLU9h0q/CjrkNfqeB4czEMfYLwG4Uh6eiX1ZiVu1w1qUmNJkO5rp8sVU
EaTg7btax4dtCrkR0S2tEPOudV1VMIo0qBjpO6fPGWZCBOhf6STRdDPizaVnFYTl+ZB1glMNRkmC
TayrjmGUqLJTeeZ0mW8v9vFGTPtMzMgJ8GZuOigQIjc79OSrnoGOR8Y7KIzU+DUKUPkECAlIT+7Y
l3HMthR2OqpCuds0qeNJktswLxUHYVAweP+nShQ2jIhnXu0Z8YCar2RY2qvnwRRRHh/NP0bkgRqw
kUqcQn0h4OETV7iHwvDiKfsWQ3qnQwAyBMRfD2ixUWNJoYE8bwJ9jaLoD6nzSVUcmH8suwbSjoij
mNzZ+Ced27V9BVlhBZnekNFKYNx7G3gRgFnV3UQYxC5HhdBQm1Tb4b3aBP2hHKrk49NTEemIQsEj
5W+ZXtTmQxf5DxMwl6BC2SCWZTEJrS0FMHm+WNt5/Nqsy9ZQKvhcQ53oaaKH1+3AeEZ/OgQIYrHh
3GBXzE8cZ8vo2ySm0KLjVIW3vESBq21tExKkf7L4e8d1g8Lg+a74R3tbc9Bevo3Wr7FQmC4TViz7
5wZ8US7xwokE43vlVPuUvLE/smlwDIANshxQn6MRjJ8WEnU60h7Ejk57xEfVIMvFimmGWPkrl+p8
ajeBfVKk6O43Hq4FX9oaXU92rSD5ff5AOVPZfCkFdQQwBMNIIXiJ3BcYRhUDp8RKAYI0VMW0zvNw
vimEBz5EtEkBWEO9EhNn3ZgHSZVk1VQubLZgfsdMuOzVdCd7ejBTTzGHftlMwC6QTC4Etc7VFaq8
bi7VIePRn3qWeh11YWB5bu1CvxVAWsP5kjTgOcMOD6xF2kLh/rWS+luMJxbbIynjqr4z2V0sdLpA
wjB7p2hO6u0o++18OvUH8d9F3BNrp9/z9yIp7I5V/M+d+iX0LG50Gy68VWF++wheDby/1M0YoL+c
6OS3iDrny4a1NX6tS9Va3os5c9PF0OlX4lrC1zuFJDv69jUj4Y5mmjM+e3OFFoVuaKfqXa5PKmbi
kHbRmCmS9IBr92gc1M8Wad83SFES0NIg5KWAVe8XWmGAXo5j5PUy8i+73rodDdJnQY6DBdfIKyBG
nsblPCDoVVOgBe7OTGlOhK4Lhe3CP2bdcWQqmtT1aZmYypOsPDnBqlx1CILCApwDys1oxe2aWAfk
KN6p+aKIfP4xI5UrDwCz7SBP2oM/NO0RhUx3qlkMjThb/9QRErMy5DkpFtcm8KYXdSse2WHi6MrC
dk0bQD40KhxpMu48BJcwZuN9LwJbz/QQJce5JRZVgMZCsZCkQqgk95u6AnR9dbFrhftNJBmPs88p
xPx4YojDcxsaSkKhFGixusi2S1za7vH0CzM6L3DSy9Z6c9sMVgWWTHSmEMsU84d6AZV6A13FPqiN
kIyKhTJZdR7EfJ++DiCmykTyjEeUUr8rOYInbbZM01Y6MAP97KOt/fBL+9tj4kB6NJMjqJ085oiG
5Sg7pRuocUr3qRIMOsk7tImB3GptDSORsQ0mrURKZ5VbDrD75g7xoWD0HEhy5UKxag1wXqmzl6E5
/9sfyEq7KMJDIYk06tyCkNAsRSaxcWeydlIAYYOL6i6T/Az07YESrnl4Nga8NMyI5CBkVxup5Jsj
RlayIiKchdcwmDt3qo8hKmKFMwSwIvQjOHpk43aadmQLykpsWU/oGn2MXsc1mRyAqZlN3uIVcatT
7qb/Y/AZ5h6HsbNqX6922wZha3g+qMWt4xwDeeXq1OE33nqV7DE3L7Ysj0XHhy8VfTk4sl3E3tck
FhmF832qGxcbuh9Xlef1lYd/1dBvUNNkBWpqoeo/7CPm59d1DVjd8acj0ZR71WMzj0MkXLwf0RsM
kdC2HSwYdAjCxnSRViTKSGnCA4uejnuq1rUpNw5lhciJeKKEHp6lmavMRdDQughzmu3tc3sVzgOj
AV2cZ39I5mqlJoR/0MgHoJK6G0cwOAItTB0fpx57du9ox9UrRSM4hfhhcwznSrUTWzLDQw3tZeNF
0Ntr5G12SESZjlflz1RnBGqfHlXSdYoifzDCHsHn3PM1R9I84waUDeCN0hkw98XGCas843L4rgJi
xoxcpwKEOQ9/HCp3FOSvi4AqfyTPS/F69jw0jFmCUlxzbQDn94mNafRsOF0j9zZXhjazwWk0U4ZW
vP9iwVYzZTthpw/5YWgB8cTp15++Hl+q8VH4TXgt5rKbM+1f+WR+r/b4rsvbMdBfB/TQT8dcQgWR
tUyYNIdYgN2v6oBhKHtgxyvnsYyxLsWeYHjg3tncZcgmfEC4JULrNzQ80i6km3XVTITeZxP1bI6O
dnHwrdSZ8jdIHxfB7M1fVIswS19b++O+NwxkmYDum/hsyNRpRrU1diib1nqGCfNBKhnUEyLgYfFd
e6zbwQ386WyhqLoJKN92rOli+S/92B/S9uEGxpSqj9iiUGs8FIivoh6y5zZcXP0I2QOFNutUvd6m
lskShqDP5LLdlL/XIzFhQGUedtUJAvp51ZgK7XJRZt75A0AzJ8qFjWsGVi6SkZscUbrVXitTaN4Y
Jck+1RghrYlIPSRY1nCmaaXSFM32FxfS+NzRaFEjHGHyzkWCrr4NCuquNRFaXv55awls1SXPFEyC
RG6RV5BtTJI/McE5KnlFVw+lqi0TZwM+t5PlXk7VaaPduO2G5JB5tijVoMIFDVHAFE80cnNd9hNV
FbrYBA8AMSZ0TQ2o4vQI7CWM1ka4j2ZCIwwjUg1MhUrjquurK4dWyzTeR2l05hiFhObUZ1jRviVl
SleS8eL0bzF3ea8GQZbZZPVgFnLV67MTFoW6EdVmBD+/qte1E11ASxtlyDMRLW3kkqYi6V6vanHi
DpQYzn3eXUUzTNMRzv8Oco6YoQv1JEyUV0dHufZ7gnHpD9l1VFW8lJYmDQs34ueirUfOJD0zgpX/
aoEF0ceWwy/g98wdhV3HBiZ/D2qYkk5j0V9CNMgX80jmZ2+KMWK6ilpnEe3jHbJ/JTxFi4FcTMcL
QPar1rBkqpsSkqf8gFlH953EZjtdmocOU7iHVsOhLHV1eXoWJdrUoXJYYe9M3h3f0qL5gm8SohQc
NluJkoeGCZRgKLv5nbUVJSytKOayuQd/FDSTzFolThyl+5sTf7MMuIMqWFqxsGc8EoLOX6pqjx1z
AfzRL/cUHPwEsk18+fQ+yRVNnH6jHa7hjF7or4VVcKga9C4Tf9rbv9YryEaeUg32rpw5YV0kTVWy
dnvFYQMvR11+HI8j/EreEDuRQp9leJzRL/aJtZb2N9TBYqJ1uCXKXtCZi1K+cGCN2/vgMum2gy6f
63Ul5C7hQOYp49ESD04zdWf0A2PFXphYUXiXDLlT1aG1AhuxU6CAGlOlgOgCA1K/Go4EwM4uSP5z
gv7Ti/WOBFT9w/Ujvb8ivmasfSkjgba9ID+es0C3BoRIdP+Y6kX1U8DM0JIoiZ9cgTPyTtyEumY9
T6G4CgwN5TLX00sxAz9rG+zfekr5DcmUKZjyamQv0lWHGSlz0Qvjqajjq65vSv3KNSrSa5LfDCOo
tNBbVmNlsDMHHnfy++nCD0qjgtTy04TCyuFmxR1VVZGJI7t2MtiDJh/ak9EG5q3tjNbliyVrC7iK
HTjbZrGEN1PvVPpZY3mAVBt2Ru1ovWyo6GatQa0tKDOa7H2yW8PA224SfaFytgoJ3J2Q0efQ6DYE
OpCCiIVxIdym6BETBiozv/aDz2PnYpTgQXcrqdBcQwQ2ZWL/GJQ7t3idnwc1XuO0SYWMrumn1e5s
coK6PkZxxj6N+EncUGarDzWDRqLX1A8YDiKcF19E04EAt2sVk406Vc4Q8E1H1U08d38Lhj/HCYyI
ID6p+eeaX2zTsm5pr5sIemIsnqIeN51qJurx/abCoxCkVULtQXfKCLfPV7fN4ptM7o2QRR9Kg3RR
zg49edr8TU3z0AyW89XvzheZGhEN4B6PpUpx+/yThWPj8aJ+lP/GCT7pBMhncmescoiDaooIO7Sx
GFtaYIisIGEI5WFER4X6OV8NAO/C3xli4G2kXK8tFj1CPlEWcSyxQEYUOp4p/olx5XrxCqsAEU6T
ypnjPdxlnyNSy60BS8y4F2IoDwqA1Zw0rlu4eQtDzunrOqCIF2sZAAz/w7TCEio9Wc5UCrgiGtJh
wzGWKBLZJz/Xfrbs1j30jVVvWKJhYYMCfLXmVOil10csH1OUTTk2hUWDgypY4SncbVoihJoY3gOn
x6jOmp0x3j61wzCBGp55rpZeWmPuJ0Ct9ipnJmrTpxkkmJ2vrn9iAlg4adYNA4UqFJLc1u8SMhyG
vZ9g4b0+0iO/0BtU2TshkfaimxQi1CorddljnU7dCmeoi4WL1JAx2WbUNhpwzs0PN0KLDIBaLrOd
1F7MCvIi3Enx/TvDd0YCJMogzskdIi8E6mwFnD4Pcf12QwLiFO8VDS+h+Z21uo/I5sgi/D2g0F2l
3/mplOzkJAmSVEDZ1DhzbXH7ijAnZ8jrWvTCl37/nt/XcTBU+k/YXjJB+ia3DQOeT9C+xzpbf9z5
Y46j/2DHLGiM51VvpL1eRHzCEXb0jMaP3Wd8O8GfgFrPSfKDriD4DTNh0cw0Yk+4Vk8I4Cty1NQh
VB3U8kyOKD+H+GwxmnH10qFk0SyAHpZ9j5ms+zRp4h3ZnQb6TiXuLq7l+4jBlCg64OHlA3a22d8E
1uHtU88E5lu0/NkKL3eOZU+d2p94zDktiKFYPlPIrpsBVnis+Wy1K1aWEE/xqEZOfLDjxDMH4YIi
HRU2hVWc8fYBeFRpWCCbaShuiYodNkpGzqBulbkbbNyTHmoYUpZ3w7C0gN0ZxXQc4o9ZEi3EoJnQ
hV6FOl5QpnAtygvF7P9znvvLvQomna9vRu5+naKLHO2U2e9EBjF/vLGoLita0M/zhgGtitdc2eFd
uQM/GNunKccUlvaxtoFQz/UUEmFUk0bmHuqE+ei2jopjwukC6egh/XrGRz/eFgSLhdsNbq/n+br9
MFN15R+E+oEVG6bHjY8MT0+hwD+jTO8vxBsAvYnhsvc2qxBuMo/gLm5EvXA/sXn97kgdIJojHfCI
080zordVwaiXax/PewDh1EUj6bULLYdtD9718g7oVy9JpXL5cKKnSvE+TUtDMs8MwnCVDrVgx7fq
zaXCjQC5sd1HJ7/YhySeKXTtvs4lD/TAGbM6npakTntJYUTGC4n+4b/vJo84i2d1jtQatO2pZXX+
qkowVOt4/wPhpe8o4ng1njADE+I+BqcnP0HCMlqgEhAPcNZ4GDj1nqxR8Ry9NeDHaRdLNLBE1GH9
OpzOYnujYqEaFM96ILIt6KDN3zeBBP++Mvv/I/stN3FA5OVDRvrSm2L/IQ3RZ0HzglVjuYwGxC4t
yA4E/a7jXM5VtpjJlMMtftpEpeagMZcX4eu5/wVK20J7fBlFWm560D55Qi16eHwm2lwzuIVLcweO
VcNEXiQ5H5nSvQ4AipR19ZeuXXsipMLgI9gOIa4c+1OKNRP0HpWQzCmWJnB6e8OcNq2D9DKZd+ce
OiDcXuJlZ/vGcfeIn+ehFmjSqNHrH1t8qoj6NhKYP0mwaV8sRz76ab/0UfVzZXH624jiMfDbsEHs
NQ0sCkDVSvFokhp4oScBAWrPQ7kIPymdZS4ze88q9+z15yWIh3WiE0w+Uy3Ev8GlcjCPTN156iZY
f1gUpNY+PW/+5ecCqaJ/y0cSeXPsvLuSQCKzfNwbE9TMjerUqeUT7XI06/i3pVeVFynDyKB5n7QV
w9JiNz1tbNtB1eQxxMvgmbOw5l05J8npNLI/GW2TKqT6fwqckxRpH9LFRjHoWp8hJPYmJqqdwXM8
C1OFJdZt5cS5YMVA0xxcn0gVZ06d1lBfM0gq+U8s5U5iJtekOuwLhS/MTTgTEwx3cpEEz8HsIqJ3
ZU7/IpyYFe01L+NvdnaZm00UenkHNbUM2EwtwIPD+8DxqalCo+2fqbPiUH9XKzlrCfl6Kk4ovEea
29aBWEe480GsMqieFsNYJph0OLGPe+B5kiP+UCKXn/O7/izQG1/e69iOm5z4bT1eUvCerrWfvbY9
It5rKyf+S4sLw1sq7ws2VYUMiKa4IW/4/x4H+i0ihG7b8YRqAV60vmkCLRKSfgX64cEM0jKQazI/
+hb9/5cXb5/h/bR8Y2p7XavHFQstPEAgTxOkecQbuL9NBdG/01H8wZ+nUEChjTCIhVvt6jQ2Ub19
4OH1g5hUPrh+JdU3TKilUq6X90sY3ATWDrqyW2VaQpCpcr1L0eCEkh4lKbijZ1FYK1TJPDhAuiyz
lMI6lyCR2ybiiT4aY/jspKu1oYRbH3mEwcpFbXXDeShun6TAqcHIpb9hfU70EyRaQ92R5sScvb9/
D+NMkGNzhB8pfQzQqnGIltbj8G7uumK3EuE/0JlecTUcEf1o2j1b4+p0KOYnd6w2ioYzAEro3Ask
ZB+fOcZr3r6tGBjIw2ZsQ9FXpPlU5LICAMhNo/dihJawPirszJieOn+TRFB0WcI0D0h5UVX3Co0I
FRlNbJibyJnERaEC1UjRw09wLEg5KSpoVSGcZ0A66l4B9Q2pfTy39dTs2QEok9bazg0kG1o/31Vt
OhyZ3D4FPtcYmwlPpKDapcpzwQcuhEJSWvynPCxUs2qbOQ0fRLWVs9Sq/x2dhc1NK59Qe5n9QstP
s337TWfC+w7z8DVPwjMeyX/CmbBpT6qFYxEfNVT+55/SiH+d71G7V/RuLekUCQIAE4pOvNvQozyl
BW8d1ocB6rICcBbtlnsnIfjWP/PaIRnTeTEmwJ95OSEXU3+5rRYcBhjIXNMmZXjCe7xmxKBnfQuV
YIbScGja/9bXuUXlHXiZGGX80h/p3sizuDhFVIwJQ5+YCRysrcxNA94jSFq7iVFAHejfiVFEeHF6
/ZNJR16xssfaY7QJImGZsljGqwNut0PGU4cUUw/xtLVo7Y7fD+x8u9x1Vpe+oD8jfAuZpN9fZFyl
5/AjWD10uhGXqAz4m+g9m2MySH2U42xb8D04m4P3meIEaaOrudqunw/1U4bzpqmEvpoFTBOs9G3P
L4EljuJg09jr/0dndMqYA9LN6BX+kUm0tgqHGIrVQDtCQjPldqpTEvHcEFgZhtgZgXtEygWRJbBj
foR8voN3EZeyZ1Z9BpH6qEgx9jqUj0KOjfDKJXbp18J2o1g4mL3g8h/KW9MFlcqdXLn7HpMfJqKn
TwplRPJVax/ajbi8rf2GHYrt9wcNxKtq0PTpCNmBImC4bg07nSmt6VBPKpAludWnjoBy5RjMcKMh
V9qye6RYEqNPNeJQRXHIuKb7AWTloV/eseE0aK+GPxl+p6vabnHOYiy11RE8rRfVgttLxt/ehuV7
wDihYJZhvdt867pWGOBzfT2xxHwZv57VasCuHnVGhKHv4AKiB3hiNcnfAdwXBj/UCQd1Zu0nbA9Z
xLL7EW/zqUfEwZuu/dbnVIfk+xchxB0MNP9XPjTCt1QfwF3oGqm1S6mUCCv//ehajFNJJvkqTfp7
0rq9ubY8UvQ6iHX9+TqjYs5Ban4JFpwdXDwn91d2Tk9KomH2i43kPq0Or/R+NIa9wOxdqvdFfGJz
x7JyLcXd4/MDbpXDYRsIt+GzDTWG4rLekybKphp5YdW0CI4SuXT2f8se31g+EAJEB/1qPAZCuaoi
egnUGyHzLYk/m7EzTmY42P4Rha9ppDd+qQRHaGsqYBJ63Y26E0RnkL1Bsfp21T2AJ6fQ9GACQLbi
qAd2SBMPfpOUArDbmQTCtx9csCdEKycCYPEsNDrLH+jYxCUUCeeFkZLylmHc9wGlJndx9ETUUipe
fh3UoUWB7qTzouWl1ExsZ5OgYKoeKx0abagCQCw5T8FiR36KMMLWVYtsO3y+VZCe0Np/odLr6BoB
/Oxf3n1Ht1QKYbWXyovY+HIFrmWg668MwsiXLBqXMj1GeeS0tIPAsJ92kPFEaqVWvUwQsLgbE3tU
94Mbxwcr2eYT90JAU4sZFYN6tW/YhAYY4J/eqMfCdhYQNYu1zOxw4oHm3ah6h3uW+9VOxan51+DS
ilAlfUtq8bD8lrwL1GrR6wYjnhMbDj6LKrDRSP/zBEN52sdM5vKpjKPp+27f40hHWN46/pn/mi9U
OvSasRZELwWXH5NssoK6pViRRXj7scQKUWTX252lBu+38FG1pJEI1NuCHyonkpQFAcuTLusMGV7p
DeoAOnEFTgZSS+Mm2te4I1JfbchEMvRB9RDLon97K//LtRfDKmKbKGp3YCsS53PSc1s3bBZPqgbj
48rtjkrzsFsb7aYEJJXj9+ykEdGVod+V4g5iD8D/qrV1oynVYYb96cFdXgKp7jwvuMSjNMvSzezt
TPDMA9M4NLouYoBLj7jTkoKySysCESk/XHqgQYYJE7LC+eldqi07UzEwI91JvR1qDj6jyiOa47yy
QnIo4OVgA8WZTyeSDFf4uY5dGF39AMXIPo5KCvtm1FT0HEKxMNLiw3GY/csLLzaVwBw4F7apnV8V
O9Kp6wQrpNdONg+PwIaIPYo6A+sr9SxRQ/a3cT6MtgmPH+3I9tJrg/sDwIokULxzoinfZl1cEgbC
qqhZAonkrhWHJaZFS/Sw5Ga3Enuz38Dzp2A4TdcKMbQmfB1Y0Ks9ltZK5qUkZpyqTPBRBA8L4mRD
eHEWXTRwUKTD/3I7v+Up69Wl96v3rSSCGK0oAIR4d/AJYZl2EmUgd/LEY+rx50F6GTgaLWVv+rFs
t1rEuxHNoRRaNnC1n1ujF+W3x1/dBAfLOdfPnwxuXr94qwDRraQ2cKY3PO0GwA/G5JFK42KSs23K
D5UeYLzeZlwA7oAko/lLsgfjV8TGQO0DILV4lIvTTNWMpyfOnUlbxjn7bMBKuEi4Nlg8/zShtzWZ
xfOwHsl8/Nzy0EEKOkhHhsia78RU+mMubglYtMsN9rWDTlMdZ0CqfAyzHKp3a5u94yNTQuk+xeat
CopLe95vk9bDHckh9wnpcgNLXe8wJJrt2DGtqnDK06VqlwYSbwTsCeFerrM+W6NuvCHTLBMWAaJs
iOR84cBaL7G+URfXWNbfHTgit/JV/mdmI7pqdd5EXlpAW+CJ/I+dTAlzCDiw3KsTRLXQvhUfd8xQ
jfTRJcWERHu1HdILJXre7IOTdzB3Ww3oJGNN1GgkTVnV9Z2nWqNsyeN4G4Gh777lRfSQ2U9cDVuh
EmVyy3Izo6gKBbmbmoWR9/zmIyxGXvnW5ZL6M56LaN2Fc+nerkbmPgxVHs5hOpXBNbcGPvYWri0P
07ycacUsoMOyUiOs2z41Xx97801YxA8Dy5LA6xscitXj87OZ4PbsrWr1yPldfo1PFJP8Vlmwl/r7
KrQEcAqtLW14ecGynpqA7/P2qmYmsRNdIyS3NL7cpYMmFU4tGGWnFF53wBP3N3KmrxkDAwOFLbwB
2z0YWpgpRkweFOG1qvvZozy8lCw5TC+n7+6EPv5DViH2adehflvmux8fFANiWTaIEQBy7PEFxVId
ZpJfJSVHXMTcKgWw4dI/QiMwNvRgoLpUnISKjXE5ixd1UI7x5wbdr/pOPOhuLuxiXz2KMvlltCm4
q4vhcOU7Bgirt/txBhFBt88dt6whGEfMaJq9bJpBXvfKy0sYSZ/0uDtyHfNhmHarup1j6nTwVzX4
4OTavn3CdBwIPrlaK+QnoQRdXwWvtmkZ4knOK5rQW3gFExWzrAp9jtuX7SbCX25ZplBYSfbFeAkY
bIKW+jczIslZ+q+JUu3iUQQnfdq8F4PE4BI37TMesTYfN99vbURSqo4sRlxGic+b1XlBZFk+BqR1
5tXi43OinLznNwHXVS0Jo8g2i2K9vB6NWhJUVrHgaZu82T/6mxlC6zW7Ul6YVooA8UhlO0jvRjOn
NvKK+Jh/Jq/nKFHb7lXwfnhIdovPx1znf3Dp7lHAX7GWIGLo+ObdZVBHRgqaYdtrxAugj7Wrk3xq
k1hFwy4zym6fiSQhCTLfR4jbneipq9/DT0n2czRxUhY7MiHkVhFoBUXPwsmMkRYRdqyluFpqecW5
VtV19Vt2vRbLlH1Qzny7wHsiaTxrSNL5+2YchfivMeJJ8MwWahd7UYdSYUCvtx/FGVL6f+pamC5b
m41Tz/wwVVagb8dhMKJrOW9ZEwdrUPYUcAT45TSgNS2ibEP9k5Nagv+crZjTBhWOydvknPHgznu1
SO0WlJXEa+Y2ettIUOTcXL161ShePnouI01mRuDU0tAZhakBEvylwfdXqj2NifNPcGiuaL/xk/ej
tqlxX2+Vw1t3okLAA1HEw9G3SYQvkgWdj24JInXKU6RTAMyzVNTxmsedXlT3N+8nFuAro6MQMQvE
28T78z+FycO6tbqnzbOmSnlED7O+wXA7HRcV8Hde2pqdL5NTa/jKjNnkoXedZ0WVyVQvPdryZjht
Ucra3aIN+B0DzhkJe+Rd6w9iXFxT4uFut/kcjfGvnt0nMzBd14MSD7A+DSkOIP/RvdwiHT1680GC
+s4it/U9cdk9VxoXLZUIllLYIWk71C4hD8kpTJPdwH8pm94RHiN8+NuGugMtrmZxW4OWl7zE3CXf
tDRl6zFonKoT21Q8anNdU3Y7B5jQDja46MsJYaItVDZnc/Vi6cUZyOL/WYZR7u9HYeJt923cbTtW
hX78saPCFyqKoaLuFE+hjAC6vYy8CDFxN9Tfvve3gC/dM4cAbHML2Ap+Yo1/Q9NaD6OQ8f+GA0bP
a7RVfAfpkMWa7vbVjY3K/oMYEZU6OXW+gFvj/fDhTNt6O0C8+xV/RRt4Psl4GjQW+PNMuhK5vq3N
NmxmStK6fkBn08++2FyR8TLv/pb1bMZgHkpr6YIeAhc+6I5sB2hKXlDEOMZif7xTDPOfXjVCrFT6
yBbdS574uRgnLCEg9A5hTbYc7c51aA1ONyywHnDWJfS0FV24m2JTEjyItoV/EeN/zbgBKxLjx5pM
rATLvPRK/WNmWA605V05zK2x4gK2xoKPlITF7dUHuQWvD7AbF403Q/Cs6rl5tjQSSVLTHUhiBISm
/HfrMMKvZI5qk1qLHD1uz1S2LMx64HtT3Op9xARXxA91XKLSLWAgSsE/kCx9ue2e2HLvngBW84GC
UFrCs+mlW0t6QDPRflsItNzrRV4GcvYpvLMl1QEp9VKV8BYeSnvDOlzfC7HJWYTI3nBHhSUwZxYW
4WzFg29Wfi0ZrKrm2XFAJf8pofYglDoTNQ5WVnmGujHvNcubA/OKHNzsc0fhvNANgBjD8bRncSYy
0BvgYBDd3sZHprA5QZbNzZacDEvccdieg88s4H58Z0gJyqCFiEZ79es9DpyLaZSP+sRYnBqwWJFs
8z9kyO28mbSfFv0pwZla54teabsA+OUlVZgfTwDdf3jgJXBUZJ+jyneVINWRwm0kGjEmMf1WnOTK
2wtwNKrM49RjU7KbaN95i2LwqmUWY4rwXLElpGFmA6dVSanNUKiSETOpMZLzT/eaQuN3cg73MuWP
iWAMAuwAYdxMN2rZP+ZMrnMLiZss/XEuQ8A8Z6A//N3CmS66iXu64f0q+3A/o3YFVcOsoBhjfg6F
m1Da9qfLoweDCaAmz6T95o4PE/f95nbv89lzjSKM54bg2NlphKkr3x8ZdI+uFl7yJHDCOfdgPVYg
faycBQVdmg4udBmy7kpLuXENBJHmtj0ruSfKUriANBsEv5prbOduJAdky/Tn8T5S9c4c9rOUvEig
e4ThRJMGMLAZXTsDQdiQ/jg12vT437opUtG6s2Pfs9kbyuWbGu/MhdqdQYDGGGYjjLtJBnVXhFi/
wmazPbg8LxRIFlShNy8pJxpJi932uAS1voDsjE+VHrHxvVndbuGsWJKa3n7AQRGPmobJ7K98saS4
WfgQr4wOHF8oXQ1oX1FNnV2ZUB/Z9IvbWYlZQoY2HqXtxJWxtCpF8jPbfLqix4n3MqRlB46gj6lQ
Hdr9
`protect end_protected
