../../../../../VHDL_Files/V3/gmem_cntrl_tag.vhd