`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
IMfOuVszrCgH0ngu1ouJoowV6ohQv4V3V1+Gazj1q7/NtU/bt/5hbSkxOIH8UY6CuIrvK1LP8d5G
dzqe6i5Yqg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Rj3sIfrl5jIc8ouK+xGH9+Vmb8iAA598D71SREywIYt2xeXfaqopcekSzKblJJjcwJfZdPL0dLXy
9kZiO2mtmVgdOmBXAe2YtOT2bcKuxpS6fqwlM2G3v1wW7Q3PIYgy1mQXWjyO2jsud8mSIcZlHuWR
5DtyHA6yt3lm38DHV3k=

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
qpkKci/TPEjLiZ9i9notBn0cPPd5yWYioHamDNIDovefkaHtyEsXG9ctqMlttCIlQwTB1rgpsB3N
uxFWsNGrYh2VAwhBSMzkaSEKPC/4zWWRCf23uU1Dm/QCnGSkybfVmlLVd80F0xn8GQCkhGdubqgl
PRwJQoCgttQUmYoIEE0=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
G/QIk8ccKB0XtXQ6fGfHb+EPAkk6gZMzkFTIZflabNi8KZ9oooI4ZgzE6HKi5upjaTOx0Mr9nkQZ
+d2ytByhIiJagHZ07OuS9gpp/bpbXa+8v4rKXSXdl+9wCflZZHkHW3xrVc1RTLpqjqtfZm75tm/5
/TJx36ynWxQO+h9kctxaZd6wweRE+UOPu/xNRSG+6s6N3yb4PAUCs4uRzDlhCRoWcEMXWYU6KnsT
oa8KPuXh2LGaD/U1MQFRYl2Iw05SWdpwmFWX+XalxTIPOVfTyDSb4m9WYtIgNW31H/oLWD4gOQPn
dy3k8qJ2TkA5fgwhFEmkmycIMmFOaUse+mNywQ==

`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
jZ26NORpmZKspxhxy8E3nuWInS2v8SVmkJW7YbNM5w6seYC6djix60+PuZfxYZ7kYFJ/52hCpUm0
nlkFRVUhh5lOsAXwHOUilGtX6crbX95LdjWJpcaakSXkSao64l///V1aogbquQjrFFMwDZae/Itp
GGStYfEAvZZF8v2cuoV7CDCyqdbNflaLJmv8cNY5vmP6WyNlo+r7+YPm1Z/TCSJwjnIdepeTPWy1
kQm3+Xyp30gQq4l15O2XxlnvMSx9hM2Hnkxw3sufl+8Nif2AMcfY+pyhU1SsIVi/GEXBguzhdTXz
FC6SYAJGYxKQf0WBT8hclumJaE4zNictG3XzUw==

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qcEeIzaptklUrXjzLRqVvKspVtzhkAnZvVXPm+n5SiD2fptgVEbzwyjbN0JRRJVziK3Fx6wqypeb
ueCQWnOKML/tC+M1ajDJ22dLNEunTuCLt0abx9vGEyxsoifzV8Dy79WEc6gj5QBZvCssFHNviiJw
pJ35EblO+QKdVSQblS1KBaiPQSTQkiyaxz+/Qd3UeWb3mlDNdNal5m8ORG6qevEbY1xRDWMR5LRC
7pIj8KyBHZoF9fJvBpVW0kgh26pl4BE+Ys5l71OADSKmQsPX5UNqg2O8G3/obQR4JfiUUmRME1ze
wTI84KKJNC46jimrrZOpzLXBHkFeFpiZnfhkJA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5392)
`protect data_block
Q1YHzuFrv/Sszj+j6NP2B0oxpvgw1c73Lv+qItLLRmmJbEj4BNIW4e+cFNYFsWOXEnnTTU+HGb2d
M9wIEgHkiR7/d18rY4oPgGpGh0dGhfbEvmKWWt2KwJOiPrM761JjwQGyiLHCJIHBDAQAHYqeFv5g
B7avqSCmtvAewDSi1SHfhM71pXPN2eGIoY1g6YifhlsLjMXqKqL9fJvfMILDwOr40OzEChswIr/I
hJDHXEsR5xw6GP7QLRQJTFYtBC9J60quuQT0hmNQ9CeMeA2TD7TfPSchU6MNHrNyHI4AZAuHu8tS
9093cuKsgcZM3/pG3M3mtCOc+Svz73Lp8zSoKAzNylDlyd8YMylrZ54K40h8i3+XUGu7QUHsiRI1
tp/Q/3m9dCh0zm5EEdZJb7gNoyqgvVxYvSh2Q51HUVhU/mo8WpI26rFFq9AySlPHL1P+WJJYHj92
kNY75Hno7/y4V7K4szxQwqJ6vnOn3Dcv1cIveJcRuxCMvrZnT0cC/YV3x/B3RSpq6iB5ujhYMIfd
B8dbEc8MjBjttCQ5PfJ341xi3JGXxe4KW/S/ekB1qX857GEribTj1NqY1lnIZ8bDryTxJno5C7mi
36Y2RTWSbv0B1ZGoCh0pi08NrO/5DXU2aJBdp83gmc90agSZjs3s/D355UOzNZrakG09XfN5Cf42
WgsgB3+aDI16OPOq4yRXLic/6qbUPxvateUwBLlwN4tGg4yWO+dSDYY/Q90f85LiHJ8NEC3J5Z70
p3CWOGgQjP90p7JPrV4KPYYHDknnssdOBzMh957L3yR9VYo7v71sYz35AryuMLImH+MfN3qgti1N
/TcxvVQm3EYbQQZgLvmsB2l03G1vMiajuhTvoBGa6kP7EKYDEK3z08NJ3Sq7ehN0wtSH1ohEK6ZW
MniD1tzZ7S5ukWPLfF5tj3gjtgrPl6EjfRtGfH3Dx0DX36w1/EaHrH6qt3/INV/WeoU/QEKjaeK2
zZPntEMANyffOqonQLBHGu0NZUABED7boibiLdNSioV4msfCodHShhqK1gmOABglf6QfK0Zv6Ja7
aW0Qf0RAaBSRDqbrY3Ybb5nqN0WihE34LyCgAZJqITtbN09EuWPWhyTE3e7L7BMf14uV2F4SP151
m5Eo/w9838NaV/1rdDInPrMmLHvv3cqAXW7jpEOrYcZ0CP1EGJBy1tnCuz+x+z1S0nEWc1Mayndr
vrd5CZ/FDtwHMg6TYM2LkiGN+P7xDJix0FOpa/fecvPPz/2tqYWebuz7cStfwAGrfH4Ei78uBwQA
FVcb1/iV+tWdT//i7B52jVVYYR9rNiOXitgxKGy8koStRBnTeVkaYaiBjZvtWyKnMNrNwSzTPUia
ma0x4gEs04Zp/KQsjOe5svo9L91j9RYZfy2HOlxFYPwCnHLdVuM4j/HBKdp4C5YRSlVPlbUMer7J
E2zomEz+cTjZ5I5SNXz7d3stpvpOWSMqwtiJYh6eIRq8WQjIS9rq3hxoGLksUVDcMuxlb0FkM1Qg
x/zECkR/M8GJ7fqKGAQ00SsWAdI/sqXIa/j8ZZ/aD3+SEYpTpr03DZldSkRjfidrdjHiiZ0SZwcs
WeyDz4t7e4BRk27vdAM9UhZVAfBs6luWzeE1sUT1ej1HBB9k7dnPLxvqFJ6K+pAMCgdCBBNjUSZG
XLRLGMhuX91Ew7lQ6YR7XgU34UkPFYjpg9Lo44KsCwVrcerYuhE2Nq+ShSQXj4K3LSnxAkimb4Zj
OM1AiOuwtp48uA3tBgqKB91XMFGp6H9Z7ix+6sfFgNhBOyK5r6x90qdTHQB3ahfxCkZvK+XUBcVA
saKPn2Vb+r9Wh6HBFeHILBhym0kuuqd9NZ0ZXCTxqlWioINYSZKNTUt6V6HDLHwgcS1PMrzXN2s0
0fRs7MKuz6J4JqzXFhJcYffIxWFWAvprO7BndkTeaJXd+9e03JbQMzi85ZXW2z6OGurpTmG+6S08
8GEtL4KRJPoXdbfm+ayiR/Nb7K68M4z8H8PZtIMcrWsSlNaUCxY2Ppnv1TVPS7LggcZbS3BDwnfs
TKDp5LZm+4uXIaSHCV555Q4WNBGq98IlkJqDQ8CDdcs+pzqp19KcgmtYA2BBfmiBFYiKX39FZ+0c
9awflwQxT4g+aNfH/IegrplQcZgaKz7RNMEio4JmX5rq2SEavBhYQ3YU/MQLxWSJAJI12xNWFsXI
rH47bI9zKtGAzLpESP54hL8oSao4vJIFSftw2nq5yk1YObHnmeqXaIBf2uqvIMruK0xjGYwqs/Rb
LMxSRxI4+WwOdxQ2LMKnzO40VM2akiQQ6fh71iWjNp5h7C8UFf/wI54Gbl3SAB0M6zSTuI72Wtx5
0KClcqItrDwuPeLmFkxBFWKFHR9qYC+2Kw8pYtfOS6bnr7v4aHoMuvROQKrRAO8JCopekw8cSCIS
pi4S6lNO1cFpWNr4oeiXoWKv9BcYaXl76TTfEjv7heKxlmApUpRUu2RC4XqVrU+Ra0AXK2486bB9
Jg4UAxzpJnEyfAj8iMgt6Ge7uhrGFW+xvDPGWEnfVn08QrlJ2fgPwA9sLeD5UzqnOxs3wOW5mVgO
voE76G4L2cNifnwBdVOPBMpCTSVhZuryEUOViN2NknbyKBWDOmPrKw9eeofjBN4FtCWrQuVmO067
TCTdI1Q9rL2wF63mRAU4pWakKLtE2BOkUgjMGr9Lbgr89qjGMZS2/HjVmSK+lVwBhiAPlCcF+/oJ
52IlpDKTv+xS3cOTIAF4yQBwnl2NH3FEENDt4qgp1EgMqZOOgNB0dVLFZDfZofe+yl9RV8Daxo+X
9FdCgwMOtKnDfFqsaYURNbv/bmY2yHi0jh6mohD8brYp7gzdHxLazOyQ6CrM9aY9odq8c/QRTzCE
9kfJMOX0buf4aIDYf+JOeR3Id/kAu0n06l7bUQSywjaHvzT+/3NPeEE6IrFQgptSGNLMGrrfDt7V
l0YS2fxigEiGPr2ARKWh80jvdnxvWDswFAXfUO2ng1WeI7A2f/Nrt1dISxKnrBsgPpyVXqLG3L49
RUq4zQe+qfAvVCKRimLy2poNgMK6ISkQiH4cSSi2149gdYsLmPx8IwTyEw5RVJt4QsOnXOL2iCiJ
Ioc/nbZlJP/Y8P2GtUXFX1W5dWy92awE4dydf5yERzThGnlR7S6ldyYkuEaUubBMDU7O5B3xrldR
XroR9m6lPy/E4KVvUVGvVNhT2DS/H3hhyP25VP5N4hzSjz5jSU+IR9QhuApVADeXwxDQV0v1LIgU
1Jk42vPIEGARXk0OqtfKcDIaRq7zuVBSDBSzTAAGOr64/kwMyEtngGBb03Sl0v7eEqNjvnv42W8D
JOYBTvP56TU1ZVvo4wpTCpx9R3a/fRtV1J07PEdSkltH+PE8VOb4nbBltSQ7HBD9SujiFFS0xmvM
8LLe92xUyXBsXRY6VqAG06OfBI6i7IMd0aZhO4JRK3317W5iQ0Lwy5SNQm6F+DMIIDvE+Kw7xhTG
psXl0dMtWfT8aSqKqiPqryECS33zpISkjxIEi1PuBmBIlHP5GIdWlU3QoOcY82k4X/ym8K8tQO3M
2tgOwXFzZsQ1XHQGmxA4FlnXLejf7v7WImKr1/BxE7UmMc7FbRr9FjAh1fFDqB5nGa1r7QoHuRKT
IbCYMj2xZUDwzM8Sa5ndQciBBAE5yJ0+BH4W+LIglKQ/4TIQiU4B/psSqpbcVY8Hv8iisJXxNKDD
P/bt1QmKNzXV1QzhRk+RRk5f3Kf/g681iVTxMClQmvU9anhkFxxqifb21rUlvv7nHdOBNmV6HpEq
466x7r9EeGFobdQCX0W35BZ8Yf2CdRDr88cOdos9qNgcbCBDkM0bP+QmsyiWpG98HmoZJM5i6kVa
oxYu5S0XZhFEsG5HjPXo7cYxiXv0qPbNsmEW+zRrnzHF/TrM3y6QeZ40txSR0Ci1d1pTlCuOqYTe
yXl/kAt5Gc/qRUXJ/oswpIOr0Lp+8z3FuMK00+zUtKWftNRczVjs7NDdmgLddinMvv3kOQ+j29qP
ex2No+OuV4eVBhymelhufDXu2nytLo8WjiwqHn1QWoOibe6fgPcsjPpgfj/mVK4K0X0+QrEpga/M
XVqzqY5FDzZl6kqyHSAhU/huOQuFG4x5Q9akhehc5LPsDPlD5d/aW7U16PKEhVMyClDnlfQrgsbt
K1UP5uNUmI0idOEWCzMXlEwFX2gsbPNBYdS64kYRYGC6/10PUGCc3ZGhBTrI5049xXZV5pJUcQB4
rLDYbuKg2mDRZ2qNgpkfeo11wAsmj2MDgtT9V/hkQJXs4juIzqBDDyMEFWoc/049dMlngHfdXSR/
jy1Z7/jmGTK3hJ5TR6p8n/Oq3CSF4ZFlDBIeIDEJT+5XxQ11/iXAq3uV35V5PLk4rWMh1pzdtx/6
TyDZDEh9cAUfAQqDeBYqlWBlvEyL+un1MneSMqNlxNeg4lBeWP6Ai9aYuwfwl4Xq+7xtkPHQYy9+
09tbx55gpIZUgYY/cKFvKYoPq3uYCLhNeeY215iIeune+qPMN69TWr8gcMz8EZnaJnNPGgEMEo1r
H+4AEtvHHUCPNWFNhWOISa8KG+vd9yw1jM70Fd1UPe59c0BguzvXVYyao6DOE6/f0N5CMVJ/bnox
LL2PH6/xIEB6PmLiJ9tQOqs+ML/2N51jHyL96jMJEEoqTSHsbU+TUe8Bg5e9djR+9c9KZijKiDcR
9THchzU1JG7PLmYEWlwyD4+hIwhbKQ6Z5/tfUZPs/IZFBhN5s0W6H4zZZS0j2gYc89/fv05srsxf
jXLz6wn7jfXIKupcRHCxtP2VKRIN4m93IjX8KtCAqi86bXlwKU/bVaX57zBYZxGX5FaTsJH6DGuW
iHKUMFOh1F3gl8hoWvIzzIVx3B4AWnAG1HUBefofMbjx1iIO+WA0yBnBf6KSLKw7eRvwPkVBxKrU
Q4+rfAF7iVNimTYHcQPJXnbyPp/hMESuo8d5PNYnpULCe2VrH9o4KK9OJfte9ocCOMP7FJNOFHSd
UfwP5N2fZqmFeQ09ROQ9GzaJmfWQIFpD7mPwfczdStHnsmc12UKlFEtU+l6IMi/dyRMmlapD2+cD
xskUxta0cs64jV2MNVmdqAXUy81OAOfuDGZ7/DwvhWg4xPnHKprQanDl7DrS9Fbg9cO6tRGrxdp/
aXa/euYkyrIDf/pZ9x53gcgKp99fHN/4TRJw0TysYvwQ3WGkhGm5Q14a/kH5N8trnZ5QWVMN/BN4
rLc7XTCerTGtB4l/U6T8OogO9qlEJHgLTsZ5wttRuVWJwWPqpFD5xtVioPVdlP9AGRwrSiNSVC6v
vTuLFDyw9CduWvbhwUU14F++0q4fHM5N8vSpGA7yKrrmj1XCvJ/98VIgR55aa7MW+qNPwlooYgJP
8vjKrH5viulAmp5c6oZ5Bvbdywi+x6c8mjAHeDcf4IQKAzFuJS6YNKPadrpTwYYEfJ4OxqQGBP7N
iZ+MwUWoB+tNhGY/EJqTrMt2I5KvM7EPARaVgsAkFYTupH+MUfuSTBfVJIq5dVheUWOG+FCEwoP1
uuVcLlZrbuRmIDmS7EKZChkbBEHw1LZw4S5BxOu1QIMC0TXr0wMMnLIvMkthulW64e6OHAs9pOah
udFBp+afpYISGqhI4Sf0eQN7k59Yw6CusQPg7dlVC3VbqvfNj1PDon8CsahcDOUkWIBOlrTvBUWJ
9iU3D4g3rLvjtI4MyAu29KpwIrwmqoblhHhSyh54bGZB61TWyjIq0eMR7jpGbtAmMuH5ZX71Mx03
o/P5rNnGuuYjYyL3IEnQBJmJy479QRj+0o9VmrBG4xwEsikEhLddLty/njrZaZUdYEtSZVffLzFa
zujIZibGlqEV0lSaszfLrkI5N/Z70pNJLC7neqjxdzlQLVACRyXS+ZHjvWN8CVXFSh8CixetbuP9
Ficm2gJHkzaa095nWIkA13eYNJtdnN2vNOEdT2FXoELhs/Tz6WDOcth25fYhJajcRZyNfYt1VeUT
u0f+8luqrzzP6iZKDDf0Nys6nNBBCiwer46SYtZZCzzc1o0pBekCGjAAy6ZfpPgndwU3m0fXU/Rt
snhB3v4kYnL4Eg6eO4v2qMK9CCmxEWfqQG/Nak0KUgTxINaGT+jTL9PG+lQvW36vp69QD+HJqMq4
hkNXbJ6XJ4KsiIPPnVuJwUnYsc7SDs1/4nqejfA/RbvcGLqYOieoMUf0S5AZoILvaXM2t93SrWJr
oljzkfSqUq5MBbAk3rWFQ5RPJh+V+3crJkJFvx/t7XxaI/s1RAFc8Boi63K2TgATJAFBEwdRnL8G
p7G+sjcCYhy5zxgFP9KHC9JKDSw2uqgvp8Ih3dPzSOZMFrZyQEtjrqjTgY9twaJ9dN4PFobCZXiZ
XofPmgyDAzEPkDqkZXhzQYTjhfwuYVsyyMShtrsm7AIC1s3IVx5RLThgtrNG16HhIYTasDfLctby
SmSZXLuLf4XaLQsIiyl+IVTutRDmh4tpJpiia7C4n+yUv4F5yYQL+dHoODa8WJ5lt0nhZ9z0dipV
q8BMnValSffj1sw/d1qUOs/Onn9PqEySsbiGMLKc71z0/90PEFEXn3gTltrWHhawNpplyQwh6z02
uTm2idbCgjGC/jRd7/2si6ExweBQYDECllHzwJNTn8gzx706psdlClXOGW4zzgCIZou3xksgFCNA
KGciQvKGK7X/YE/u1qrmHQDo9iKNnMyYPI8duOT3mxisAz6kaDbN2Js6sSP4vgcc3dFjy1hqd3t6
UrwdriKF1TfoQaC7B4flicyes3a2Hd3a3KNEHJ8AQmr/+OVSPzyvHE4X+PrTU6IIX5TNPwce4EIr
36DloBgxFe9LIHzjVOh61ivCm/r9Ejk0IFJeSAIX9zvFD/Sb/R3XS49w9pKUtwLbUOiDqe5kW67R
hiQEKyJKEUKj/wMbrNer47YrrZb1Q0Z9qp6rDkfaMh9Rd1VFJjqcTqfSvkrC31KojX+bKgamrgtU
jWKjDr4rlDoW7z15BqRTgEdiwG2TclHo5IjLYlG0gjXxvl3wbjuPaxQqmHNjgfuSyFDOCpewqlfF
57w5cDpfik8fSSeZNfGcumFt8ISI0PZbyYBpem3EmThJy68P+588WWPHvZZfNr+cTlZyZX7cKZxw
5zU+bJvHvsgSni92U5+nDuAuSjxwl4Id/SuZhAdFW1y5bQ==
`protect end_protected
