../../../../../RTL/WG_dispatcher.vhd