../../../../../RTL/CU_instruction_dispatcher.vhd