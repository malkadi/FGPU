../../../../../VHDL_Files/V3/FGPU_definitions.vhd