../../../../../VHDL_Files/V3/CU_mem_cntrl.vhd