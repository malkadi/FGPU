../../../../../RTL/RTM.vhd