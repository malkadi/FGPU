../../../../../RTL/DSP48E1.vhd