`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
pg2rOGd/KTcwDdRn8tBeCboOFrKztHkBJKehCtG5izAvyAC/6VXlCu46n5x8UdzZVRb9oGGVlYYE
EPLaBek/5Q==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
E3aUffY75oUaxWz5xbDFJvSgNJuxEb/vF60QmK+TVvXUT4kO905WjogNo/4uayw+RecdY/ITxnbm
CtBn9t8q14n4cGdAAdXMMc4+mG6cUPf9YQmOBKWmQbz/D8tQvTYba5pqTk+7rNV8R3tZbO3QIGv/
/GW2wfn4eyTXlNeJKuY=

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
qktdtfJMime75Ja10jhweJniLuEomGBQKIRjLt4/DHxBPd4f5v6IMUBc/AAL18Le+q0RBAZI2XYg
LBy71Pq6DU6GKIEvb1CXCPbf5Gc0vUcJsgT463ap+c8wSl5XhDplpCFHmg2AhwRj9uZLrBunpyOo
emofTHryL0pAPlGSCzo=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
DlreQrg6ErB/t+GCadQbLa/zqOHNaBgF+9roqR+06XbPb8dCiQL0ZSQRMJaGVi66waqEoPiqnGl6
EuEPEwu4o46cAQIw9XVZwnXzXl1hqYIMIEXVCCMDJP1gNZ36RbtWoNOfCJ+SsMlYUjyFhCfKRvEG
z+U/P26U2lsXBAOo0xSAptE/xxHpIEJ6r5Ggeyi/UljN5bOvkRvML0+aFDAxXqyKDB3MH512oQUt
HogVgoz8pIEnRD86bmxVcQ5KMsxicfY8HJ+BytWdvviOTqDPh01oEWKMAwUljKONAsRJjmczbNuU
+U160KK6tvUtKviO6HGRHyfZEjfNoCG8fsGLQg==

`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
fMaL/MA4P7FVFo8k5xbhVzAYHxt1F0VSt16y3t+grpO0DCKNxMad+MI6JoNXUNsnJMjjWvrnbp08
CXvzRQrrPuxA1P8Gn0GJQCTsc7aEeiqrU7RKAsUwphxuQ+dp1YBpo5kfyK2UJM9Rqem9InrflA8j
qCQn5gY6ibJJZK1kX3sQ3tqzfcC1gNskNbkkmPOxJ7Rh3ucQB3d7xXO6tECKoTPUNnDmKUotkcuT
28w7DbbZi9mKw8Rx7b1+i3ZLvOVbrjTEEpdBjIMRn+7NFO7OUeTeTa7zKL7/JZLs0JrQniolvYlt
zutGAXsg6zBHMCDdn5O/QSyGAkOuF9U7eOFFLQ==

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
pGCOkKBVsmzN/NTvFyge3xNTD6qIl8MVQ1M+wFxHHZ0wE9rXiIt9vwLlnfk4CT6zfmKxBzuyhMmE
jialmhLvhJjc/I9lSWrYlcBBAD+BK0cPWeV0UtGynTZQqk3P0Ja8Ah9PgcIypiXysNFbkuALV11h
fTeI1UyErbWB9F9qXj+7NgCJKZ5zwSDDqzH0TfIg5ykflzX3o34qK9uvuLdy3hh1kD/HB6mcUXcz
qc2hzC0ZBQKni3lkq8LIguAz5qVDTUyOhrEPKar/mgn4CGBEsjY9VT0QLHk3O0CPeKo4ydaEzf9p
XbLY52GkzGdXT3er2G5hU6HFgylStOK2fRoGnQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 62080)
`protect data_block
0Ep/dM3ZqQUHqQzsv2G+GW7WITnW64fCiTvYuXdtypCMIcknbyV4WxtA11A6EaBlV0IdYbsbKbdV
TT+ISlFzdoRb2YYIKdugJnbVzofepiJ0UXeuV5gw2sXqYamCp2jJtOj2FIUh3bY7cKet7l6Tyjgd
jLqAc8WLAIXky7DZOs0hfggMXU8z5pj+CmSrqJPbhJidX8MCAccgLQgWe9l8uQxEpNM2lCN2+/pS
0MtB/1MuUlqocJbHv/Ln2j9nLEV23lBDsedvlGGvSXDt7+N5OpGqG3jaJ60vF7HRHFPYA2NSYEmk
RY1JDEuw+BuTqAVBbsjkzJddn1SDgC/DWyIKX8B0wTCJeLZ1xImKR1/jykxa2jr/ghl6aXn7u+o3
oK/cg/kg6dWgnjiRsUESa3luWONnXlbqAmY1xlx5HZ6l4YWoEo6sCtI1gWNpcyzzcVarr0a3hr0O
eZkyfcna6w0ATWbfj4J/0eK/TwxnuY4Pyajz4OIWRDTTnJE4xwgGwynZRV69+Nbp6d8w4Obms7s+
keoYCI3HZd2kwJnAIbc9iRLST5eS24kjn1D09BgDWF9csndI/qsW4TOreTTLsUEiAF9c9OgMQfSP
jQJL/niZLE+oUxadCnH473MojNZlFK5mrdJYgQf958MZwU86K+zaID6/GKPqoTpv7MlxS/afNvot
w/AHR0LGn2NQhuWtNayA/bSfUodOZzstuOK3F3xcW/UU00tJaB41tL+shZNtHgUu3Xm2ggv2WU8h
2HsBGSGS3G0gGd/YUfTrPpRbeOlvRrollHqsVzPM75yyLjwMRcXvcvLmrKlXuGNiDsqGC3netSSj
E3dzDujhc847D/1H0255D+TzvrdXswwLDTJ1NSCS3gLVOplV1vN9AZYCMLhl6hH4GTQf/M3G5PMe
KbgKQUePjwJMgaShbZGm3Maypuhng0OkITnbS463+gfF76UoqIiisNQ7LFpWWqWNiuRKrRudddc0
Hzy4czHIGlVPEKILtIvg9OKnlJzZgUe/aZ+605k/J6zPyQcrhLhK24Y/OWMcK/8z5Stu7a4TiHuR
DdUi2m5W+hxbSXh7Y3MdFOya4ylVCy5IeWTiYC/WJynvTF7dP69z5/FUbGOC8LYWK22ids5eteOz
Rhs26VMVEz1zDmbIObEq/WFHO6AMSvgPha/na6nwwQOG76JcdRsRxdm7+2qnuFqyPT0A7ai4rQoq
X0CoiXB4XL4ZTAIcVEUPPN1aV2PB9RfABDKyeM8RuWFwqJcv4rDnSYrwPWGgKl/jaSu3IqiiQAFC
olX4EQzNW6LQy64as0nso2UqgpUtWj1NyQVXWO4C7pL3L5/lav+ZrFY/cUhOfOWtfYPvS/Viv6uF
iX7FRyXMpFjnhLfSEPIEn/t/bWDq/WUDOjGu4I0t8FS0UEWcoLFrKnSfLkaoNMty26OZP5Yu5DA1
DgEGdprVQaC/Lcl6fKN8dfb2GT2mXPzalxWRbckXT94OJDufZCmUYzA/7p1d8sSM/yVhYPBJ6uSo
lxiSs0V9puM6OPsRmeXYjWp56FqhB+rtI+Qx62vRXYyco5dLqRMTeNojAt601fJFuuXmKnwU377M
Kj88MvnakZVO2+ltCy9T38JVX4/TSIao/eKEnX8OCzMqUoQCuuR8BHXvPfax1WAAwSEm7Tx+dgOS
WjGdASFRv73T/HbNKIklj4X+xje03jBWiC09oXgPUggfxy2ekaeVh2kmSobkqZ5Bt7w+nL9zEvP2
wOMWf5xNPoGOavWkKvA+r0MN4KaChcu/GeluOvOuUqt5Nz5267E6oZMLI5oB9OytgeGwdAbdoklf
EEkXChYb+QDPKcugtcOeLIMuvrdnnEjpnttbVAwyJtbNBfCy7NMUkjFhQY6RGYrnQKQCpRspZaBU
vgk1tpWU7uNcYedcVZ0g8EIq8nNPIwwZjCE9IBGetIzPRRz5MtNvbPXV4CvVrg3w2S+MToCoXMrd
/B3Gu5sNw9FMDIfbiJth03NxmPvuVNF4mevK4E2C7cWGnWm5PzAAqMpfBYwZLfxyqVy2EKKkIAYA
akH4/AZe7pPxqWKjtbeMZArMdp7QUf/qK/LoOFZk2H8a7N+lxiYq0iD0VTauPUpoe0kqif3sc3Kb
oL2hog1phsj3hKyPC1kE7/YslD3G70Jx5J4ybLZjYv09RH6FPr/+kzGghsJIzSaxAhZoNrSyPbXd
UqCWQSUiVGUbD3tVfXGTD1p1nvE7iLYnSGuT9NtVb65qzvZwekqfi6SfjiYIHDqmuLKKMHulSlIA
QoGrHUCJ+Ka2o4ZAH1OVpCIEP7JgJv1/ZZrqrY+6Nx79yDS1HaaT7cwEFqeF5cSWCu0IBtr+jvaA
PDS3zivMfXZ/JFpjGLnzHERK1vPGysvcrt1DCdHX+Os2/9cBuShZw+8gHwR9qUKWatCzTNXPEXqN
wQfwoNmf6XZ9K8bZUHpA+jsafblhXs07uO+2YjL2w9tsXabajejXCQTSVz/XcPOqRTYKHsp3yba/
LG2q0jvSWTeKFfrBxx5HGNAimthSbfhEMWLMdX8lsE9Zs4XiRxs89i+1gBC+FWJ49ai+pg8poGMF
JcaoO8ceI0cPOsnpvV3qoqFPBqGtsraEGusZZqugi6lJEG240PIkRhVgmlMGJc8T/ULJtfJEKA17
ptq9QmtxEZY+d1VjyMcYNtv3+1yWlKizOJt0RUbrIARrjB/V+thr+EA3pA10EC4RuD37txCVEXmO
UFLX3nMzwB0EoAMHFuw+AkwTkraNxAzxwELHmUiPI5b2PKdfNJcEaNZGHFcGyw5M6jAfGFLIHmJP
PjxBbFe7JqsYnpS311DW9bt/GTqupWF8NXpPucMF4EMFGb8i/Szvf5ZcHQ8JB1P/kXB/LX5EY6Nc
SrDd2FFwpUP5ffWs89rx/q1O89jqMSlLxJim2eaWKFvzqPyAOekK5dXEhJ93jvogco0X8JQ7c0WD
00KhR5Y6QomGB4Vex6R3CgLrENWf5n9AUzZ8Wc96P2yYDP9io5L8iZlsDi/7Fo+cpgzjfLykYZXG
vUUieClaIQV5taMag1w1D1ixS1TB8BhwXPZHIAdleOJoB7cciKGkc0zWZUPArsfM+vZVVzk7Dhxc
hJWeLjmwoOOSj+IDDrhEmKO3PpqlAnxwHNP8S41ML6WlXgBe5esA3TFENliPpyuKp1sotrfad/fW
36eRqrCknjbohWIslIuvjDkP/E6es0NzQiGVWvct9KoQ/qlMdOyPJImbWsbZa0gx4CF/sWjQ+LG3
vSNU7FEoSOF7FYMbTmdTAlOeO2AmYlwDhCjwCmlCfiF2PmtOlqz4fO52RJGDpk+UVD8nEcj9MR+R
QxUVQ9E/n4CykDBjzTyAX0vhKKmiv9BP4y1PCwi5s81bhvs6SFcuyUDtEkoOmGG645TIe4NPqq5v
Lvn5Cn1OAGrYLtdKNpkKRSSUgTi0zgv/DNMDdBJQNEVpwNKhIxnSId5668m45eSgZc3F7YDkLfzZ
uZCedHFN4+bJAIJYTVIzoVpCtHISmGwqsx4z1iQPIz7v6JkfsWXQ0Kzdk/dyxrvCw6urzfeRHO9J
zAIVNsdhjW18KXYEA2QFhOX2fT1LHZ0fL8YccCJnJqJSCNtuwKl1st8ezvBnY81iX12bQloT77dz
hm5yjfxlGH36+EmVC15dgpgL8oMOwjd19RNvakeyP4ux0mFa81DvnY2IqQP/WgXhLrmziwmWtpCV
bHL7VSb+5x8Ch/ZQRBzn9ZMLqrlkFczGsc+AWEUyU56C+0faEIm4FpMbVAJFjE+krihGdsuA+xLe
hHmDK5WbiaznfeoQ5knS7OAj4Aq6I+fIBAvw90Cdo/lpLtghOlyyvapstq6R2eEjrErjeB27qcdB
rvjDnsLTC3GqmAkbcYHsh7Dzr9luv2pulcjWh4gF+KrQkRMtxa+amLWnO3FiDkBZZCYu8yi5HO0B
yUP6tvwQ9utsek06clegmRER5ai3bq5iFaHp7UGY+U13v6/G9TLZd2+4OGTh1fA48oVae9nlmY0s
B3wATBxFPp74j89LGd6tQ6XsrKk4Y3y6rK1iFZgk7qgujV3uwMjXmMyjTS7Q7MUTb62VkILDzVbL
J3gzEbkvxmyYxPX2YMyXsVZSjy3/4Viaaj86wD0mPuEhOrCckqRFyFXW+dEpXOKRgFPb/n0MIgAA
to/kWLwzJFoRmEpS/wvk4DUj9de7xtg70f8osgwPjbzzWkYNYMbvLKZBUE+fOkjOwEuBR9NUAPed
zQanKjWFsmpulPCjdPC9ihmDw1I1wvQ8ITdilJViNhEOyMwq47sDaiHMSVAu9nfdL5axbemQp7w5
vIE8sFFmERd6Owl+AqXMGbzRFEVfmCc152ywicZTZcDu2kQ7UbGnwUgHhBcYatvbCJF+APfw2Qmn
pGrrgcqqcp4epMVLTzjUByq1vFvz7ivENdQf+DLsJXTcaYoUqRFCS6deQe/YVB06HXYOyiu9cKgz
Vaz2BiR6ru5VqI2n8PI2jZZXd3o1eu3Dez7xlLUCVKUBXxkVU6kTQ9jIrT9iqkJqJurgxzDpzn9D
5QUxQiYpySFILORSUSIcHGDH5Vv0vifuf/nqYZhkbWgtaMWV4dExjgFykuZ9xddQDRchc1yLYLc7
qQYYx4ZOMYahw1hnD7rUV6PVV/c+j0KRiB08dRB55MFBFHrmYHIAzSeyQQ81OeTdpXYpTgZLPeY8
uzAAonCg5kkqW+/yPm5U7Uk2+OdPBYxJLREtVKNIy75DwDpTEkUkMEgdbx+IuEffuhzKjcUoAGoF
qGSjm+OGmINM07ByrBajRf8rgnixTC5fkQrbY6FwyQA741NR+U7/csYhzwqsvixe+ozwoGuqOJco
uxX/zrd8iYLJAhR77dVn1PGRZNAnxZVvuDR5BpeUkELgur+hn5G5TDAxqSp0/ydpyLEzkDASG4Kx
WwYUV4YLMael/Gnjquv9c+J+1XCGIdLGz1QIdsQhySyBj7qVQvAU3aRYkT9V4yvzHRNqMEgRmCWx
AGdvqZCqrxF6PuFSGhnos2s1U90BRD7EiSpM9o0rQx3wopFUR0Vlr6HALNu3W1CzAY2nPO1LS5Xa
i1b42gfr8YDDyt4DxebZTGvZu7K+wFv7aI6hFdH97KQVzQXb1bmZaPHeA2HGi/VJz6TWFNZe1phz
TAbLdPSwBWXHLpXxH13ZB1J3+EU7u8hzq1iON1tvsUL/1rSHVasPHb2BmhlWb25g5wWtfBJfTMwu
3JehFkRmuJgav6I7hLtALeCldD5ReZ58s36z2ylyHrI/Vu5k6p72fMhANep1oboJxQK6+qDpBuWi
sbY5shSabeC8t4zBQNIcx9LnEaCbyilD2IQffuGdJQzactEjT9rkIhhL8PAuXmfsmqc8QwYV9R/f
efztWaLlLTgmq/xCVW3z2UVkFZkmXJWQqlkYh5/tyk1UOiRvqIPcNpSCXOmzzzEPWMXKRNRMbm9Z
UosPgaWNuhKdejXFjcLzwkWLVy8Dmng9Q6S8q0FH1PWmxZADKFPDRLeeADlunSZrWpoaP2ko0P2b
26lr+u0GOlvkJkEgp/XvzU0PNIYf4eEMF0UmxkX/ukiiLsp7tNj86nNL3s0esVPSWWRsCFSyrc8o
U2PP6fpkRZAwXLorfFOQBdNPjU47EkHsWPKGfUuQQKys8Cn+5SepdhSRtvH02eWym5gOzNrqQPxH
/LH2p9C1R7UZ1oO2NAlJp7pYGSrctM1SaZpjWpj6oT17g2tN5ijYGgDEl9p8aSLxDA52HnG19bEq
LwfwU7K2ZYhbct3mZOVhL5sY+ataAD5+nTQ2DhiGSky1AIW5c9A+Dkg0/tirKlMRCMtjeG1VKqch
MtgvyJdcqvomPde7xVcBDej+lBbk4xA4O+ZEAg6jGrkNAb4onHGIkAbWa4FWJzkOJxpJCnj8Ui/R
GPau0DGgkRShFoe0f1VybVBnt9c1gNUj15KVnS7a/R1xB7yf5jzeLRaWJbluBzaf8Nv/Gv04ThJQ
7/YPzUyZ/mBdjUS/XhPslbHVG6yw3JtCMwREhJqjmxiNQsEyaC2gFfEx7VeD2pIPawqQLzHRrGtv
RsB4gefXf50kfvoVkaFZKF4sCuTVYBg4kd6hUi0CsenI18LSihnsYd3GQ6H6AYYmQXfZPCgzxLlO
V17Jes0rKTpvO/w3gW657c5m8Xiw2/IXCtBFq+0YKFZsFX8BUMKR9drMW7k6tORB2Xv0TcMgfzDd
x2wnXKf5myIbEceWWIE8nVotI2QpY5Kmw7RxS5VLoe9hRz/3dbMBx+iGvduCmpBcu/E6DnQU4Zd8
oGH5SKg/vQmjtOUACj8HQCX/3q77p9cKfdr0XbTX2S6M2I7UdOk/2nZkb/aDHopdgl4yWhBvxAXG
c+hDqJV+lRRmT2vcPB/XTOEK5NdyiiNWqcrRhtJW+58ooSREdyNnySq8hMIexv9rmg7sIEBRmzbI
U6LykjFxLR3zzElaVnbuDlsg8va4lqEWSPd0kJcbCRDoAi6jzrDXFMzCAd1UiYD41C5Bm7Lol3Cm
4GnnnBOVTo4s3pc8MRsjGX6bymCsWxjmkpttQMgjPq2nIM/E4j3X9sLAS4xNkyKjwnf6xxTiSi1O
AoV+NybDL9gHMNGiI6I+c/O8ELuV39DlJqrwnfbpsZRz8lNqcDDfsBBClfbjEegrbmPSFBvhWBZx
AQVvq5bA6O46MAOADC5hPeXjHOpHnbHgkBy/dKDreik5vuplHfSyLVy5A1rCAbWUEzXpb6EC4xdk
/ntxpZlx5rGvJuZN8cFG/3sdBN0FzDbnF9h+rXre0bkknp/WZkSl9uYBUctTP6a6VP+F+4ra3nHc
nZgsWgGWnaCRXIMVhHkFGHETWpZzP/WsML9pb5FryOjQjZnPJcSLJ/NQvUeYGB0821QcRA3DfM/x
pYKlz9Ulg9Ef3f8/Zr90uqoBrhucMqBkXncYWBQaxG5ghKI/jaufXZ9APii9C658hWNxHxsADaNI
Rhe0eOHJZn1PXhj3p671l/ZGfuxewPEQLnHcE3OWQnp5AiV4EzYhJR75DUWZ0jBAhSFP0SxbFqhR
tICvWJJj9Yi+s4PoHQ1Lql+hgkdBcptM8igfRnZ1TdgV827/cCYUte0n9OcLbeO4NmIFde80ZbkZ
pIjGhK+hpxurrcPRhQwdfSAc+N61AjvUpTm8+2c8duyYDV7Rbd0VvMgBKZO8xBdrSWUBFVltqy8D
6nwug5w30Rv+JEOC6G+BsF7Z4MlFO32T/lLcfDMKtHnDBvV24AKKb9Osk5YFHM17kUFrz8n7VhIQ
JQ4Vzlw/8I5W2FgEEBMqLvTvowtAQF/Px6T+zpkTH4sWc5qk+KG7w1neZSWqdw9Olo1rqTd0onAU
0073oMmN3Ef9WC1A+wzp+SR2y27fUGNlp5mccyJ6tACTUzI8SZFhrTp4WT43Q9dKZLkdX5NDFHnW
04Px4lI+WLoY4gFym82NwkCKWWTykiahb/QqFk0PrLYpED/tDUJ9Mt67hkUvg3ZmbxK/quPn0p3W
QEws2p7anPCoTNmf4xiv4fpHhtkryIhFYTcggxbkiI5jnc0LKhghHa9KVniOIBZpDBZ5+RT4fd1q
e5lmsTwwsmwUt8EDPfkIWjMjOWML5js7xJ6IVtX33Is7tZWnjn2DIZYPPo08nOjQ66sLjwkAkzc+
6hAbLdiL9VV+PMoFANzF/hTWJ14hcsirAO1/q7YoRa6DfWGABA7fzekKd0PpnK9JRNKdSlagoHy+
6NPWfGaO8brogLVgsWjBZonO/yLnXZ20AT3foz8MhzErdQqUtdfF4royrtR+YCr8mQwYS+IFAGOJ
6DFM+aQa7MEC1YgV5Rrra59FrEXZc2RDjcukvIDiuI8BeZygARAmtdZXOhcD+Kubyt2AfkazA6qO
vksXTORQAMP/XkSjcLqbwB7HB8LNQ+5FxUkwPa8ehY6pDevT8V2YRweD9Qdq3uyj9jYuuSXf+4fW
1YIAn0ZVlEK1EfPChAjdfSgWkLSeilyzYXBZAUo5P4pO5gu/buXgWKlGE0Dvy4h5eGSuYayNwxHN
cB867gPupNVlAIdRxPYximC7+wn1tH/P/LHz6y95K7LLPkOBnOEBHXnY/tPyd/HfsX9fyMh4ZqXh
Yb7K8JaeYYS36LZEE/k7MU0RUyB737lpMJdOESf/0KZQSyL0RXA8QaB7qAz+paM7xFdB4LJx+bGG
yt80qsnlcPigRRY3NjWBEwMHRVNnxIqO1Sf2r/VIkA1b6Ao6YsHAQgNrPpmUptUWdw7xEtn1LkTx
pO49Pbf2O5xfCO5PhNTh12tDwF/IITsx4iFYQEq+DQSjI/fm/fqA6Cj1MdolYZXxQTya5HBXybKX
PKGtnnAy+xHTftdK8EqQP5pyDgiaZ7CkDosJb302O30thIbUkSZF/M4KI4o0fZF0vj6cRm/NhnsF
HKnbXiHKXNKfj81o3yX5gUtFkYMe81YYsVlRGqVXO2U4LAlavTa5lDSRa/DdJiZgecc+j8gxRcbC
IibqBLlgL8IJI4OfZ3xj6aaxxzHzcSd1x8mWZsmbba0crsLSEDNZ0a1NBHO1pd0HldRli5CZ0We3
kykiKyl0vyvZWbMq+M0pov8lEGCNM4QRkwArzL05Ez9twVoUp3UwfPfUBft58tILNJ15bIJbFih8
CUrENOLHdvit90uNf0i4gQMxd+CGcZdvnxzEL39XYN2AH7navat8KJCq34yls8mnHitz3O2Bn+q8
5Y/v9uRSp1eWY2hSXMEuSeiNQO5wT1eirkNCIMlq1qI1/JkT8kIT22JEnguFN3SeKT9FssT/eUPs
E9eomgI8XdZjqAaLZW/4ezBgVbNpVCgYv5mLCkySYwiLzKfl44KW+s5TMd6MIlnj3L5fe8X4KhBL
4pnJRi332F3wuShnE8bh/ogThuuuRRufY6QwHUycNjWaJBgLlE0xM+Cxd9kO9tYNB0TPPcs53wT/
vRj3QOUDilKAgaroE84xVxWU05WDEnGxR3idgfZrPSmGLh06GR8TK4rCwSo2hZdkIdsE9lA4+w7h
qTJrA24nCJOviyFAFxPPb9zvFG4+uXKteJdXRyRY781NAvI7bEtM4GQLEw+PvbX9V6T2Bfv9QWCh
8PVuUStQ25Fo5Tk6u50pMBbylr9IYeJslotIgLxgXiK+jD05IZiBT/JrRHCGYGlq9xCF6pPaUExJ
/o1KjCY/2MH+TVJtUT0it3URTN/rXjmTMiLqQdab2wrip3R07EAGqqHETOHduuU9ZU+eqUEKINyu
PKJWLnu1ywT8aZSrK0OWThJKe7w51GZBG6uus63e7Skprq7zBVEgN6odrR/Zjdpd8OXoZRIt53Ga
gnX/fhrbFyK0mkfBzCyBpeXroz4w3PGbfNjjx9kfZuLHc3KN+OpHCHTUyaODxCj7LW9m4nX7ZsUP
4AueLgsx4ceOkeQ9u3ji/DcpuxRs7SG6jkoaRKNbza8OSHXkDX04VpyEJhcGKBK6owfVgh0OwgS8
I26ZqibdOwYmG7Apl75xYW21fOLB/g/0/XbS3631HhGFCsHYvh3FeAEyd1MNuBFmYQoKtGIkRvEE
51tTtXpPxNA+r7S9/HIPqfLtYN4RQ6PjxjOkW0kwTucaZn/NfT/Z+4oB0R0ge0LAqvvB8irfX5xl
aBOjcKPBdC6OxOyjDz/RKuddA5gSV4vxQrN2Vtj4dFJZULuS4oO5gB7+vOomsSftj9zpEtCaU+/w
cIhRfI/waz8+IlNaAcWHb/nsl2KaeZG6kSSJOCr+OKJllcvZAwd2dcO6s0pL2r4q1zzFznxGm5Zn
t1yC9h+UxguNzF9MQPKSvaYKIx3WN1+loYiINStFWiGYf5HkQ+0Gseujwn4hCzAgGS7tn8FNRoPB
nP1w0bmjRIixkrG5DcGfTPd7gEtQughcDyeSE0JKCPNnB1qPdp0h78j5vL5HA346Qi6Ff49rTMkX
137csfxR3IgcWjg1mvI0785fnTXoeBR5wFAtlzEVvwmyJFYTMQfPjsCTLq+OxQZgNyjHIfvfb5rr
ZJHKm/9lJCD+J7QgdRyVTvDhaJ2aGvLkDdinXDG5VuNO1+gl8NOf9rwjOOpbaiUttPKd2uyMTy/B
DLp/+P8NkrhseqSmAGqprxpNLGIr6B83CNASst4KTIg3H2dxAnFzuYDJxh6XyBiuuI4lJbIUIucs
9lo3Y16Ypb/wQpOAOrhVaGxALgCYOwjr/W6Clju+yhK2B1iijnzgcLhEQUlTaLZVh1bu3eVfn1O/
BrAZ2R40xdxIrQGBHk2u9f4UMQJkzarVpni1RB0sTE48VdjtLkhV3x5EkSAtXP6wLgqArLH0v/ut
djF0wOtx9o68D+zPZHyyU0M0g8vMy+VEdWnhCr6qe3D4wdO0G5V2gfchOrQzwnGzxev51p/iAZLI
KIM5aNoNp8Ciu2me44PdtG3JasUHPWLm4RkcvQZosno/BAYT1RVkjHzvgBQLtarMqwHcOq5erC+i
shyu4g+uCFRWPDiNsDvwEOV9sUthhodEiwYtqlxsGYV9jkM9aLdKNgfJP8R8kNFUcgjMR/dCj1fV
TvLc+7kH22YWwOb9KKmxtWY315GKQlrtT5cK6IVT//rQNLtDAOD7rXlNgD24SM8FMNU9OQAmy7+Q
AfIJl5p+YdGubfycp4bri0qK3n/W5PS16L52gyHhg12tD6Ct1dL8q5YFPNqqHF83vXUi+fueXvWc
Zcm4nRbg1hunVxOzBqkrqGAH9VO0IZ1uXEjP1Dugmi+2DZ/cDD4PsamvgK6hAzJh0NV1VnVGEeCt
8pY1QP8426gWd03MNmINkJL0ZsHsiPcOBGH8rJJ8WC3yk81Hp/bBgAWG2r0BSEyT4IWJ0HYJ9s4C
m/3J7VcZOnK+HNa4B1CtYELfMGOQANpoZYdcg6Q7b0NDRdOCjs3SVIJ1a/WegFfUqiUH7i4dyfm1
Mpp+hp3+f+rXCKwWYYyVVkTJ3GPh/Sx4kpYEsWyMmuC3m2H1HlyWSdYPDRLSHbCINSXYWN5UbYMu
OzEG5xRN/jVoJW0zBSEDNQxcEz016dxkEq0YNKlv91qXFVDwqJLMitv1wwsNKCn8bteOqNjMXk+a
VFjYaIlOiRFcOD7+cuK6tLppiOQXe1F/IfurMHWZ3jwkSIZIjpJT/Gpj61cFIqq//6lyV7ueFazo
38rwGwiGb4FUz5MG1U3LJWq4zZtCsE8OS2h+70ThTjNX3uuME744AOT7NiMFKLPb/1MeiPhVQaT+
zk5s7fI9gG1/bZzd5qCOfdxLj6DCbX/Co2w7/uw68RO3PGfMOEKAGdu1RPT54VcxBvp/zP8IFD6W
81m50s3sU7p0der+MXdwdF14SirZ9iVVidt91ehdpenEK9xgX58tE8hljmhjXP5NwBUcmUG8xClP
sYyd2nIRoOzru4qagzBIHQF3YE8+/SxqW/iw1JUWPRiXWAfWkuCewAjdBtdg8uJgHEbr6XcDOGiH
2XAafzYhDgrT0QPpYyDHLQJcwxdafRN9/fumM3WEdWjCoiAJT0LkOaB3x8VRhPlm9RDuRqKgYVzN
zcILalBTcwkvZc04yxF2+iPZhKGxXEvGO4XGM5gYSKKuEOFFKCQQS10jvbcVLxn6ZSn5YX8ih3A9
TgGheZA7i6cMfxVNcpRh+xnd2GzCqFOW95ckxcowe3GbUCuJ81wIRf7zxDLzDrh8KHnxc50/jCHC
pADhV0u2fbW2vyTci/pc9rCewI8ULSGPMg7nCeQE6mWGLpi3JWsBsvhyPDXLdzK7czC1Rokf+D8I
etsYZKH/FxxAcQVZV/OyhyveKPWoHTy9JEZFSvqWCmLFCLFXaZzDq8wgTX0kZ60uZQS5wAyuJrbV
txb861gfv/fDoT7uQRn8e/1B9H50ggv6TWcALwY9v82xhFRGeA2Sg9QBw+DV7zWCT+WpyjUgxm5l
kRnNhbG7PzJviREk3kqBU9LytI+ziTJXmpI9H0G95OnXb741kRfKd3PvBxQzyrEMA7ae654kNLia
OTWCn4acMvJmLOd2PW6RYnCpKsvkql20+Mf0dq76YfytKypp3INcVLh/3yE8N3ZR6HVJ/wrjYzCG
PTaGSiumdoZODdohMsvTmW37hgF/S0rVzV0r2pWzpqe8iAfzoCNKb0UlcPg36QxuB+EzRMbKj25+
WXaQ6hX3YZXMFBPdd9NKrQStUWCfvnWj7Qz9Dvv2DS77GWx8mF6SSZ24iO/O7G3a7dJIN0gOmheF
jcpmTBUsY/zAUSid8nfM/Fvs3azlWqXT93R5LPGjRo4fvnOz096G3ZDv5aqrqZKdZcA2n5N6SnOh
Z5ZihHWWc3wP/MKmXabfywmFQbf4kEONKmvj8h43Zzha3Iiso/p/+UtmEKtHz0opHDrd3UANUYje
hjmjLn4MzXIJZuQB1SMIGNLYD9Eggks1E2popx3vOim/WCozIo5TNRJMypditd76oypfK98XdcXo
GJCQOZTrLe8c1GAabtcsHIoVs7YkBsd42sR4iC45jLbPzv78MgKt0/Ox9vOMFY3Jd+P0TpyCY/Qn
2oGTqGYQ+7jlKnYix/1JOEzjX76DZRvn0GrZ2N6u0uVd5fQFVvAsnmgqbm3yIt3jaa1zBVHUM44n
RqIkg8STbGWl195v4Ei44fTkukvQ3SbzZf3wUxV1tJhNFPDtDEv0GgfxcWKooVB5pn+IYSr3b8VB
p5mVYKr/ybFl2UXlp63j7VU9JW4OI2TxDzKJN5Z+2ZuujnWha+HT2YfoQl0UCl8euXw4XTXkTO1L
QaQg3saJ75KhtyRZ/pR3t22jzOewkXxNeJdNwSz++gmv2dPtN6RR9/qL3PowSC3xyfVPoFjCvMyz
UDtVO3n6W2pMvPxKRgXcjJE+4dg3H2U3Ng6WL3UT6pGlaI8k1n+kOjuInOBm6bralftVuJuvUm1H
cSXTOiMJcHJCvIXIZD9ZtJDuR0vCYIBrrrjbN04VNjeIack6XUIPnO7uPzK6HtA/9SncSQ6d0oid
VG5sRnCymzRq2CdV76X3I+gs+lgwjQH8cb0tFRVhxHgII3WSHeeBktxLRX/DejtQDdGNwbSlTrZ+
ch2/vdF5yZrQcA+DF04lT7x9mZmICsxBZoRNIUtyqFulLJTsJmRzDS1WxzPCrZY5zRFCLItlNMT2
v4SzRHHA3FLFnvjzLGeI6zJq8kF2iSykpVfc9/Ci9om+zEH1Hf4n8ILbRp+6ilB5aQ+37HLHPw8j
DjR239xUvlyDTGNyuKZkXK6u0wGRkg/LvHzL8oTuXDRpLjLj64xdHeB2YIqeG33y5Jk4mZ6vKQ31
wiUhw7r103JaQUW+oI2Cqbuy5sEVi/aCUPS16BActKWPOZt0yotk0h0IUeyc/mxRWL08FcLPmj9Q
swXh5i4+YlJXmv8vCOTI2I6HB/1FVQcuSlbicIMG9oFqvCNhcrzccnYM5kgwCXoBP+Sn9TYIIJ0x
DyxsD+3LyAH0PRVveJlbeeJ8Hd02cFLH1LmN0zaLZ0/7DehFi9CuRHSviGuquGR7RJHAlVmMvlRQ
E/IWnpjpHjA//IFEUce6qFJ8jaAUwccy9QjycKlEw2iOFTb5LJ9D4QqD7qalTFlnAxP6nPeMezCC
zu4FNBhRY09YE0IG/BLtLrHwsVQxz7K5djqicoYG5JlfWAjgIRnWhEUo+yHos8qtpfbka4Q99a4q
5LeMemnT73u5fWGRoiClB1TFLfw/WgHIHOqFkKgJuljoFwQaWJRKHQmsS3XNP51wxQH5Ldxs/igv
xFINaT6M3XoOyjWqxO0Y0LSa7c9/Ec2RDe9H+cRcaeQ3U7m9ISuxPy+KkOWVOXbLGvJ8eZfkjMXy
2tMUI3Q/zY5fObTr1wsM7KfKASvpyAi3eiNxV8PIinoDer5FavSn24tSnweGkSOPF+aVtkn7UOCJ
SdKwVAXOZaTgxh/GbMJEyzo6EoKDFJ7rYVC/zFNeGsSPqIzQo8WrkHy7ejnk3LydLK0EXQz+1j/8
BY/NoYfkGF4YWJzLZD98O7FH7h9NXP4S2eH/W18JxCQI9Dz4x60uC1dk7iZWn+kXsT+3Kl6GhT59
cXMsUeMTQpg1Ss9BDd9qCLwFPn4qnegHruXM8EdFMhJuTgOwxpWFRZ0EFNk1nbNds9Vs3k0YDRgw
vIOrYefAsvaWvXcFni0A0rvdqN51DCNoOlrjwsLXC5O6zQWtP/l75DMImHDjnjXHO8I1oYkoHJj8
oK+ldzcqpTfOp7tfd7BAbXXunHyPRs/dhBM60j6jUiRImqcAerjgohWYyK2xQt+kmvKTRGLZoQqt
6c4QQdqEEr39v+K/9k/3FUUpZVR/rnrYnoMSDPc0oXj7wVL1E2bTjC0uPWj8QqnG0Ye/t1OfvTY6
5udRDjVFk0gMCnmlir1z3KI+o5gcbvvxp+/nK0XEwpgzMuTL9vWQ1PVpUPtgbs+KZGCZpeH2FVzZ
EX019Qsmu4Bu8Iy/Z32EaVW0Hs5hHTyvTh/jaCEdGYmPtOCpcpkr+Ffg9DyEKGfbfPCzoTQLl93p
4+iActdht9CZlSUNRC0EzeXJzMU07+wvon/s53MK1Qhyxf/wMiYl+6S/rRxo5nQ2z+tsMFmETaKd
AA9VkcPCtFddgK6roPFKlc8X3PYKkrb9Kt4PSu5vrTz9yOVfnBrSE3fpBD1fT8Y+dQ7mQEWI+NP8
yNG/dEd6wLgy7lA31Xwk4SPwBOc32BSNyggAho8Pps8oQYtiLlBQpi3OGRjG9ShOsEV0myPLa6jb
qiI9Qks+aVwxquao2dgCNoGNOSLuUCa1oyUstrjjOrKaOPLIGFo2x5WeGkCuo95p1GgYpFkldWX5
rSZarXi70XwjBAYnZILedRx9GGnrzsjBE6/1bjJnJtc9Ig/4bm1MpeoYLSZt/nof4kYgJ+An0OXs
GJt2usg9B4BxVfnlH7jYT5+GRH4FpCdoTsC1xIF3f7Zi+lELaQNKAZC3X+XT2I1puONGp36vHljz
I6pqyiGf+pRW3C28OxKKyeGWwWUh4ynMSP5ziJF4tsZGaUreZYkVr/DgBvv64O7XWiIImyHMqToE
yttITyee4eSC11rkOhNgR4gUOfJ9n+/hp6kskUI5h5UWUQtF+eUwPDeFhr04l50CunLvC0AuSEd3
uDS/uh5HoGIzJX2BZDcGR+PeXFf8viFAHDMcqzg6q++JPhC+Pfsy3gR/PzbfiXbvZ+mRMgb79G0u
/P733ub/hZk55G+MXFz6DWZCUnICZtN97sA0VV6Ega/aEVkI1pFEM9Bf5mumT0M1OUlm8fVj6HR2
46FXZyrwZgxPf1qeGgHScTXnLAgnFPguxZ0Sz4UfIYiNI1Bm+u7tPeb88jyxhZU9cboYcAa+5ePf
copx/bf+iUENTcNei/VOmZYNvC0nk4FcWpkMGEHrAX3kBOq9OeRkjV2p7DRElMhB7ZEUBYJJXGZk
Mcd+Sgl8lQfC6iSp/vPxzvxWg6Pynvz4B9w759/6WkXzAZzSjBN3RI18mOGe9RcqFHaxXij2KvZg
jmq5rfTJhROuVKstbtxfr1RdSJv1z0F81oOoOfQs3PUNAvy+Jsqtq65lhDIW1eXg9J5qbM9515s4
ua1ietWZC0xmPx3gd3uDIdabmILEwUbN9DhNXNAzx4zjLBq6qLYlO9Cw5JmTa67+/f9Ji0l/OqWi
MPw1NIOnGnWAaRbUO75yGmpEEvQEy037V0WNg+gt96Ztk+XAB/Ag9swF1Sau/nQ5pDW6Ai581NUV
6DkY2rkQBfbU7I7sgl6+ZW0o5p1twSg1mwvqCRDLvDHIZNaV05PGhmmuVpXdgwdvAXiVp8rGMvH7
W3gC6oCTN8QVy4mx7+uGO+bH3krZUUrN1/b35p+vsXqfSqwsH6zKLXtH49aTtY658IFzaWIjAd1M
QGGK8s89rlSrQur+aStWb44ZXXSFUwYLfoLALRpAPB6R0XujCVKT6s1s45emfrxXRsRLNuxwu1St
M0D41plcmQ0owdYVzfin4Kto1jP8Q/9b9jrtU0alHL4TLQuLtj+n2l3yrzC9MehdE/f6hWjDqSbE
JaIbLjmyScdW3ouYYPk5SV3LQ68YgSGkOE4+48zPtgjcWwtXVYecstupFeyZyTBh5WNDf/LIu8+B
qKnU6ZJDnfaX62npRKqqJT3DjUnjz/9R7Di/SWLal6UCyFIFZJQzp2tpMfKG4BgAJIju1EIV+8v0
LUt46rZx3ZXwq0y4mh2dFWrAmrt41KsOzsMN1/lf7tF5QZu1xSNQl8qE4Qh0elSAq0UC7GYMWdDM
YllabUIIHSfhVy45YK8T4Yek1r2VnvRNTDTq4vVbvuQ/DrKgOlhhT5YB6pZgEhOyt+mvrDMFpMy3
ngnJ94oC7tudr7WILWvvWlGX3nrE3otKpe0aD9h8c0i3sj2hTnx9zghUjIVGWCsKFoEtj9VW/AGv
z2BeKvtICp509PAYch/gq7vphsRNjgce7RSI9FCapaMT8k9lss7Y53OFy7onOOXRHLEelBg53pkX
rXjRnSNSrHin+roo09N1Q5ryVSqgiKLPOFEM9hXOXz1o2duTsQV8wveRkbyQ+92qHsFEuxExDCgj
fwLv4XDhddIonvdW+1cT6TLUMxZY5Fs/n5f5wQ/6ZZMMZQr0Z8Aj5O5GBcOgiv+IAkxNT7CKEU9c
J1FftRekHlnfPfBCS06dLGwUs67WZgEfGC7qqXYKT4D5SPRavg9i2rVf0jYD6NytRwjtKAuEjNj6
HKrpzskuzHDJKnPZ3Z2KM3pSDMobelgk4yGd6gUb+qaqPeDu7gMTugOXd0VCygJHm+1m1ciN/9Eq
nODZKonMhXbdpiPYEDE+gKs8iojkk4E6o0Q2Hu6vG7P6Squ2ll3dXJ6sNYF0n4Wqg5eiDdTr+blO
iWk29MfiRkDG6pPEVYdGs0eql1b66OYun7n9IlajKjsH5wNy8xZIBZLVkZBylPIUGuYciyvkAs3s
RFTL5BykkqdAn7THxOJwJ9ifMlK8Pe3xcbhiBFjNv9dHHIPhuOCtCwH6HytgKA0aFxI1bZpfdTJR
DkrGL5ej6ThGqT9vrejoYz4ChSMaxy58YDQjVJjUrzV/TGkOzwI9Jx7H0o0fWiEYlJNz/xiqE/q+
5fYtPHqbHXzPZa+58IXI4UYHDiXXluvmdFxEU+ZLqGf4kpOUChMmuKvOcnFExYPCMmih8R6Kl/RH
72uSMBrdKNvkFfI71CYvJsjdMq806/h58HxZKOaE66qL/wTVFdZyBcutyf+0XogDLgdT49OdEpVo
rjaittAU5qYC/dR4qQ6tEBOtDnWdPrqSW5ufxzBdVt7TkhP2DjoyJtxhJ668SN8dc0+5fUdujqlx
0CQfYgaXTEoQq4bftRRVktcK1cZ3CuPRu1OM18FrY2Gh6UkHYvOle0kMs4yA8JAcCfnj8gpGdnFg
XfvJE02eXDG7qJXIPBh2ZnBJ6UXALnr4WeKwKcdsF+4xfbcH7IsTbSR4Q3CjT8eLX69/OagoY8vB
o5N5Ys58SR4jjntyYx+/q9BztpqQV5W8wUCNbrlQ3gtuZFfupAheQU3jICHPqxKfeDPh2Iohl9Fi
N2oc2RRR1c7dz3xyyAj8szj1zt790pVL9AAVikWXkbcstoDqnK5B5YvaNQuBJ/oN7yvLiouSC778
l16trnyb5aN9HDFFRCJx3fnx0WYB1T/kV5Sa8h4dN9oCZwswcVVrAKeVoXhmIqM46YfggI7z4Czu
X8CAjqcY4gXSNfMlV6paXYBtwz7+/d1VbeMAvOM+zlZ/q0Nme/en6Hx4Zxx4u0JHav2mJjZl912H
N/to7VvOL7WB4YAOQZ5Syx4KpUYqLQpU5M+vKVSEu6DW7TaucRxH8AMcEtBQ0nAYyd/uuMISPTZU
zsDjXFf7+WQefdWMmClVi5eAJKvPwdgwgDIrelbtAffocW50XNfxT0A2dAHN9K0uj2FXet2RScqU
/qd4Plr5HLR9u4X8Bm2ugdXdD+qB3c2VSvdu9dy/XYz03YdoXUP05a32sKo9H2nyW31jRqbtKpta
X7px3Py6CFZJruGSpA9nhQJYfKYT1VFJ3xuOiDFZ09gW5YsgVK5bNb5Ii+0ib02llwzeUmKXfd/L
KLIe79xRswyfXaisxpT4SGQtp1qJ4iPM2GXp5grm/jldh73MyjIy3TH8QZNhZPUtiPE4UM+5U1H5
NqQKibrAScPtv2XryGYldroSuyx/x2MpvsnIF/JUpcLIXXZaxWwRGH9elKz/8NL4Ly4Nic5Vjnga
fzgmjHWoESMkL6CodKrVrvpX1IqP3RZHr4E+FrSMs6VvKSOKXja0+BNsJ+S27No130jKruJqDHNo
heN0bjjK/fBkjGh8bDWJnJwykV6feGAtzuqXNFxtrhehqudX+uWC1+5bevdtDHb9bk+M6iDc3Cg8
rnAPYyw3IEfcyepRloS8kdThix3ukUGNIzW+pLCEw79rNn360O8C07vY817R7/cTbnObSGVPYeoL
AvshcnhcHwbHN5BQ5sJnqnYuhGPXhC//s7i5v97u35+Hq+FHJP2bEc5TLEdPzF52NN6vQ+21ytpo
3qbb0Y6fap0RfhY7SWA9gAEC7nK3de7DY+F+9RxW2MS3n9KRG6EsFQOKl8dsuRxB6qGEBgp5FANU
p2OsbMIfoiHhZixvvqIeDL0K7WLbaE99T5rHZ17ou4I+2mWHyKs4KAcXXDLXv4lEV073SuzqTOTE
q3ie9uXo+f9itap9xgoch+5X3jFdeZQ5Q5GYoY4QclFs+JPhv2B2PhdGMDq7Fulu7HA5fjeGJ/7I
WqFru98XkgcCzcZTX+jwZ0GJLz3mgVB2NBLcbGG66jf7lGSwkhg4YQC9G1RTc1MLJmRy00Xm7YRU
7xVdWvtlDmGgj/BHLONYh+6m3B0Tj+o6qbYkkSMbWE5n1AWwWEaUMXcIDpREzidAXyMnD4RNgz8n
LKZqnCgSGMT+r+kdU9OVfTP8W/lxhckB8J4GV76G+/HHt++QCEsHOY+RL/RP63pepYjX3hm52RUD
YkGmcVYxF1nv+BSKNnndhZPNPF9bW/2BeQej1INXZjVbcTdSURO7zD/YNCMkGy8YmW0PMHpvFg/G
JLjoiqE2KCpvJsee5G7CVfmKhAuCgkAcbVaKJ+KowJ+ZSpf0qoo5nh03P0WAWd4ZJMf6T82HqHEq
Or6N+xAu9w9mjn0hdMqMxhzciDJg6psc4MgcpmbS7bJCwTR978o+S6ZLJ9qtFJCiekvGeUBM9n2F
On7WVkPGanzqNXl9FwTZIA3VyUMO+W/wOQ4kZ0JJajm1k0H59g80I0OwnJ+wYQWAzNOlr5qAWzfF
EiaJXw5tnQqSnHAdEe3sFgMAGp3O700CWaJUkeO87kY0LbAJQHZNAhRcUbAA3D7fISX7DIOh9VCH
wAsDssqwbJgsFBtVAOe35JmHzDMoOyVfSakf3uzXB0JZJB9PI+PJrJWxCvWYLvBWzrkheYU0p3Fr
/ryhSZFjSF5GHFFlvYJgPHD0EULYdVFLBD9IiIhc6ehMuNPWkCpstBMP//rbsi3mnXaBH6fVddD7
KGyOWmae9KwjUxApcnzc6JJ0QMYzQXfXsbplD2z0SjLv48UalDd5btPYGIZJJRApGeujIUGci501
+u7EY0+MeK9qlL06YsSWk9PavqPkUyzAGUl17su+dW3pmbu8W6GFUwyoYkLyn467RqwWPtJvcGMO
i+II5AZbpZUXsFMqXnAsFOh/IX7EBoMtZLarMtsABl0KoBdEMVWoTyUEAyT3N+Nzuu/tJw78126K
FS1XkTDr/VjzxxIqgILfA7/TFH7V5Jr8bNRl8IvkvbS8MRmHBE8GTk9WG8AenygUHA8YKpzD1lHT
nE342iOmKgF2w9wJ2Edl/cSjAIRFLGFfp5nW/64r0adxzhvxKbp/PSCtyDixWOCeoNH/CwX2sI+M
FyKdOProVf4b8PeIvbc8KNjsWvuE9y2kYV6b0gEbKESXi+EVN0daMNIIzaEqN0gUxelpqKPyQWCN
bX6uw0sFdfcjxmNYUsFmmEQ5kCyFJVZWM8N1G44PaYA+T1DbkPxoz28ei+k8tA9ZEzxO6ybpYlnk
/jEuDMsKfumyS5EI1cDX+iI4apvIEzfw+huco+R435EnEUfK6eocCTY/HKvwAn3ZMaoi3CR2b/wM
QRG55fIXNQWHpLDZ+NAdS+U1Pt/ALk4xuWkk8X2LrrKnefiZkGhU9QddE+ZRqILii8lxj3owV1B4
UGAon8ElcDhtc1MneZjdkBEWlKodI797YRFM93Y/IvZdGZatQ5oEIL366vuz4fy9eEJIRLfsEnDX
9xBp5yBFt4+Qyg0HX9QzmDWzbObg+WhpikKfUeRtr8wTmdLzwkLBF6nqEUqPYmSFMrR/41eZkNVs
OiXZE6Mh9zPE9HnfcQrRtV95R85pbaQjXgrjnnLqpTxuv/3WnIWqRxF/5u/G3zcNCjn2xWjtT8cm
gGtQxQSTgiEn/mOyWH69Z+5PxhmTYCrB/bRwXW0eaGOTdJta7Q9JEDk0eYryelFg/cAwWQTCkomz
8ATKTKA1dpGZqMwXIDVBpN8gIaYa4oar5hb4MtDZgVAErBqCZl/USUoY1RazBUk1qPyCbNuSPNTV
7GMvJoZm/3blFZAxEtl4WB6zvm55euhk4hJl/2LekCM8shZzmzYrVwIC0nToIC3mZ1qR5LjsstlG
hJHnNgq4L7R3vA7Q1RAhWYcOvVJd/ORQs56QSU0i+kaH/YZMJXFMtfCeYKSnbvhunwLFzsXNge2d
mtbHWF0QUCUTcCkai0cjYQJoPVxuay+nnaOoz7JZjDCflBBlpVo9v8A/98tgYVY7dIb+xEh3cKBV
GkHDPb+f+5I5fxTEOBUFBAkUckmmpWrBswNkkmXjq5bOO2AyDWCOLiRgWX5ANMUGwivzR71Q/7xR
ohw0v3yB3Jy6CUAP8tseixXXvSozubO2vSmIsj0iFDFojSa8O3huCXuMFaZ5KxBNWMCb3NZ8kvOP
tiIRfkI313/YEUrzMGSEr3Az3wdWoHSHllegLgHe7RxAAEOmUOevafrteQ4qOZGyB97yd/J++RrK
mlz//Rftlw0W4nbCuHE3GSOxqlA7F2rt+ZxpTEBBGnKz3qMYKSB6gbs5sicXhm7GlSMI++rB6ZPY
PljtESjhJEOipRxJt5AA5JHm7qZ7/vvruhlpCdXgs6mk+5obpLYLWjHwlVEs2YAHAhCW7uYxiJCq
SAHEM5n7vdsABMIJpYJGYtvP5kqrX/lS72PSyvvx6iouv717XzbrxhYombg1DjrIBgVEuJ1gXdEc
B5vQ6I7uG4q2arDwWMiUwZK4iunE9FCdo34BPeoxeWlAM8JDodifTHcNOmA+9jnlPQRFEeif8rHj
Y6oUWSKBmQ8T0R4Mfz9y4uneh9azpE8Gy33V87397Sed/02eAY0qHVV7vzdA835ktE/L1mIdDGi4
U8xvk1cKBIxt80LS5a+CVhADaWgkTuyU+mEmFrORxUFVjKYMfxCutVc8VglkuzV7kwLXGjrSSO9Y
6/usBFHK/qDc9ArE/xdW9F/sGhE7Ro59QyxrkxjrBM6cepn2BI41Kj/QtJpa6Y2s8F1pjBeuX83a
lQHnmG0/StYT0yUkjq6mMH5tMFXZ76/P0AwHyK1JjWhb0GCDTaJld8Z2Q2QaviU8j0glxSQ2wm3z
ORRPXRt5IcZeebMhiRWruo5rFtAqLBVbr5wcsy3pzZmQN7vx0y2RMJ73pOcmO0E4ykN1XEHf4VNN
O6C1Nxiux2HcGqSbdrf95NfQu7dgeZf2RBet5vYYLvz2+kJK5liAVra6twRudNSQQynO8VH6XpRf
S2RDYIjFvGG+56n3pCoAb8RJEU8ZGeTziCwE3lj9GuSHySAdjBOQYAZmYSZ7Vv4vxkeKDSO+A+5r
aVUtX+bECLR/2QlyQYhFc/+ZcQWuU/xaM0LhpqIrG2ac20DsH9rPLJm130KM9smfkULvClzz64cI
SHgWo+1egPqs/Ov6MGCkwBYeVUp2h3x4mDLp481HTqAy0IuZwO7iQEI9FiK2u2FZTgB0qttKrX5p
C3q+9G1wODb3GVtzmoxGzuTj7MHrasuQ2KHyZ9ZT5YbNfSCLdY9q9CyD7QEby4Zfy1WB/e5+gyca
kQGKOK2P9qY8kDleDCePayDh6PQOtOg4rjw3H9TIPIsCfQ4r+XxK/to1P3cCeDeZLuqIF6X8vU1s
Q5q9ZwCQITwO3vbD2jeO9kYX/T+utxK1si7qVDj++3fXoEZoiSxHuqLGJf5imU6k29ZHYGhZCzjQ
9DGIH4FcBfBZrfPvDugHmagI7nNdB15Be/OjSsB3CH6i5B5Nff5ceaZ6Jw+yjlkYBeV28wKBy1g4
pvUzdiuQqxXBy/QkgFuV3vIYpgfWPAXFe2fPwhjdZNqbcP6xJJE1xD+dv0j6dt3X3FaVg64LRc2U
ZfNz6nD9jYeGN6Ug7j0mMIIw83Mnw4nob1uwrXFkKOwCLHlA08cj2HYK5ectIA3MsnXAFwzGvALg
qMIs7YaaIGuzd6Q67FNKpMToUbnWNTToxYF/KdHPnjgM97kyDu7VYSyDfBDY4+Qcl02t0ZZ9uBDu
koRe3CJC/Br5MalmXEm0/aW19GYfVM5lLBegUjKsoblrVupQkhdI9TcQPAkyXrUCzyEhyOOWTakD
Z8TtTRVzQylgvtzBzWa7tQIhmCxf7OqC7TnuLJBDpoDZKzts+IQFN5FjvO9bryGDAkby/U/DNBjA
51vcFYOUqfxUP8wjHODU2bvs7igd4njExNPbt0l/0+6FDN1tVb5/+p1VaJ6MeKkeuk5orqa42io0
DfDxxOi42hS8uHfq6Ho0l76AD10vi3LzTvKA9NlIW3k7ZkfGV/GyYgN3ue9fbCgF8lRDohOSWgro
XKp0c33NqV3QYYZDsSyMvCziWtFC5aADJbA8N8dLalqySjzBaqDolI/otan13iO9PMKYTeSO2yh9
SgJNMlUhUs6DjNDJds3VcdMBo1k5EcFcMt0rwTwUcw5wX5bIWztmLxM/coc1631/aNdNxrFTQdIn
I3n8eNm3r2k5jcswPeFp4PcGhzMEYpDAJ9UBMxrCy8j/lmx94JkBi2v2cMScxvVdLjImL86SKIX9
xuOLj2m+gtVlKgF++sx3mieGkL++2wQVzwXyDfNrP0C07AQHYtJANYAMrRQb+lQjbwUq5bF/Ajb7
3MG3Z24oJ/+SDyy+zvbcyyNi2Bt6S9GpyyklBcScONrVCBPQaks+lMM2Lsj1lhCFUzK6raI2t+2q
B+6yjgw0YNfz9+JLpj3qtQdrnZ2Jn9dOjYY5fpO61eWpfT8xSdgV7S/uFpcqXUKBF+qqNLLobyhE
OA6U/NNvNXNmIHRu4JlXOowJWWyapfY5bXBDLsy88pzR88+q21kAp++iLFcsdpacSPV/NY0kDnjJ
5VHYGqmoiufoIqbZzXk78SHqRItLckJRrJMLNQN8w019LevDL1IU/WMQuHU7/DP3AJPlVICpof7d
DAkQbUKY+2v/YbMb9a3Q7m676gv0Ssw647mmoEZH8iShPvEZNdzmoNYMIH9ityL3T0ExSIvH9Guj
eK0Rh4iHwjHhvaXbBlMQNxULWx8TSbvEDHUTlvLpQvsTRQmV2dWJOj5RgvqsyttUYAx9toG18CVg
kV2ulFrHZfSwnfkUapzkrxnHxkhiGgxs8FyoHfXykKQPkGRxYWvuEUsr84DBnA4LeI3TMKDsbYxm
+RQR+gnXngDJwikoebn5rK7cfxHixFpnvdNoue2Wf2wXMnfJ5Ydxpp5d8O086dB3f5fl59bZ1H14
TJpyMngkHPxvMELpJTKmeIerlJxlXdSDrAQNK3+9uSk+xp/ybtJIndgad8ZzV8K+mlICHkrHpe0B
p5PMo5BGxfaOhVQLcu3yzYc7CZ8m90dkRVp+9cQ9x0WJTTcz9wtYkY71oVE61/+I9yyPLJi0mnPA
0vP0/cJO5PMLhGWFND+mN0Z01s8FCTT239u9zluZjxNx0tVxWvnjLxzw4HdkGoihsj5LIvYV5YDx
oxQ6gCzwTQHHmsi53xQK40rE+UqsUX/aBsloBYT8pUX+nTqGSMdH9X5qZlFLTl67XxRPoW+mvleh
CbIw0HMSayP/2CA8SvZoWnQJZrj391nxhdLbXNoE7qHf5dz4rc6+fChWTS+V7hEYw7ygd4MPvtJm
0d1Wc7sfenk3zkg6idM/kkVfbEqLR1CFNZR+jI8KuubK5rCTYzZwrnqWE5M2qYP/0mH4i3E1fEH1
6xFEKchgiWKeKg0EG5g9tGznXtpT1bm2IzDqLT5Y+7q8FUQUao501tecyQ9sfuEqY4xTBkzipG/j
Yfn0cvXvzOHubHEr0mzMSJuv4AToPMl2+FwFS25BuyBIcYC8sJjxLTc6T0BzBkRpkmqseiUmcpdE
mZPpbi1YDhmgcGMAOBRLlwS2I4Z/MZA9A0xRxpvReeqf7gEI3pvUUSTfebhP+fnq+cLq/Cbepo9T
0ODGsMRmM0ChD1OANOpkIXzdj21hKT0c11HhPDlucz4F7PNNL+dYKz6/mdUdsA9xKgxUN7xCDv6k
mJFIu7Zc/Q4F7x3lnpH5IU/pF5RN4RXazCxHhRBcqTD2d1jXHACatk1EZ+zOx8HzBp5xbCWxLxX3
2k0vLN4vRhMBaCFYetOlB496TppjSK4/D2L4MIXXN0KyfUksbgiF+cLVReh6LThUhKuFfXlwTWHg
+y3eqiIYlrjHnpmP3Efy73diM+bSyyvJimmf8B1Lt5fSMnzuUy3xl7z20LB84K3OvL6CeNAX1rXX
ADeCMPvg+Mcdz63065S1CCVk/hg7t2A1yoYbzP6svwu9c932BohOw0oGPAyjlDoUOuAUtQJdVps+
7QG7DCQ5dnxnyn0Rdblpe8P5OAGW76b5M58sEGrkx6XPSHkP8tySpAVPrWBxAQoLGfKLyV5Y2QWv
duwDBhpLCcBqlpJm2n0/WZVSxpktnyAMcQxz8R0Y1uZ0bZQKNzhk4CNL3BQEU0kJgjY1ZSINAXt7
pTa43OVmrq+7OVGHeYNCPxrEUMQydWG3T7lH+NAxe6loRXrXXl2CFnuQ463BL2nYZ16TyAbbOSCE
TChCO20jCo1a0RtQ8Yx8fQ14PL7wxS5NmJDWRypRrz/jxJ39piDy0L1lz9xyPuFn/pDNp8zeCJ4j
atcyaEseg0AdthcuLWy9NvL+e43BAu6NBfg/EPCshsg5WXC/KvW8f9Tn+G6x+ZTcb4HklpRFvE+r
gOQ0bQi+N3YVCCRCKQVLGwhOvuT3M3vu4RkEhSPOl92NQLRRTJl0F7cOiD5fdP5VVpUUJmtiQymR
04EaU1tzdjbzcz9GmAAusfbZvfMjwIWXYLRtbSVFNvta3Qj3uD4/jRjbN6GRecJ5GDlqQ6wUjJ92
kOMD1PX9QvzsYT3Uiryqn/Tp7s16tWfnZKAV74O/oXXXhmYyU6pf6Ml1L/7DhqRQgwoy9HhKe6HU
vTfI2JDlTvi1nct8CI4ne+t5rKLVcm/fSW+q2IKXeN5HQGj5MUPcu8o5B+WAZUxNL/grgcxbidVN
P2GlzMFNFJKSkjzl4N+40qUtVoODWYS8FPKqFpAvI2xQqRs3QcLApOujbM62j/5mMPmTfK4Jqbn/
WXbWcuoYrVq5eTm2yCb6YmLF32S4DfnMdQaIYqbF7c14UYEFMDRMrvOTZg1vWhpSYr88Gr4NCLwi
VWrTtrz1PZlLz9y03q5NrXCSKK3lqU9iCvzD8mbR+3JCSqpqX/q9pK6pxtoSnTjlXrt0CK6bc/9Q
LsNQFlHC11NqFzeqIfL3pdXrVkMWR2hGPOZFwzkivgJP/X6AeuKQ4sOXGPTG8ycmQt7JJ+fBvfbD
4egtks2OOf/DHOBcilvwU/XPPvgNNftlToiLMwZ3r8DKc7mHjDzG5Tspup1I1/Z8VTBdIqGAyFVJ
xvNMYzF90VQV3yrm7CiSmmReVpmjuHTWrSVvXbl35lPN0YYZmNCgpgD0laXljKvNM7YuT3GFsJ9+
roto0BRIYsnWQ31wKd4Jvste2XF1fw3I7cl0/smqUfNTivmGyadlQn+0NTG8E0HzHm/yEeOo4NJQ
1qitHlyYxK09JjB8VTR22ovJMhviCbLmZdLWVlTla7+Hltq9XSzLUTyZkDrhrahkJmBZvPvRMpU/
LCNejA6LiuHjno1GTgD3TjTt253GB77gdOTTSRNkXW3IpuleZOaw9bRw0EBeVqYrrgrpnvqCb18k
P52qYAbfH8x9Xa5Ur3gZlMejN303TFCeuSA/sJYPjKFtPsEF1r0Pj6heswPnxGIJwRecJNz0hsct
8MZICW8GvqDRFtdHsjbS69n0KfXzrS97o1qRqvLnZSTAnMTAmNgt4DffJSKaBqMcxxDA7ViP2Zcn
TKVoktQbv3EVV+k3t7obLCaHjTho0rM2cc+yTqtUhyJQZqEQtttDEUI+4KBdjIgWcgmOhJfQfb+I
kC1MvlyUZUsaYv4Fnn56lEONBeL7dKXWnVbtAFvSlWvZIq8upm72uo3zbRfn+JqeVGQq/qEzZwo+
6jRhIKsUbJLELElo4NvAZ5KJt1h3LW0Pc1Srg5gbXTd4sCnUtDsh6p0IMEOptuVpyOcp+aT24CNC
sd9lA+AWa1MR2zeWLGeXY11lR+tgiNkTpWRgn5qVYBZkr4rZCKzNyv3bFadRZR4TyZ6z6YQKOu5D
FlHCC6eIG7MQpubZ6TXPmg+YtF3xLc1quWj+wgu8u/ciovCfs4Zms5w6gwW9eE/nv8YM6iHvwaoT
eUuxW4WbnkTK/cLbEyW58vwUDJuXAOQCqu+ae++JMS8Xbc/RZMfl5VNfhs3mKuY91kedsrIk1Gaf
BdvEtnP64yiwkgzYShHjgC9F5rfVrf3E56AAKe7/iqEYuKhQLg1NlOlIHsQNOaEBMOCEJJahfvAc
9b1S/2Qq9gHVU28+E8nkWlIqWUuQtMfeMxC7p2T3tVgK9Rk8lLb47YxFzI/L6Bl3/Cm4IgzQ0IfD
AO6urIbt2+BFyPTRryFbpnZxcwnIU71l5TswIdQs41DzrraJ4sjHmkMkNm8crzMRC2mSI2cS3loi
eZiAsrKWUzokMzN5Verz93PP/0eMjxLnr87U949m983f92XwSVFC1b6+gjJQt1PsJoB2yQuiVphJ
N2jlfIPNA78uv8TfKp8AiTlzxYYIgOgIroyJe3YLN7dzLURhGh5jOG/8MigePKW9Z9pfeRaKpnBP
mU+6G/vceVOj3nxO7GZHoPki7AkHfrMN1jwmytEjO3jVP9UdYX8uPaQo36amwy5P5LiNVEvQJyFS
W57L+AEWQ/ym0GSwSl0B9aXRPu0qVhBfAQpEyPa5WoDqqUNlw/6WIqaJNI1ipszRvkbKeOzFR35r
m8sUm/hkBfhRcbw27lALyR6RScqveqsJCSt6ho/HDsB4Dn2gqWgKvdpQv/ArZj1qWCQrdTjlMoC9
bzfppk83jXwLLCZajGENTkQOLnUPiSsAEilN31/yDmH2+MCvdwRg7ofwqPIhuH1j8W2Efby5uVi8
Eb1RvIOjYuhDR1HtxFZ0OwKKds1IhEuLTB0T6H1JuOMfiaDCPDh3F08ozsjm27uZvLi6bSPc1KZ4
9WGBWYdZ321O7W3zw/XmvwZF8gsHd44R37TajNeMDy2etaSC/ycaf0LqY4Ps0dbtIyvBopW7Ios0
VOjmBAFsMydb25W0X2omjn9YMpPSlOB/IKrE7eJUpzucMScm7S9meM4BPt7YIrUD+Ypfhy3vvY0S
NpbmaN+dxwOe+w+JMPQOmKYvwYyCTAQMC5AeRVPYt0lnXEU2SQqXu2FPHRqS10Ycwk4L3BaY5HQW
0B32BMSOl2L0c4HElB5iZPtcu7M2hVIN85yMpA4BECedmWBFM5uNTmzF+0vYnw/QJ3WB1qpa253k
b7JdrYN81FGFPCO7ky//yuVAmRqZudQDUFse39Aq5Mx07npn49+2n3ZSEnqv+TrWdIb2900YIIeA
gKgy2MLhNCpIzDYIbqqLTANeBvOS/8OeIZsEJM+t0A1hnH6LAscY8ki2lnEMDutlG7gh5xi3Syu0
tRHVbG9KVEy4owh49ZIfS+4Pee6NLPRA9Ki2gFrMEug8hhsfluCp2PUAgHJRoTgEU6jJ73xvKne/
keAJ99wSbPL4EZoeAQ6BWAi7CjGGSRUSiqd//bELoB072Nu+q75/c/2TYpT8oe2wAV7554X1+9y0
hOKu19ipDkaaQGyy92QSAOA7pL+xqzEaOFy3lTlSiDh3hO/7nNXw5hB9lvAihWrtHezQ3L0XR2tr
oY7II84V+cBvi8OO17yN71VZvJYrSz+KwqzzvoIeoH6aIOmIbPNn1nOulPolSD6L099k5qnEQP9Y
hhXawdYOApOpTWjX7a+UHKbqGKhemz3HL5vbYNJA3WGtgk+cwOI0NYNHCxpscjl0jUrV8R/hOSFd
xwSx1aY2B+wyTkPlz3dp5t7J1CZe16KR7KCZREtemKxtPNap7PVTqT4gzYgzAiePCvuQiycTzAd/
AhmHM3+3leIaxJWjSfCZqv+dnfHCMYpr+lqR1jXuLIUBWKv/uF3d4F16wdx8S652T1+J7hZxZ54o
L/FaMKkSLy6mmRq++dey/pg8svil+LZXYxZO0+Xh34oMcTGWyiMSKJ67r2y9W4Lbwk2aof1Qyw3T
X/WIygeb6upQsdALlw5iBwkPsuHFooX0qVyMCVoD1JJmct26BM3agcPC5C7TVYBOdOlJ7ow59ymo
afP8LWz8Mi3x6XAdgAP+BJHoLINoVo2qyIsLt61hTWWChcyLrQCqdZulymGMtdS5dAmIy5KpVCzk
rAhJoDGUZUux9Dtt3eI2/tQmUop5Ap271Yd9qSDrnE98lUb6bAPNoSmWJy1sKpYpN+7FwzJ9YNTN
CKTfs0+vdYtdgVkoXtuT0BPQi/12oc/kPsymZtBA7TkUMQnHHlvbGftaIc7OElPBN2QofIu2Vy+8
nTzrvql3BBF9EjS4NiK9PRwBBTTXB1Jk4QbCMDBDBQ+wgfxtQsUdK30sqKHJadsqMmAAhUWyv/0E
p0rpwcqbpypORCVcsqyArr/yvmea8m7rn8G5x2Tg3ONFdHNlcHyq6KDXfasIr+V8oR/S7iJef2m2
cw2SqKLq51C7KqD+VAwE7jRA5fG5nJEizEFk7rmpaLbTbIz2b13qwvbHXuATGjF+kjtEieO7JVC/
3GgcN4Hn0OF4PBsYFZhWtk/VKnSs431Npp8QobH11AQdcn9d9Ma7tksnFcxVsBksNxEdJ91Hqbo9
OchZ04u2+LKFpRfxaB//A0o0fmvX4yv1TYKwyt9XEcFJ30yTI+8N9DA5LIf8nkPAC/dor+cgYZ+G
pyodfzM6v1P7mb3t9SXbiZWsHHM1N/G0JZ5k6csVztAiLBMGsJ+Y8VIXtrZdQzvIZhQggd3FmsMY
FtfAjfdq0tr4ra20ps7a+sNAsZEAFBpqY8xEWm49qHY9pjfBIqoYPmpQ3PZU2xlgHXi0mgiSYsk/
URdTusyczXq1uQyGUnkBN/sVQjHpXcrsNxqdYZM8ufzq4hqaV815MX/eeoV5PbP4RYSs93GXZGvb
OBWqhqOK6L92t9FlM+ySYBDBOd3GGQy3+4V6r2bFzYXtVlSS0KXUujIEz7mg/J416BX86NakxweI
w4xCzlO1G+dt05On9UjP27A6/5+NCnjcnM8dHLOO2k0wmbYFygs+2UQtxN3wn1gTbrJZK/SI1+vH
ACNIvjxV1Rk82ZI5Dt0SQa2XB4Eklzmo5xS21b0aaSvF8XS2CAO/PmzFo8FUacufimySMOtV1ZN2
c+kLJRYgsUfeNkBnBeJ1QIImSr6KEjCzEaZ3gM6ETq7K6EcZTYDFgdUQwe7x1BU4EvfMlWqyV6hG
An9C0qB2nBsfYGf/8uqJsKAbTBKmG5kmofKqGFyd8VqQ6iNx9BMiNen+e8bDynbrLX7UKk+gWwbw
5JGNZPlRuM75kljGVXgHuqFnkkNWyRSH0VRpDpO7MQMD+HDesfEGzRmoGhATj+o9WlZaOBUZglUD
CvqoMzAB1hlFuUpJoHFmXQPOPbRBYBMvcN213YNULxrIib/00oDCnsUWnjQurLn6CkOtUxqACRF5
F8ojvqEMuZaKRB5Oh1zhPXN12Y/yJ/RhZ8HfOL1m8zSIJNFeXBEgCKObeK0hH6Md5TkA1OUpQZAq
jbkJtdW8GUDs4C/Roe/yHEqyUcUCAA4+j38q9sbL5VM2V1A/zKJKzDbzmKWkGynuz7C2HjDbksLs
x6Fd6bJYLmn4U9VK/iJMsYz651OIBuMrXvOR0h5ZsMcb/vmojDEc6H0mwNyf076VIbSpMyn2q00/
iLyUwv1RJJfvdXc+zzIgO5svH4wrcYs8OAWrG1OHEi+dINIjbdff5ZH81Wy/ibSad/sn9ni4liBQ
8jRo5XgO9qy0u19sNwes2fFHjaYxEVHGr+2+f1w5y6aZSaTeDXfstYgn1X2LOjyAzj/huFaQ3cUA
pV8jWVFFFTIoTKkYvP6uvL5kDG77U2SIgyyvbC5x1BRj01qOqZ7TGI1omWvKbbgV4mFon/vQCbEg
VfBEyBIelXmEWVBXVXD2akYEiJAFyfWZyvtwC9RvJVzshVAQt5wPNZhIIQ+lKwR2leny5r/GYR3i
/sM9pnLDSl+kbo4HfW3p04vDsh+/HXMAvHSaH9RbOdvFmsk79dVvTDYS++W02VU4KUes4PwQkxeE
QE7hHRev1oVUrZM3hmJDKktKy5+5y2gLFK3+mKkkPXt7oXp8A8gFLFjudmwbsWvtf9wN4pAQm/Qt
w7z3l2JVobvw+zLFTbVtNFG2xVfckA1joLJ8KlYjlZ/mnkXlFGC0LmKea7Q9PJif/XZAUkJscDH6
guehuBMMhdjE6f2wPnjNMO1OnHpibL/72i6Y++fyJXyvbTN1TJ5wwQGEiddjXfkmM2/3iaoacIbL
QhsZE/t04D0qBuX7Vk+C6GDFU3DzR+eXv+HaTzIn/UzMfzgjXcp7x4xrpLakB5p9+/obxoFx4G4V
aoRtplOGSy7FuPh4Vww8hW1JnmDdsR+utwROKDnYSTbze2Y/GNaO/IsfEdbGy981dZORBs/zmry+
GTBp216yaHG7oZUpdB0CvvIDqfEIj43mXLsuCN30ulKVC5LupNNE5omSxCbRDhyO3/pyUUWBOPc+
qAfqX59of2XyFjrwOn3CiBLKbD50/iOlHSznJd6GmSJcapKYSQ2mXAVWcXt/y+S28OnoUqNk3HZq
b1rKS2UIbMsP7+4kr0ry4oBzZnFErCuq8KNqJOvkv38LO+ipXdGF8a6VdcwwE4HwUV1Q7KALTME9
hJRGjT9sojmVVieKyeJmp9HVdsVhb4hpKywBo+NTZKvwwPg77Gri4yvL1aX6wtgWr0dyDm8R+CQx
BU3oByWTb5uxLgPr+REu6yxIG5E/pb3WPlNONHSCpzZUQaW/16ytIyDTWc/2Hde3/8MUX7RMAghy
gVxQJ5QD5iKZ/yAyocpYRrFmkIl/zYkplB960wXABrPujIeeU7qgg8z00sRO2nDklxzx+FzsJk3i
Y0c1pV1FTM0u1Nd773hz6MbM+5SIHYrvuO8JTU9Xjz2BK6gAHlmdKO9tK89P6Htlxx9L7A9MsFty
OBFvf8nbcufCk6ZWoXXEtcw44PBrQpz6yrPPCDQ0KjMPWQGMG7kxTVgT+ayvQy36WVfiM6M2EZr0
KHePJqUzx7Of0SzljhMvwdYy2VWmTTUqnd8kkM25NnCMgD6WLskt9ei8lv4h0ST7jo5m8AIFk6Fl
DEFPLEwq4s5X6xeQO3e6c2ZXARBoSFN/3ks34k+k54ll2a7kDfItN1ViddcHR6ESbdN8I5V0ardx
lwHpWKy926genAjgyq6mB+jKimx5aGI7fZT6+huTzukSBQGUMmVXafcp/AS9rRvTIai3xkRxvDXy
axyPREtw4JMf/n9nrcfxU1B/K6MVNVu4/roEz0pNsYOAUfpVbrJVk8668X/5DBtWkKASF3zCX+bY
m2W7/8Oye34MWBSdbPBs42Fkj4uUXBm6xXB7hDzNfrjwn7lFlTPlsFsXDXj5Vl7/kbp8Qgeg4JoC
539ppWv/gBLQrPsVbZQsduJ99oCGUodbQIv/z8Sgmc94qZo5VtfDbLsbIutnN3dQD8642Ab9GstF
jKs9UpQj5wr1VrM0Mei2JwN4hkt40SNx4eNWZxRAtK1Gs+eEVqi/90iguBctjYAiqoHp/kabOj8Z
Og+uaxSjotNrQ0MKP/yxDOdvD0nmrvhVPL1mBwu02KkQ2rXOZ7POpcDoXxnz4WHeXOvk/3MtOsF7
MXIA/Hw7Baz8ga2opYsl9r0TK0lMgdBBLnwpK5Dn54EfHQsEls++9m2Q5Stlpd3Ls8/ga0DF7Pxt
gHp5MwJygFZ72UU4bgaPH6fpIbtr1FIPAJYo/L1KlWmkqYae+AyeDG2xTn4NafaDXJKpy80gwfzH
nlUbXxq4dM3SrHq+BJkKg+n8V5tMScI1I6lCgbUgylYIxMVjZiNMf+4dkjzkLSIy07waf+PZ3ybB
m2MUdaF39f/2MJ3yn9JeaL3e1JAdDh77CL1SG3CgR9kX8YNUdpfBeazmlZ0aJjgnA6AMmzayKabL
blYKYLsQvbg1v0x2U7I6GUzKlbr9udwjvpmc4je/G7hqg4+QyWuIV7F2YQUAnT4hx83UZ7pWm8Nz
tEqivkDngclpKZKMYFh46RLTqLOl1xb7BsrRwvgsHRfI5sAfig12JPGqeMVINBF4OzXcPDMATdCj
Eel8QzUnZemcOcOABt9G23DKDtkbQvLJLPruHr/mAm/RBJFbMwzktJFWKmhFTZyFaYi1zJKTyMmv
SGArKTg/az/MTGZlv0AhzCs59tS66RgExu5TH5q89QlAfhyI0ITkHBDDHkF8wGxzklCRPkzKshtB
3X+BBxDoa8Uh2e5SAOLbkfsnWf23cmOpfFjuTI8C0ZlF3WyDcG5R6Iug688Vnysc82Txp1y/Sbi/
tcQX7/idNwwBSLbbdOumD7U0uAQuaUHHyeEf0igxKgI7WjNcaSyNf0am0jDabyeYf0pBZrtzlwjV
VjqGf2O5a0jy5RxeNVzMNyXUi0ST0g7Cswa4VGphg8ey1Ija2pY2xmXscCT33V1KpdCzr8c2XKYV
3wSnvzQL/9RW0bYIYsKeBRZrmSeKuh2aS9fjw8DDV0c6Nxr2Q6m0STSaaHuQwWzPNL9NGHTpaz7C
HxsmvtQQJuZCtcJhWhc+K04LbHNZqifa8edKxX/lFVmsa8ctMxjx5HQiC+ymYAZVLzpb4mMz9I9p
mb5y1V6wLTHMjBdnIzCP6Zc/1+GCvIB/ojw5G3E11cnO6zQxbxj5aUOOalQLsjB4favTjF/YHb7W
MWjNpqhAqJLVc9zYAw8EMotK8ixaNEMq2svPjOziCuheK3CbrK/XPM2AaCMj5HneLZ/Rn8ZDpT5C
HGiQtZx+xhIYMNKoAHQqZvrN7X3Q46kfjKKIIt+Su9Js+bceilXO4DTpWKewNjgM0AyBky6kYHhN
6dbbGIMmeLLcdMGkmAm/GOk6E80f0FHOdGJJIIFHxAZ0wbfcPFATy1L89x47KRojUeObjLjZTDYS
3BeZrfH866cGvXB0E/0eG3JLIsi3+gP4xmQ1jIu7OhlfR0UTwG8Z5sIk6Q/7B6hFn7EDAulVeFEx
ds1saMByZOOlKuwQEjpmHz+Z/M0kPOItOG/CMAiIFFgK46NxCLhbWOrTCfMlBRN5UHQ90zLuHINb
ItC1VGc7zmN9hbbi6Wo90X2tevyLD27o+a8hUvmlRRHoTh1m2iFb5xslRO3fFFj6nqafOG8xP/vW
LcUvux/fyRMtyyqGLQybsWhWrEshqQDvSpnblCDsz566DdriuX/VY25Ks2GXixhgCjQfEy5P0tdJ
mgV22tVt0EFJmhyjn9zd4Rykutx0+zGzESjgzk0XGOXBoVugT5gw6Bl6qwMB97CK0AjlH025o8D3
0FQQqdUVyEaODXVd25aEMXIb9j4znqgXnLs6jFXb+AyJ14j7LiGoEJKnoHDgc4Ix1JyKcSd4b+WT
DzymWucq+Zf2Ijlo/cdHx0ykLv+e33q4bgGY/P7g1d1zFlZxif6QAAeuKB7M2vy99CoVobmyQI2O
KfHQ6NAmcRjHX874PDTDZglyFX4T5pwGsIuRIhHlM34s+k5+MHrirwPkIOE82myDHx/xzHMx7SjR
v0U0/weMs5XZfJfj4RNmR/Ha5Q3HhXb+MeXJ9UcUvLFtmXTMjda1rxXHTiLaOsd6584h4ql5OM36
n64fuqWkSIUvpjK+TFO4aY3VV1ko8V50jXxYQnQmcdnQIJ///ag0dc4HHtbOtsxRGaEUM+pYFkZb
DerhjA3q8I9dr1y13yRxWWpEYnFNPwVgZwyxhEaLi73if8Ev/pcL6jHr0gtNBBvSOXqxkr8uVXpD
fdIT3yjoFgV+b1lD3rjJA3qu/Vfl4RiBC6Gvt8SM2Skh+HERTtYtUxqRqt53sk0KYA5mRwc6c5W3
u26+zybHwpvPBpFAM14WGdGXM8aL+9R3nGuE+Gbw6Aw8dmbRLstSinf+t99F64UH8cVwsLzHJhTU
LMFZhlWKJw2ikcmWY4SkZ/4zbrEKTLu0yXCYTnWJLXa7THwfubexSt/dyCNOAibm8JrArU5/Lvz4
eMeBfQaOSV1EKbf0Z9XZy7ItdFbwFtd7xhFp/Kc3U5O5kDWzE1tMDdvzr89dfJKmepdJo5nWO37U
6XN4jzmlHxu9sOipAosOlAvfjYVehvIAAkZPh/XI7WDnk7xu+l1z7JgBxeOZVy8WnGqMOOwmh2T5
mTlDV4aLwv1qBb9WhYrJDKWRVbhD+10ZFPSAVXy/H8uXyKxbFKPAwuJ0J0P2ekfggN+P97HSddBA
r2ht3tAhNtFH8Cv6Oy3gmXcHTnYGlfk8Kw3+r/leVKxo+pKyhhhdA/onu47X0bRSVBDV3TWqttIU
yxdERW4CCXcU+piDl+YFNqdC4r1RcPWGX+XV9aghLIRToJmJOI4t1cMM4ip/BO0ELHmhMRv72Ncs
qywCtW2+70ZpM+cu21Wkvp3HxoZ1877l+Ffqy8Ii2DiKVuz8XzQ/nfi7ub6cXogAQIJrQwJ045Os
neTtNNiCCWJlF8WryRnEDlfssKvvMFz6Woh0f7KssXm5yH6RO5ryqDCEGpk6gO/v5vrxQTeGJm0l
lxG4jAAEqOMugKa4l+8QygaABap7LDHze2jiGuNIN5xsylUBzRjqDo69SORCF5IgucRwnuyWSOz+
v97ND3QhNamTJxhzZaWYZs47mw/UqFK4E6j+tWpftuf2uFAcLxGqrVUMvWgQ7fRkxNCXyIPGrVqN
gqzC99yz29d3MJ4152anmnqlFMvKNB73DBMbSWubMyxtZF9C45B/GtcTAqMC5sha2Qqrv2gOBtFb
h2hR93H3ZFSnFSxi2efmoS8PJhhecfgMQ3+s5aXmVK9LQ2OWO1re0lYMK7LfB2BIk3z9MKZXvnov
6fdxzKKmICeX2xGFS4nB/betNVObWnHnEBEwIeGcHHfl4ujN9GJ3m+yOkYTzaDigAy+EuDwUGYA5
KbeDjkz7z9SxLXLEyj7Dl8mjA0Rs0XUbc/5ejtkmRIXXya9Nto5M4nSyao1xvXEtYgr9/9rVw0uU
NXnjnMFJjmXALxeQkDBhz8/T8hVzGlo5iB/1cIoTWv/voV+WnvaCgyAQ/SbfpQ3b2yS32eltBdDP
STmXMJooteOFIHo0kRO93Dcz8QvmFO8LWoZmSxRWE7vpxGpE4lzTPI2eBUyFGG9YcsOEBHC1H61x
C3XmnfWwbIyWdyxTdDVE5RXqGLhFXGx7OXI6WLaBNzpjC/IIdja4zVKN2BrU9ss9hmTY4npq9dOK
aJC1FwkPG/Oebt5egjq5ol5gdP7Xnr0ipT0YRcoAJIMDvFnNwpNf7+EtAKCcPWYlBgpEIU+REMGe
j9HjnnMz+ejiA5ZRzdDMyT9RzwbRIR1q/pwcfhFLmcCGlNAaYTSwbVbJTGGyRu5FjgueUdXOYNYr
59GDE0W71p7SKvAkl2Weap+4MutVjgb2QL8KErP4KOtuuWAxShsOdipXl5+BqQgVlYxvRd53jgvm
6IMtXWMkJmXdUglvOprbXL809e77VV9Uw6pAjoTV9KT1qmkZb7fRAg8kA8b7y1BuGZJvsG9UeqRr
zESYauZ+L+6zV+ouz/t3gVoohz55+y54pxgKQpunwJFldj7YOxrPcwyNaE02c5DIIc+b47G2u7DH
r8tSPDwn7Jl60LtsHwtRzQynuUbHw8GXm54QJ8ZCNqjPACp+Guf2a5eNeYjNBIEfUiZqIrJZaWTy
tCk+TmXkrawvVYUDTIf4ilvxs4SJfqc3/yvndt3r5j1iQnxCAnMydfu3WEJYa0myDRoTmOwjkB1r
oZf5UmPiSdN37k7fc9xiTKzIy1j4HV9PwKxRhKlmljE3v0yobuCNzRaYQe9+5Bp4we1FxdHsKtuB
dzMp6wpxjoMZxXFLGG4ZyMSHEWFOXTF+O/9NPSgAsQvcBpek0FPnT66cQf0EAbgYjMeAdSf2E5J7
lWdZ2a27DVmiJNFvHlZzCNGsqCKm92TjQPrtsNiNivZls26G4C/OWtrnR5dB4IP5ZtwY6BOk9Qeo
H+VGgX6fNx75tsvg79eiXmxcCjEAroo55CNsTwcU9kAA/UJmGimYzrtLpgTJ+1i2+LiKQSk+07BV
SrbFxbv7mXELENou2V4fT97hP8JRiFlHBGmibdV6Ndt9TfXw8XysjeCXtDbZ6T2l8BNkWb/IfrZd
j/02Rmt4TYkr7ZoCqAxxjT53+tZxgNu07U/CPY2m9sAHOxxj34e5rB5X090c5tt3gohDOoN0e1u4
I9w5+nlFJmOAubSW5FWAuJ1wsjIvyhFNVuhC9O+uFZzu+UwFyE3pEqbDrtU6TJA+RzzLoeHytc2n
pLS5IB62aauMF4rJLhgN6EclX3BEPPJNuC+oHQWszjxD3Xt3MSr3YLK8MSy8w1jtBmAr+QPkPtsJ
dRm7Gy3r6t+7P0oNveyqilqZvbRz7vkjs0i//HesiueFggPdHQhQNXXyU8wGie2P4Nabw5HUpeSL
XUnj+2Se2+kA/LHBkUQjwK+PfK8RjbV64q93RvZWPAgCfOc6sVLdu1TXv3Vtmx6Y0JTmYOBBTjwt
lC3Gpvy6bTjCKt78MTXrIQ3sjLAFgnO2e4ty0UjZ60yxOxKJHwcGsu6oJcVfPf1Radgmc2IRfKgh
ZBoIZJuiTOMUCsh07dXToUALw7YkgEVdQgw1FE5FeUo9LxyWQmmHtY+d0VmVFUsyJIhaI7w75TQa
zsWN6Pv8peXzvR/Q2Gs1Qw4Cck8E4GP+27Mc7TaYEjNBoO+JjzSaRZ7/Fm2Mefw3wkNz7WKzGzf2
AGzELjWqA+JYXANyLx/bg/NLsjMQI/3rDSO2pPHxKFpAIqlp4Bbcnnr+tgqR8C9WQ8n5hLaocyhb
VRMYaYEFKvOp/EEuuSdVpK6lfINGCbOw/0EfAfYAlE+fql3Ld6pR1/xbdMtm68NZ/Es8e5gKalie
Y8D0Vw0Gv/yRZPKK8Wgzze3vELNOHh2QLZYgfCi+z/X49nx2Pm6UIBEZ8OnFYiihCn1/TcIx8pp2
0oyLnVosjzpKXYxPYh5L1+MhzWa/QVZ+CrceLb6GWodIdBLCVpS/6fPGojwOUwCBvYewSp9EDKvc
TqjdLD+o0MbyeClK/iEt8Dr2RPURTzPP62zmKlaouAsT9hjJ9fB1aMphPL/08YzZEuiC3wrxqoDO
NWHm0FZl76M5FAgaPfqHJ9+FpVCr6TXECcuHVTtIyQBFNLHHzmuqbFY5mqkVfeEJFJkkhpFXOT3p
6MBSwpjGvMTX/AiA2QSqyFge4hmr9kt0Tyf7pOOMeewXwg8gan9tTQSXbn4DdiLr4fab/1g8ewGK
9lPdlFB7Fz1msRRtv4yC059AUmf2pQN81UFU/5DSZ+0tjWNAS8V6eQUu8SQIQ+nTGbbU0zXXt77v
hL2O0bnyN0KXj8G/pxJJEQgnrR5a2s6FJqA/aFcwWFNz0ceE7wTSGIl8h+nVj+oeFNM+tMRWtB7j
ulRgTWPr/J2vM5DulmVItMtNMYN3C1IN8QzdVBWrJC3D5NCInFZjNtfyYrHKvBdh+nlK2KKsFAUT
ggm5+1iLfjkGR9Jwp6Ga1OaCEVDNaBrFf0FTSN6uDiHLQulM3zGN5ab0eYZPDI5m5JbUquTo7h8C
STNr0wpmu0gqbnELauWtIvjZipfVi2Xq5tT8q2pPWKqHQfEEu9ESXoMyU3jUC4WAA67KTieocA3v
57J/i/XEJfFDxlOversopwmunNITqerIwPB2jtb4yGaGT0J27U/ckKMhjX5YbnWn1JvlVbTP3WXM
skoS4BQOSCHt7FpmDOm5zn29qU9jbFhbORk1QPPBdGDcP1qCvF/KVBDan4KvjTxkSWdfWw3iaTK/
mdY3PuMgI2Lo17vx+XDwbI9kMzn25LEX6L9Kt/XMN1LjjrPHHgYT4ZIu4gl8+tRBuSYSj5CNeB5f
hn7uq1g7oK0F/CNkXpMTlTkxN+kZLkwhPwwWxpfxW4XZIBzV1gQI4Ar+MHovxZy/LwkYUsrjpx6A
umZ8qPU5JdaKUiekyligSTDOrnuRT84yNPbuciaufZPN3pTRVsUzO5xn8vm7DBLPKhZZw8rH6dH/
uPBLcJrGve0AARvKS0HizSDtod8w4I7PzNDKqEGTRaGCqFGnrLEiki2RQdbhY+1C9WN9l2edcD8N
5zxz3LtskxDF/vBZJUePpHvZewIT8mXDan419I0+RkJ9FWasJcYoy0TUq+ZHy+z3Uu8KHA6E+e3f
5/LnIfw6rOtQ0rUnzdHfSEDpU23XSaxvtjP7jEUclG+6+iZYQLJOvXMvJNQuQedYsIRXdNihg0ZH
jPDST/Esb2x2uIb9mHPSV4dKkzJSVggzCfnSclMDTAZFVLKdGSWgAz5mRobLa0560QZJQVqiBbSG
ZY97Ii7LMrVouVXaKYQHAxzrNFbZgBDNsThuyQqnb8OSXuiP+OhcbQR4x8I39WKz+vkOGfTLfky2
uQim5aFCzVKbhiybaKI+hcmxMeC2C02StzU131x135cU9ffx38ld0eW2PslE4ZiFMT/ZeM3S5e1p
AdE78KisX7Aujwis3ZvPV1IkifcoYo/oWEzXSfxfUbefZoufW4ssqI6p8Yw21Vm/v/08RSgz9mcu
UON+btB/DkWWlRphZVSLWWoFGftxWW9rocRhouhJncbNxgUs72r/to0Xl+C+S6YQEYREni29D8aL
CPvjzTMh+Yljp3OdwgRS6nBx3Y5mtjyKKlARgD7Zaz5A1DN48TTCmbvAGt83jVX4jcRaQHss+P1L
L+8jg5QKRIpkom2JzJr10x5GnkaArTTulh42eR4+xMcOpBE8W+J3f/RIzFZ8b1OKZa9J+3qHoJMt
3PXNKYKxlPfUOull/v+vv9cMj9ZPad7muFuB/e2hf3lmCds68j4Tj9Ha1PEeB2fI/CtMGbLSfz6Q
E3bv1iqzXjaQXWZejiQuHB3HZlHeOcEWMHH0907PQJN5dYPnGB/ud7oPDZbDBzYiaXS/SBwCPvV4
HCtkK+lJ1C+oq/oab4SxM9QADg257v2UhJq/J6oQG3z4vHMxXRTHLUGF8hgsDfsQmxwDZkzPo7T6
TJAWNjSkXBkN16uwVfvzIhSG4zwU/KNfBuZEI9SDJl179dqtWAY5lY7rhDpuziZEb7RcXHc1sSZM
eJs8q00x18eoTQNFuTLz2mAkZ+xm3URAqXX81vo7UNQgisLuCL1ypv5mBVa8/kNyfRgnCXbt/lWY
ZiP7MvEbZiYR8m1mVEXrBpWb2bno/OixkHMI8a6/7X43SYH89359naJqLSIsCuvEunHM8QnfUtCA
k53AHxneLFJJHMAsmLDnycOaPFj4GX7xQLEJ5p0O9+TDfL6jkkZO8MW2VEUCdB2+eGirSLmcNMBn
eddXyKRObcrxKDBGetj+l1RUCV/FDTNjFfS6nc32NuE+d92vAztVpLAx/4Hp0Io2r7QA9h+Jcj4L
9k2QyjtbXrLlK7Rn8zkNFVyfw7majFZQATh/eB2XMUCLAIDKlfqLGXjs/Zrus63j5vSfyBucvKqK
rKUT4eYvoXyzeh3mV3bSflkcFtNbqd6rIjeiATbM7ysQd4oEZLJiyqyo+6dTKRRknrJHzsmN8AZk
6VTV7LkjEl4L9l8TqnSPwCubaHCFv32tx0sqyYaJeWTcxG69DD2K5shn5Plo7JVS4ANi/+N5fH46
NjPBGqPtJkFX1NfHc4awCldhq9AAPpi3nFk2tlrrfBz/48xK2kcJaspjJYeVjgdWm6ilTj5yFLVa
Ypk74QRh6L5V3rCdBn3nhEKQ209/ECLtwPIrYAjbRccfr7n8memRrgYCDXzJ85x1GQemwCl+RsK3
MBOaqqgZCLCVYFuNScAiRaOOd9CIMmrrSoBdcv7H/N4IfGoT0Uoq+ml5bcCXh5wxbeGxCFgfwCoL
kTRH8QwuBbOo/Z0W6T6+ryMOVItOLkt531GH2HAlPh8MwOa0ZsZQqoyOgquK+h0ajUexSenvp2bG
9wIfOlGaZmkoqyIWY/JdnIU2msk/Rb9ylzpcGN0Odu75AEacIVZ28D4atQWY86nTMwsk490W45Uy
8z0tPTAxKPuVFyewZZk7e1RaapzyTFTFlVdRQ7wFU+RSUiSPw/qUho1/O/jWVuFR02mIGdtmzWMH
C4NsWO5NPO1fOSOt7zZxekpE5sgviLBJK8pr3PK2GMmmYBn1dajSh1Tc3rEzb6VRinNfwRmX9jLQ
AFL2nDIr7+f+qHsjLkACA1XsyWRb3RaOk5B4VEI7CUXm2EliMk15AEEnD9JRoAncujbXFDU1bnkD
R1dQZmHItQGdLLeUPAahYWE6OdXhIjC+nZVwCoaa28Ff+7bwtpOP/CJcUycSIRgUTaf3WuB/hnXW
eRClOqIb7h6pyCtbQqFrRZ8OXU0OR56Lurm9iGqbQN3PD0eq8r6LINYhCpidz2422g3A+SB0e8YP
v+LQeg9DZpDSZbT850Yt+8hpqLGSpaZwDIsNU29aabl3cj9bU6jO8kgaAUhdohDAkljHAIbbM8lx
2qg4NWL07Ytx6Jxipb5SNLlpK58k69gOMa3mdSClTyNAPrLt6I/ow/gAbhNbW3jk/drxLByRNz9V
PVkAV/vA2FSGgqUfL8W+6oBCHDUHnY9Z6zkFfFC7GIksHQKdOkTwkkV4Q4nd/cLbc+kHAVuVWJFx
GAl8u5lLHV09QzZyMXsC+N20LarYxgLrUsGvEHE8k3wDiYhx9fBmfic5GC/UlqXzf/4/f1DGH7ov
O6rb64dl2TepWedAk1Ao0ZZ1hb6NKAXetbwwiOgQ9LoVMpt+HXdBophZBkvLPX56bNKsDcNSaWdK
qM6Q0ML9ANBYdia/KszUjcDkRh6Sfex95Nx9WimnGCDwSmVKYZa+8MCg4gF5czgE768d8YuVEZyJ
KaZLyXetnDdmNIyZtqqdh7o5AguMkbpTUEAazrMoB5FE8hj6IlV9CBaA1TVoElsJZo5ylxGghZ0K
2j0W9HlTfX4KxfOxwmhvgD0poMXIfM33vhUjmtimM7VVriPfBmqRG5JQHEjZv03n8fGfU6Fo/yl3
zr8IezMrLldloGWpt8ICBuey7BDWl6F84f+XroalT102yFRTqc60k7bv/rv9fOdOMfhaU7LUE3H4
fsUGMoEgO3Duqwu4fEz9Z7VF+79kI+YhdFhm0qodVtwqjMZrHktzT+S52cO4vpEf9phZ89xIRu16
gUnM0TBcn0WTQSgf+sXsm2Netd7HA/GZqcsVoNB8m59JQmLFkjCajQ0VW2T44byYQNk066p/5ymq
ElieUXAiVT3XXTPGzjtKZhBnhWuiQqeL9Wmo0AH71kesHCFd2p1doQRBxLfPZAtxtMf+LxCCPcfA
DcdmkGLmx7MV4pQ8x1YS3E0a5k+59HfGlmnRmRYnrKKCBIb5aGr9lBvNdLqRqW/9Jg4qSSIlOEd9
U5N9oSn2C+q5OLdRtBZys2JP/fjCbOu4x0gQslk3JlilBwg+IKTfdn8tECB0LU8jdpg6x+gajnYw
QiEjWVGdevU2r/gYwiBsNCtoypbBbrPwkbO/RvxjBSNTggQ/8YShWWMwHuYleWP4EhhwM7JHnGPD
vx0lh5UT+IebHU7ZkwuCG5zmRlu2Y4lOYj+NQSwrpA93WReU3MqEtVv5vffpxAAIHU0JxwDgSKFm
GA9UnyCJd9NhHkybRub/ObW+MiMvq09EN5ZpS4jUnTgLCSiPhxi1KdSpY0gSnfVjBg3m2w0KjMvV
AjmYm1jUrnL69FfHN6sl0TZKIC4Cnzc8DL6Cg2gu/B+C01ok1MUMFbwbBXoie67pvVb7Xz9YYVgW
xMTkeTGvLUahwI/9jx/jZJYFZ6lcUzsxEPXK1/wUwpHL2HlH7gal3CD+j6Dbqfum/mM2iukq6xgc
iuzYrPDLARm7A4szoTzM3cCYiFrvidIw4umxyFLdY3xeTMMTUBFymGMLWBRBOoU7s41gMiM+wFI/
dKOGwD+Tbg4xZ1NkCUud46PFypS92XlsivzovqVan5KvBPFlFIfuuGIyOJ+JANrt7YfuDf8O71lo
vvkatZP+xML2Cqehqs0UJC7SQScH0g2AzNgTlXMMoo0B1nWSudEJSfNCia+Ge9kL5KqycMp6l/zA
mG9oZNwxjHqv1jtb3opVq3BXvIAJ+u0DN3+IyYiHRjRFh+K+RQaF4F1FTs5eraOZTSCtgIaUMG+2
kP3ml7jQmIBk1EeXkCkDMRcAAOFfD0Jvg2nAPI4scuuGy0cem8XZ1UH8IFTvqjHeWJdWgEMBKq13
I4SYh6pB1xWZANPNk5qcrM9jIpZtQG8jsBQ8mU/4tCIuTj+CHE6tBcUOw7hjzG54ZEm32+r7D6BA
AMlvcDHBrQSU/B2tazc2o7plo5gKq36UGQL7vwp3n4jtLU36F3swCPdvInfP+9nrSkTfKNs7sTQn
0ZKF/YTvj0aMzFehnQ2DR8+heGsuoSa8In2hKuAzs3CRd8KWdsVg8KZEJB8Xk/zYL+mq3/safieW
7H1F5nZgapKoLUBynXqYiioTfmN1a/DgTXFukuKk7Omu4qnMRmiBuuRWD1gp00owCM4fsVpXWrMN
osh3Gk28nH+ne/UaFvzruHGsdXbhWYkFmktcyZs4WH8jh5mnsK7M7uUdKAnzfFEf7fXHBjVjyh52
yyUiCYy5Dj/C7yEKpgDFb2mEs9z5K0d3XO0tTTgz820FBK5jTScGVtq3KSIyyhOD2CuwETUM1vev
OnDGaDXZHuqJqqqRIpiQ7UREGB9BYuFIDb9OHF9GBY5qxw8tVYaVt1bQKEFQGNZScaY9OkLsbDGh
7WLh3E2IkbcBfi2ZDJcwrMR95A6wXoyaX0gZcZcg8DdanXDsxcOSdaJTeSPYi57jdazhZaAR5YkH
OaGaFL0Y3IPUYxrkfHF5CKQwu/fgusJdIDogccvfQO09nRm5HNsm+TmFsVo0zJ42UHchZ4gdjdj7
7UX9bs2zQUJ9q1mSNkgAzBU4+8pDBBvqtNsymnUTSrlEt4QWw+7oCfJvc1ohlBwUau+yQ9UAi/Gu
fMxF0KbUDRPZv6vX5BZIdIjjihwzmQ8rnwX8pLIW0M2ZDx3bUEMID5+2uyuaTKNSTUZSAooqhxd9
/Jc/IrYxsZYLBiU5XGEuTFtQ6hOA52xcfXmuF2zLNtvyqKo6y+y8vUfIujAoY51Q5Ubiv6uBJnnu
FpdO/eiB4d3qxv55yT7JRvIznilRvZP6p/91cQYsi8UW9ai54lIpUQVDquCy+KC++F9VdFxQRVC1
hTnm26aAwjZMWsZkTdigL5eZJRuGHhBCHLCfR+fbExeb1QE43WwF+c2/QW4wIpyebC93X0mxVeiC
UqReIs63/4m2tpHBj4aTiGtMrUdio8FLh3Fng5xrGl6RSKWeMQZwx/aHLUSUBLcaCwuLkxNY1qBU
4i8jhYsvBDc6LLD6feoacwpyihDISks3M9MwhBU+xi9fxOFF5CtiVK43y9oWr2x66HsbO54sYE3J
ank6lNRMxPNg0sdKLMw8YhgrWoHN9aI8XRKmINHQ3p5IxD2ZorEoJblzNm+4nuoL2VadpOe0nYZa
VOR3WL4P7Y5oG0BmclJeOLHv2ADda44Zklz19Bh0lCNVqzYRm4gxE9vI553qjrxeoFCrqamOVoFb
PIjHK3LdyBPDx/u0EBx2S0Qgs+hDvjCtWPHYMkn9Z/TN5wIGCpHXYTCW/r43SFVqKKNDpbKernUm
aiwfP1hMrRW+X3sC4Pnp+mghFvtvFs2cy9KepvjwTAJzu8dUsMEsHsS1h+IEhxKdSMk32jWym3pC
du60rpl5UWP2uH3lIMTdv0N+agywrBzt42RD/6hvG3IUBH2aPw/IXJOOrze1Di/rjy6T0o3+vKfK
qTtbsaUsTxDPfGK2FwoLZGXRBxJMHsm5XHA8Z/QDDSZJcvIcZIsdo2YTc88YyZbqwDqOckUbLOFd
M1L0ZbPmH/iTWr5TvE2TCkVpiWLqa4Ojyhdq0rKbu4mMlRksouUvAJBzdWtdWILUeiahySEWohlS
8mj0RNJ6R8sH2aINZr4IU7EK0/dfbmMFu+ALr+Y1FrIax4XH6P4/Ct6JL+PKyt+IUsX6QW1W14Lq
T6r3U+KHpskl+fCOQqLdV2JfYJIr4JVZlS1Q788NyLI0lpkdZ/rrYU0Yg6lROQWo1C5Rw6JEKRVl
JiY1qv+rkOFBo/oDspbB41ri5rodjK2YrZfm7ueI0wwnw9XGynzmNpKqhwnBJHwtvoy25A0OvJG0
BO+RRR90DYf5IOtfuBPHWVRtyMem5far+lfp2yxa3wVKSumeqh7uvA/ESr1skm8W0jyd4gqDq4nx
+cRuzPeEG71Lbu2Xvetdp5Lz+6piPvEeZG7PUMqXltOrxXI7dhlxDTYoFJoe7FTlqDBCkQmHUfcz
UmRQxKjsfHiC01fca8gLYRh0u4Pjf1C/qUg2oFDADkX+xYdPQe8PaXMCemSdduBmDIO2Of9S45Il
sKQKnu/rbLseC+zRyqXQ4kMrO9kKoJF25yAqxZHeIwkJcZcOAkXpt42869jHSvvtwEsTo26Io5J5
r07Qv1V7A/v1v9WZHXOsumKnvcTKs8JCjzIVLuGJK0iaGcqCk3I2BX4DryHRrxPB12ejfdrgoOke
DHh9uTwdsqlM+OgscaatmE8MAYiFETPpsqhLnrZU2DEofS+EWlR5DcHHKerxd+DN6NncSJRfzTLi
h+BPcw0echrB10JHyNUabK1OC+47ln9M1jkb06SxiNkrBTxgGzlR15i6ZiRXB8fLOhvZVJMa99yR
MrKR8Du2TPfd60dAxz6d50weG1edyUvkRTPnCpc6FZqC6M9p5WA1Pc8sd3pcLD0T+MQ9lKIRSLss
xpB7i9R4Pg64EQgSPJ+ika6auht76b8zO6sbuzLvOzMFWnYaJBpmWKpXMAS/f0AurjYSPAr0giG0
kf5jYCMxpCk18K/Y0mcAckhqrvHke/NCpBFCAAqmWNaM3NNFxF3JT1fLjcCzjpozo27V8syERNSa
/kIQZNr5pyQpn0pQCf1oG4NYp6tzLTqg0j29tMXNCp+CsbDhhusw3AtMtBK4maSohkPcx2MSustW
r1rgcQn0tVeoP9jsohr1sXcXPL6mbG5nPxVl1anz+1NL96H5KGDbRLvROc8mnDsOyMsGOFW+tG4+
700LaTOqiYK6/Z9XDALAxDt1Af3AhW2AWzZvIaHLgHTpg83wsFH+NC4jVqY2hLPrb/Scqz3sRVlS
R43esb1ssVSEFeYuxhl3UDsz7DZvMY9JZ0Jw7GfvZ5YAM6P/yTidLaz2dnyezrO01UgTjbi38jw7
GD9g1rWyoOceM7kBN5mzd17h7xFdW9Imc5zEnbxcyM0oGC6Y9QBPFuU7xp9Z7O/xtOl0wnSyv4Y/
biewcCzGlNwYRFhm706uCa/eTDB0zuRa/tgpYKPXO+fFsZ/cjTcnYEDF9kpcpg6kq487SoYTZbjP
/JEscxLXCll0/+BdpbWL9JrzSQGyZYcRsCXjhVq+t9WAruHsgj+9FsXBBj1ip3LA7m42kl5novS6
As/6Bc+MTekDrnHFZip7qAEhhi5OCIbzEFWeARM/bZg5JJqK77jlxewY9D8HQu911yrMbZX+JfwG
Mi/6O4FTEnoA8lC2rt8yF0vw+X0+1QyjbQuXPWdITr2tDUgXvN4LSEaA3aSa7rAmg22ze7XJs6Jr
d6QLomUsvS8xiKe0OI9U2eXYY0OV+aX9U0VJ+Cy3nyhgBPCzCOBrckrmjbNCyQC3cr5xnRgor+Bc
8jEUcE+dbfGfV6alNXUT42jmuZQQ8rpgdXsUThNKSoBj7f98JnjTwgj5y2pbAUkUQ75X9lLTqfDa
X2qqapWsMon3M08QVkG3wKMf05zhl9h394cCQTMFn5E0Z6Ggw6mhe4LdaPDh7V1RhxGQTUkPlPsz
tnQQsB48zhURRgV/+X1TYR6LZAQzMJxODM/1q0Xuy4FLoA1jeh4/siWbKiHOL5O8mcYLb7GwC1Ke
PqZpb5CH976mCKNiWIWNB2YHqdqrQWghljMSRHxC6Gbhqmw5sAkCKhqaa1MQE62FbgvzgEuTXX74
F5zaM2zNyf6vTK1P7BgqKt6G8v3K9GduyLp+T0cISoNdQ8SlaTst3jK1fS2syLx0iibL289UQqLX
TKkFv4hTWyk7V9G0rDux7G08mnEOGvOWnqNjEfuDbj4Nel9n2/cCDLzp58pGwSGf22+CqZJoadii
6L5r2KCDw7wnqTmqIEZlm0foivWDkP5kpx/g5lPRyPMUeue25RxnrY8TUS1cp+IbsLL78h6+QDDb
khdI1MdGRDmTmyblhYmUnxgdRKDcJIJKrjBtzGBSSi5tCjAvcQ/r8AsELQVNrmvq31/kFMwfpAOC
hcXABCG8x9y3L4Av5ZO7UhmNZ4voMnAhDaihmTQHHmQZqdLCTii8nc0dIA/oHDB1WIaRUpAY0gkF
oM/OFy+zyQN/l5uddKCilicVvbSLT18hGgmSkAP7eARmlRncgCrWadOSWkigduma1HYdjT0I8un/
9gd5kDtpRouHpmTmfc58n5q1OiGC68bGMqpuyi0KTNv4msgzL92ce0oqKbQgKj9Tkt26RjHBbSYU
xwrRDI9kNt9BL40imF0vFsVIwGlFUm++zhRGfvgJ3qdLIjKkCXGJNW1P8xKZ0h7207JfQdPVYhTF
m/U4YnsUkVRLGZbAUObXNkd9Bwf/LrfFjPDFn7WmTQb7gHuswuB3qeNqmpo3AIh+YhairwDyASND
bu0c8cfLkMOu5xogaAkRnRpGBBDF2hOiZNsUGPHyDM7UDm4ip5Axp8Ou2WYR334OdC6wBCnZzLPV
sYDq0OcPg+4lQlw4qalFIpwlSy26cbLgjXCLugVCmgv5PQ6gd1pj8Qu36ctiR2k9i0oHpzuc59t0
jG/uaD4FE0cLRvMLNHDEC3Hufc8e9HxPflUyeRPqMM7AXofYyOjbwsAIxgEyKxYWu7qSbUyImg65
odd+U/JGeL81oQKI+F/iZbmw/Coq4DL+VTmyuBBU18ErS6BStQW2ugZJD9MaspBySrkXNfj9zjw4
RUge7E2PMuyKWD0+Agggt6Mcl1TelerxL+O1oX4EBXA7pFVY15gk5WErpVZeO9yNo/VU2epLlBFG
sH26UiwmcWGnpqkkJnYqv4ICLRzd4vM4l4Yl6hhqI0VdkufpXGCh7WRwKHgnrRq12UBLKAAvM/7i
WZj8tBaW5rXXhCFL8BEOYUFuDf0dGtdM0Zs/9uSIyDgnwTaoABa5PekRen1/EjzGncjQgpC/d5Mt
Z4N2stVmU1RVUqmO6Mn/JDX9ZKvJtOj/OqX4ycC+W86bdcqXMgkMO2k3JLjbRf2278kajmkN6IHl
6o7cA4KW4ek3M1qdFEoM6pvJsaAaBP09OMuIbyGRzjfmCB6t71QNIELX31NK00kvhejT6rdMdhnM
rpta12SIpZ8rFt9yuBhCPsrHBZs7VWBN9w9UHDq4cENN+kQsakaxLlHhW3FnP/0Wiw3f9trMKr21
sKqLrbsW1bAB7Mf7zd9vXHzpHnzitzS6765spCJNGxeC+TDLNKb8B0KbLHt0yjasj1SyOiS3sC2u
avkda/NniX4yNwsuW5OxxzMuUNMRJN1UmjVFdCO+6eDuFgupvI/qH78vkAe0i1NkuqxzIrQNWCM9
VpccfDzJm0P40HIIvGSM2cSYPA9teC1Q3aGG+NRF0GJUOIVKXYj44PhCus06z1/DjsLAvMa6h9EQ
IDOc0WDa6GALYqwIMkTL5ju12JBPlObCzU80qAPEcw+EgAPqSlxrdNkN/VDkQTWkxiZf0YFD11fF
GrO1haWLpamnD1cdhqQa68Nk+2yavtTzFrYRMCEL/lw6pgFiMMRkPHqMihyHSbkJ+ZyAXojLTByt
yJVthsVaDRr9g11zjB7wiUizuLEOCcSmEZ8AzaDSE8fD2ttE2EoCjhrL9R/SDWUYDiykjLLMLU4o
U6bwAOJMEQ+60ce6Ws91QbReFMNq+W9BdTSBA5RDlvP+rS1rXZzybEjcbjbWEh3BbBHSRKiwT88R
OIaYhIKJOhwwOGvC/20dJD3o2/kyTrO040IfNG/8N7qPHfLc3GOZGDO4gDgFBUYZAuNhONs0aNSr
NACYTzognopD7kaqMmsyQWT+Q3JZm0kyQ2g5WR8u0Y8X/wU9/eAI2djmiuIBl6bzg3ol8FpkAeo4
kR69ZV9EDE1x4xbmDMx07WxrOb7BEgeAd0LWJ/YkTTcrbdToEFV46qIxjA74q5AZeMCshsW7SD8S
Qx92OvNFuiNNe9UnIFgQZEOtg0wcgWiLISNhc5sj4iIjKLksNLOnSBSnCqV6EZkGbseB2KZvGR7H
kxlt+8EPN3Mgal7BEsoKoPuvCGKY2JdSN3ES1oPir0CLL7xk4tFhHDBVpI2weoxJ93jCCtHqILO7
JqJuTu0+RVXR3qzculg7GCbpWPQenJKV4OwYeM7CGu/1T3QN6L5LZUBRsFXoaSS//emqVN0y5OLj
RDnN1VYRwCmNtb3UOiWtbuIfKp5S6L7tA5o1Q4lzkX3rw7EOjJJkh04KBHcMsMHmNjhE16PkMHWq
VabvALz6zFxqCE/o558ykUnIzQjiRM7qCJCuErU6wv4d0E1eZHqubq5UOtcYslBVGAHbWPtuk2eB
1Cf0t6WMTLH5q354Hir5HNoCngUawncQ/ATLhAK+uDXYItu8+ZWAdcWxwfbDCPT7bpFiPAKVOFuf
D+Bi2VifcNAYvlhHp5Mue059MVIVQpBn4aa78celgSqjy7jbK6y/bA3FbTdb0EVZBg3lurBn0EFW
SFXYgAk9/9qtkIvtfn7jW5QrSd/TwZ8AwJpohRl/ON7mqOE7s2jjY8ykYip7asa+z5q7onvXpLbL
fMu0rnAbAfDnEKMkvTdpxghLpHfvjEPz7zCdzD+RfedBS31P9qNujNRQYxmR7yCScFlQ2s75rTht
es++HvLua5Krc2SYh5l0AO9jq4HpID7RZpcUbQaAFUT5i9eFO+6ae1JoMx0aX87AMlHlHxRNzJYf
mH1z8H6jUWv+56ELpXIjDWPknNLBX0drRBqHaABe7rWlI6JGDWRBhtX83c7D0UaN4R3LiryDR8MT
3ypK7olyqBbS6D9E2Nu+5e3iblKiMhVU3+Td9X+Kc+7dL4ZMpxu/kUQh/99LEQHDJSZGrjQQUthE
7NhWs7QsuRRc/GzYrryWhp6NJuocNW3N2cDvBdO+dUM6q9gxLHp5KpXVw++6aMxt/s4qMQvz7b4T
Tf1/FzeSkNmYQw8vQTwgy/1twKVZt+wwcMqXucE+/yZ0VB9GIne8J+qxPAc7S2dK+Y+fR5lixZ2Y
IbMd+7U542eDN05uMZVLlWJ1cKssTCmueHxQQb1p/9gA8wsQL891xzW+5KhaH4H48QWVVA1VLjAv
8anmF887E+nn4jcwXqlHwup5ZcA95BdL/uy7cyC7pCUwD+lO3LQqs2dVmldBqfcnePY1VfM2QrqL
Lh4rd29hZz2wdmSzpl7raxfNHlqCkGmYXV7DoH73uKnIkHSic6BPv8J9n47OuFyS5sj4BKj4GC1t
APIofr7RWuHzU2QSXq3053pHFwhuMzTzv/Dwk3df2M3B8OekaChcJDDNCKS10xWKIolF1qEL9dpu
IAeW908e7ay5qkMHLUuo9l0iV5xiU2MNog239Qu7eRhhvnBpR1L9kfgDpq5m/ITsaPDelNcZrThc
0ijp4d4shSWYHtIzGKQCa4VJywWnTqds1R7SkvpIleScsbkn76ICHrnANtIE6g9lga5pfi8Ov1j8
lq43OQ8jmyGlXRc7fVeGSc6DC8QBsgm12twbdcoa13YfdrS7HePmQxArwfcTJyLPQOk3ADKYhzbG
T9rIVaz+WWKDq3MBnhfZpZgPKx6M+Im8yszHo+BcT95V7ETqxTUwOsB0gb6RW6WKKHRdvQBa90bL
/RIPYkXiZr5nv4iPUzDm7sUBpZNs1m/M1XA8TjO/q4YDjM7P7qpN7wJBjQcMjsFYEocDDDbVycZs
pVxy7DFOb0+bWQGUsB5l219246SFQvW15X+oHGdfwtKDQ8oN3t9zUqavLzvdRfLqSzVfdEWeBXSE
n/9Lo15pUQ6nmMyFhW9XUvQdySTcd8Q48/0gQn8M3o4WO1MbrHG174a7/5jCJiUPRqK4s8Ymadm9
j8VLB9fcdATcfDaBxbT4Ovpoh72pFfxZg5wzswrROOB6iw0cjLjqq9jZfGUUW1CWd0YL9u8VaCYB
7UkUax+09XCS5CnJme1CfnXbT3qBRXjLf8A2SbY9LuwbJS7mwZ4lwi/rNMDzFxSSXOpjQ6Zf3Qc+
YnqPWmmJ7+z0m/kYPEyYeyu9hgrJrSZEqP+S4HrWQso6Lxa+JkiTvh5x6KmIzEfBBnUzqlCW/tw9
lM7OYc70pAWKgMnrJX6V8IEcs7HKq65FbARbM3x9vTGsfmH7BH5Yk76QJDraTlPaSuBkB7Vz8tco
5P/hlA3yeK2Mf+Ia/HDbcbgCql+8HGnIzqlLWeu2ypYIn8/jd7K5GmeOdl6+rm/uKgzVNfA2hfGg
BQ7ysfRDetgCRsSkRXAeisnxpOL8OSEpHOqz6n+LEAh/u8+2tYRSEL/Bu2rJ70X3k8QRnupjkD2G
ZZEStjwGw9U0+FNvjy2H8xNPo4mnoDbNc9MHogTi6Z/GjtwQRPdDGXKYwqAwSufXBEuAdtS/OYJy
ykmaVLTgLr8XAJxA0W9XRfydQwSDbOZix3SWhRjXvzX9M5stwvMaQPSg8s+holk8FxP7p4JusuRV
Xbi/V/k3vV/w9ewW0R1x7kcu6hN9ioxWK77NmBi4sfFaIGYHPj5bm2hf+fwTQgB7583U6UP5wZJt
6ESeiroFUNTENzPFGU2RWCg8y7kCdRFHSPa1EJHl2zuLizcfBbkEPNOPL6zghjbYJ323WdrZOs4s
WKkc+miki3MmISsEdO3vyjnogukt9NOE2+TtNdbws8zBfTnV6YjRZvgJd6askPor1wrH+JqXnMw0
ertACJnrL/03S97zGQgSIHBspzndr0cgmNgcXUtbUTO+6GxXFJdJbqeMadWtSJHNg1oQ2NzaMZHX
jE3afSsydSZIypqPAP61pYQ9ccGyv+v8bTx6d/wdpS3eQyo6cZdGASsPmImS+HJwuggXP/MWt2YG
sgyQY4wfCCmDYKA4Mdwgl0mC+NqaZtSEHZT4nFYQlVFgIIUfQFqfqaScnPXT2gjLiJz0ADziSB3F
4mmNZb8jZHby0IN72E06R3EBuUzhPIrvQG6mrwXcuhphwLpoI2M3qyU9iZ79KzU80IW5gN6Z2eBM
0EW+NK+OwbQcaMRl07i7FGHJWkPHcIrgh4qdsZIikOYZ39xrNJoLQUDUVWj1qNCseIPtYwfGS459
qniQ8s5cCHwH7lYs65D8fGeEjCQucUO3xnV7mS/Lqwj5G7NcZIklGnGeJQK1TGW3fn71F64aCldk
19V7GECK3KrhxzTb18oYiwn00keLwjRxUxhO9qDoLgL+N8AP7HMwjYsurTGbW+tjdWbjTl9L+TID
2ksGP4BbHCqZKl2Ompi38XYQlyMA/zhtuNERMo750OcqfseMermmfxYB/h+F1AeeDXjovXmUH2QT
H2e7O6L5zzY4BxCYKDRgrq8ZYd26YX+FRruc9t/TqEvkz/kJjYf44q31rQ0vxNNDf8Msa5hcsaxw
ufAlh+w8at5fenIfcSyn26V83SQQ+kLahw9+k9+YEjlqFgZms29VyD52EERVTaHAyloerP81Is9c
mbL2ahvxXiREGN7A1DK2lRZAdZc6zC8213biBhFtKzF9QB2OLDt6XBTdSAmVA5kNJlYPE6f6zI2/
4c7lwt52g2XLPknqnNlU6HariUbqOtjSzx0Aoq6wZzr8NJ5PijvrxP7X5oAu6lXbODhwEECblWMr
HHUTldn2clOCxr5x6B5rTQIXP3ELnorhl6TJd1NnJhvfqr+5ioRfHVInGhkgjYI+1yvIzU13pgU+
G68rtoaPEQHGicP+6Em8GXS0S3WY1h2aUNYxkfjw+b3y/JlFdC3JXw+OfV/Pf71yc4aklb1pz18F
INDwfVFWl60Jsr6BM9hF+wCfm63cjvLiQr/1iIT/SBQyhH2/LCoKbm6HbeIIA35QrFxbTYm8KsfJ
rfMUGP3wAWYyfcTUHDVrGsrPCtU4Auww1giVf2b3qaooxVrmZDfh3VmbuN6yZfDAYiVEEKdyjj7L
aoE7Z0FDDEywAoH6Qg2Umri2I7iLL196szMbQvtwore7ORL9Nz6aEbCbTpVE5Kv3rLMK+lrknJgY
mx8Gem7efCC+sUpBysblS9DDNpnB2b6QdJN1dduF2cIHvK5INIGFTlWjNWohXtQ//FHTnYy5TcZk
qlv7UB+D76W8gnD3a6NPZpnEEu4xyJP5DF0ct2BRiTwFRDLkJ9+LJQk3oZ3zi/AMiWeqWANICVjY
bhb1gjdAyd7R+cixay6lZtQxKV+XU2N13+ChAy6WFQvfxqIks+EsNFp3+VhhUeizsRBuCVe+Ekxw
wn10knkmadqL8LwAu9ZLoPy+vQ/zw9yP+V29lMyKNhEKDsb2G9b1NmZCRcsuCOukkS4LSHpyYtwb
i70Tyc8t2cNP7PdMk4sVWJR7s3O07HIGoo+xgtHZZjvVMmiXeHuxWzN0yPbJRG7rebMDyIkOxXPb
yfMy2zlUnbyikfm5wEKM7FXyH4drn2UeSQM1e71+CTMeH/bng8ZC4KDDIQEcxLZEwxdDpn+QLe9R
CbGE7hSeAYJaKeE1oem4Ojq2oZ9HmPDtKP00ZgP5dQwitDyFomSfv9NqQDAZs/AuWXYEgC+9xHxZ
P6Xk06vMSmvBffNHtC8QEZTD7ncYExHWHGAQyeJtzpm7GI16rqs/Y4FtGeovYHQaqfK3Hs/nsIFT
dnmn1felhTjbiKKPhd1crXn1ijnXgrCHVGP4FKG+MpzpfWichKY0+doQpWTWh1EUWgc5LokRsNrL
IA+gjxoBNVhNsIiBOzmy1GCyes/jEqNrWeLWYD6M06GcGQ5c5XCgCCKE/q1FwLX5kPRlvDmzuv2d
2evDErHC46QXaIbDldCu+QoVSLnB8PlquSK3mxoYclBPG238NS0jHc/W3RrTL9xC7Beg8eg/Om5j
J2rKRRC+R7ch11thAlVsq3p7gAIQO8ZOIYuBq93L7RSV80qIDPf+6QuZex/bikdudPUxvdklz1Bh
8bWub4egnIvFm+dUe0cJhFhxNkpGAdX2ldZ07x6EXnXrlte/CDId/irS4k2qg7XTvcFCOtaDX+0h
djrn+8leOfJQj4s2GzJkJ0wfbJDm0OVspgNvRzj375lme09EEfjpX2oo9zPEhKVObc8SavxYlnxe
a3FxQdkgIrQHaCtmaJixnow2UCQcNNQuty4OGW1sejo4ram4xHrv2UbuiSvjtp4Rl2qC5ElbcEHZ
ylTaXdBuNNiTY9vTRmTS1G+kTCccwxvuWrfe/8a68rSHoHvyefoRPVmFB5OPWIeso5+4jJifGui0
1NvxQ6nH6v/lmYDNWv5rtp3qIdD/QWxv3C8qi9C6sjkeqnFbbR80JKdSQkjiAlB3jN0z5KV2+loK
vZNLi74DKSCnmAAG+wOQtF0/zfesOVvfC+YmcWQpB16g7IgNcHuaTc3XAfzASEIMJAtZjbkq7a3d
FuIO/rzYi7TYznh/dmJoWHitgm5jpYTnlgYrR9N6A+Alg6NVEb+SQsY5d3GwU6mZpGy7JEK0+E20
VkuZhsy+rhWzYMMNdET5CA26gzEF5seg8t4lNdvr8pb7NnqXXawR70BtOz6eVGCbSjiL2Kg+duhf
Mc1k82XMrABv3H3LEzSIeF3F1sppxZQI/tfvkBnpvqVYKKyt7JevBVhqcJdmeDp7S6OASTXh90GI
J4D9FOc6++3Fy3ZYCVLHQ1xpjJZHExeZIokn4WKFXSf3kgDmuTEP2Ch9VMHOQk0AmFVE9qSDyYjI
G/uw8A+NqPKRHxNLBOI2lnvDcskAuXTtWuoDlgor/FsEd3jQzpdc9j6S0BfrKTaIyICDnCnXOWQZ
YufrQrNcvqOmadtgiFTETJ1/eMYPylW1snXO4SyvyfKAhT5zBhF8BbsyDNjrmPwp2pnx+pddf/Ic
EM6zLMQAPsVzMicBd8mqtmxN5/CYxLN1TE7pPcpTYtm4r8c6RZnxjxMOiRvzZqZ6gCe+OiUjQfmn
GpahWzi+uwAWu/VtYTeD3tTpIEZL7FmhYemP51LrpbLRX/bOq10nLWlj+J8Y59kkb6woUhtpa+op
Otq+qCqwddLFh3pNAz8Ec/Vlwh32oDSZ7H4JUM9JfVsWfZMgP7dlV/7Nj5ruNSqvIfJCUINbmTwS
vT5jBhHN263f8fNydJcKGf1QIC5zLPLOM84p5lcGHrVN7TkIF6+CcnsJLQs4N0UjYB3Bmh5DeKMh
IIFTNbpY/bWkI6anUTkdEwEZB3qreJjTcdOZ1VHrESS52Xb7L7JjmQVaYeK8sPnpBp6GqAVbCcYA
zH4Lf2+KKlWINWMfvTVjDuug3iXZ1zi7YxHqGemLZkow1QB16JQiUiyeEuvZAXp0e5gZ26EyzAVw
HpJHI77tz3szHI8SnQAblrHYqdukCj3wvCrtv0460pjPA9kT7Dqbo+KJPU/jYFBee3v+8esvZysx
G6LIljvI9cYK5ilYifuLrK/LFOLzPESF2stnOgVUYUBUob8Z8WHnE9mY2Sfx+L56kGcPFCnrSyi6
qKpuhuO9ltxeWE+h+CkQYikYXBxMKGfZq7U5SDdr1KPZ8lG/jl1DKyrG8hiZtG6Uiu6zZnN+cKkm
2xQhSpmbVrRJ7PreoiWJxIoyd9BNnQM16EBgfUlGz0HBdDBxVE68XJyYv7K1lkvrH9bMvWNh6dqF
Dlp2sMdDFy0jlH4axKFU6FJZHhaOfDFdjF0/Gji+kPVcV8s27j1HZl4fqcQpNInmmETHryIKJhRd
c2X147eye1J8mdPBdhruEGBo/v0QHlyEsrmPsTaQ6v/MSqfPmPOQn/pyExXAzr/8Y1vpPUtq+ka0
10N780tt4z5Pj9sSDZhnUvObThnYoIpAPwNpAt5Ie1S4XPvpUOa1P6WgOkXEmEk+Cv8teQ3XPW7M
q784wqaKsxxk09j51KyBfzLPHXKweCMqJCoxxftX1WM+iPkeRpKxIlXB5gdp8NJxGaWqVHGmNWA1
iZHNiJQTsqaAqC31HXNJZMOsA/o02DwDbWdySB3hr62Z8WQJ5AnExJr3KQv/MMXSvLUHH+pPia70
BKAjSykvLd531KTeQ2IevujOo5I9tUzYD/xCBbyddffnDhNmoS6h7jrOUSrVZDgKFO38bC2MgT3Y
zNAMqWxXfaw8lvg0e9SCRG1Vjo0LzOaA8IvA7BS22JPGrnLPdsSl8tUJV4O1GswAQbjcTIDwN8dS
p4V+TZnuRDOb1f+LvPyGfIO9rdD/XortCnFROJ1PNWndhv562uLhBcQTeJuM0rFoQ3Xuiamj/kKT
9az5Md17uEuQlFzptYhQmJrkN1gNPggKa+go5780gZPbhCOMKdN0dF+L0E9O7JnZ5o0o1cFTGl5O
LkQvTGqTcoxxg8npX5rbpb+JvJbsInnwnj/wUYNLuWvEtbHGwgxCkU6mF4odU+huli3cx5tpJqh5
Ch2sbkW1pVAZFxsK3tWBX2/Npxh1w1AzZN3gvrTf/OvtbSPlK9pcJpvA6Hs5QU0wa0sxqsPz6iEU
VlJR/vhAtE2GBHNXnzx0FcOS6F3Ac77ojXSIBMnvhK+gUJ/8ONbPwR/7vOXitbGalubAZeBG6VNK
W4i29QhwVp7vIJWfDgPqmkgN7rPNPl53QNtPOeHLKSKIuIQ0+BKDtDp7imtxozwCR6Zsv/dSLOfh
FMv24Qg9tyRSktI17Xpow+YsWqn905rXhqMads8v7C/W2iQG2XIqBVhLTCDXj0c0cImUDvhg276B
EgMoitjANMsTOpBE4zM6gzcL6T3VP1Q17dadvCDksvmEEX2NI+niZh0d9mSLLvO0yy0JcDMXo8mi
14o9+ExaOaAxzQO2g8ekXSlbZCnz7juZapmncfUUplbuRIUpoOWBaYxBXuEE4zdKAGspUeL4CPPM
LA8kbuzweY+TeSs8KTyCQMdNZll0/Cd1imbdLPhz7a9+RSzf8iTc0pnESEbT6dvubrHHc7vZPcHQ
QtQl36SBIAZGx/Ucc9tsC77hfbijtFvWMIpn91utrKY85LALUqpXVl/eMRtKEMxByTfNp8yTwyhc
bH/ou5+xAJDVjqZp5GgN4rcuOq/7n8cXmZsiBNWDPI/POdfT8rT6PaoGu+8EGxiDf637AG1uwBiB
QzLN89n62vn89y31J3p1rb7uLIZ6lvfHKVh7ci3DBKA6AUrrVBQ8da/PTvPbncDFBfaJsn/7gZvY
l0ZzVol4R7I/3IZ40YISVGDOEm2vJXV9+m4+y+rU5D4HOnfNV1WsT+zxFtLiUWiy5NZtcEePsIP1
mJ3I1Ai0ZKBuHH/BzPLMUwwqDL7ygqbrACPXMjLymSlpHjptg47Yhjw1AF53P5dnSsChfX3uCdpn
mqojLOVzvXMWUnDG4UgrQhcnGOmCzGc3Zlfb66EvO76yeI3lU6gsnzYerYo9hh9zWTgjQqtqAfk/
ZvtIjw7iF+uVoh6dZE8FHFdyrO2Rtco/XnFaFOf51G+Vc2sHqSr5peqM4+BQgmUxo9Ndt0GYdk1+
3hyWSCxKrnebMkcaQ1qZMufx7WTHuo1o2I4VUa1dtSife3GcKAjWc67WUmzF81Rvmgiz/5AdSgeZ
bARPQeQqr3Vz5EdnVd8/hx7IKLyajYQePajsIBZlF4k9zAnu6pmNDY6eILrDwfzfoYTHLgkHMhXw
lI3/l/hYxSjBGFxWYK1KK7Cg7yD90FY87hj/CJ1QtWm3HCIssHtLm9ssVsrg6lYS2bXP8++6IEuQ
EFUT5d/37zz6rSy/4m91vJQOEqc48TO3/FGPwDgwAQjKahFQuxA1eIOJWcDcQ3kQJiEVupFCWr8z
tU/jOyH46Wk0P9jYmM1HOvGPPi14wDH1wOMxksJeltPWTWRKZAUaNK4Piqm3cCuRxdX+m/cEH9VK
u3S65IBi00n7zwxb3yYbjN7IqVl/Dj4Qg4ZTF9FxVdx4zjdV6hLvcAeWu3xDyultjAWLgrMYU7Wk
ZYXi5mS4EkfRo5NBdgjy6bSbla+kj8/hDfPzxxaX313xJwbHIO/PNj3ysWSw7MWjQc4crPhbtMcm
UYToaTgWtrhQSCFJsDJt2UmtBsS6PrZXxXZVYu1J0JEDwoAJSm0AGZDCzGsabwNpzyjDr4Nx4nZK
fGQczO2sskzrW+i0Zzn5NXu0oiGN80JTtLZz+0qBKZ6fQFbXR0ko68ywEonrXQ0mrJWsuWSemM4G
Fbk0U8Fagu/sjdNoxiVlhKQ4pmtoMO6oQW1/6PpFG/bCbDXrOTKNMIuEj/yhTu2o5Ud0DJIfjdjI
lY3HjJsYQA+IVVvOKDYCzaqHYBc2KblyiCkXxoF1uOquSy0hvYHCKCKrFrOWuZ42I+pTFuKSaYbT
cWh//zQYMC0nSn7YWzu4hQahnyb2z+4hZZo1q46Oa/5PmdmRPkdMT5HwO7Wd86ypP1cZWW2Cs8ws
KUm4DNLlfHy+P9ptU5TZnjVSTDTnc+UdoL1UkxrbiPj3oJdr5Bws/I/D7EE/AFIjr5Uoc5tDK2Ef
Z1ij6cmdUJSS7aMG62Ywsx1lHzGKKyiZp0BY4Yb14S4bIV9kWT9fzeIfmPqK1H+HVYf+9iLh1LeN
FtyIbArPdJRQJFIpxVIRmzRtgIiX+IYHa+Fup3y9qNQBJZunea2iuAXvKjtSa18QuubwRBjAYkdy
ut9SebyrWnK6LmQFfkWQzcmckf6xfKjhbVcWzz2u+9jamxLQmwdmWZG8oGEYWB0jNjGis/aCQvBO
Sjd/LmyqpMshB8C61MpJUw+gpXoJ33WJ3aAX1fEMR78ryOZ/EBnEvaKQvahE0RJi31p/e1tDrexP
Jqs3y0IM3xAmeCXhCkMMCW93u/U9n80gNx88aJT6Jgc5J/wbSFAE4AaAQxMBGODpyeNvBAcWftXY
UO2LHMTmNdykxlCn86M+cutYFwko0/P87YW6RQltdxz7m/k0W2/OADP2NCheRkyrW1q4oFainJFn
A0MR63+4H98QEf1hsOtUnwV8tFSU3uPdHIJVTQVAZdYOA+jQF0DV54xDjwMMohfDV32MPeljuDLR
/jpRxgnBIy5+MZJkIClcLXhVToghRegAEvEyQfRWb5fjfRjwI3+X1r0Mj/A+mX3iW3VzCl69wseP
+zVuWI5fEcAYJH0zqDi72aT0q07trIRF30ZMSau8usPY3DvhCo8xnLu5KRPpc/TFl+woVjp2LCZA
JRgC0gpuQ4ttOe3h6BA7yMH4Qf/ONLPn8ivCMiJ3pTdIa1MpvJ1g07OoXGbL6TkGA9cmnfu72/30
FQalJhgeyq55DwI22D0uiznpdX6dljrPcdWSp/CH/e3tPCgF3FnWhgGO/3kr1CMMWj2rn/GhefQy
ftAFGAllrGg5i+0RZrFlu5PMclbw4kbcpjQ1Dgtt67kbYszOj5w3eI4Sbfxki54jQO/aQbBnmvsP
zjCUKLAEcxj4ZtFPyhieRLobPHSgJl81qkJ4CTyOTooKUjKLfL+reYEj7CvjSJplgoXalmddyqL/
zCdphtm69xMx7uKLw7cBLooqzUZFdsOHI9EAN3pSnZaadUSKrB7ncrOiBy4tkCwRPKKBV6ySCFy7
Q2fKX/TjH3fbZFPxzMojf82hKojjYLOxKg3org+nRrh7R5zgt0ttpbC5O+bl5pJAq0wolM2ZhVjP
/bb3LU02BwbMBzcXc33qeGUFU1jn94p4neuFXDNs8MmuaaAd4vfk7cqHjaDkMV5EWZyZEk8DfB7Z
SNTSup7FB8eKVLeetizyfDjdh4ZfPzBeNNdtNAnoTRuybOY8czGFb0IFOSd6J+pHKWQWdyhWECnT
Jkz76u2J9dq9H/Db39PwCZuxuLz2qXqIKFdIfn61d5IcIqGyVLB2ufl2tbth3JduH9CBuOOVvmxL
3UN0XnBIrBl/XGU7H0oj4uA3bUSLkXacvPKwhRibXHNFWWHmW6ljdb1QtzHcHRol6MVC5/2oXIDV
LpCZJnlx+JFr6Ij9qjIdx6zj4VR0V+AKO16/RzETYY26S7MT6bGqwoHqgdYekcKJil9ErQIowy/k
HeMIE+hClgFHokR/bxXM6NJ3Yj9+f9HyiA7hqUVAstftTn8BQVvEeKZhrmawcaQRYcF5JlJB2yEE
mD2qdqy7I2ICyx2a+nZq4TuyNQihD7UwK95fp/k2ag5QxEg6jP68n1GNpzW+khKru1GxArnj/EK3
29W3pW1Yt93tOrEmijaIIbTEot3rZDQj6KJ3T3spNX4NNKtWSl2H9wj3F7w1VZYXo3tgpriHw+Pe
b/uBOQcOUFzVDZTNk6jQ86zqxLparPUOSv7Q4d5PrVuPs5qBOD3EhbCsmTyzDYzbRRahWjfB8Qkx
7bi0ev9U96vgNNHWMH5suBHhzfXOx0IXpHLSxBx/uTm8x5d5tdE01Qs+RnxbFC5Rqd2L3GxiLstm
slPPcBjl7uM7A4NNV4VRglypj4nznrNM6+2YTgfcGpVuVNFy3nSyUBIr7aISISDfTulS5B+wZmvk
BAP+iJcVEd4C+xWojmPEYl/kFEDtfXavy9qonkHpAd5jYQeXOy5n4pfobzdWacb2IpXR5gFAJ7B6
hqqDi1/cHkZenaYaWupalc1aFX0k+fFabkdzTfOIrw//mknXDFcqKYjdu/tek6Na73tAmYiQGNXa
8DYE6WI6sjdr6q+E9Lg0McJlmv6ZmL+ISMxeyCS0+2WzfCbqaUQWFzg7JDPpSMy6aQW6nlHW9faB
y48sjbMpG0Zo4Tae/K9Hvokyjo0HSx9q1SK15dFce/8y0v/US+wyoYWgrkHjul4UNjMNtgr7Oz1e
iyrups8FhUr8NskpLRDtEN3n1pgXBJrX388Peatn1jgN9sZ92wOM4mP3v91WhP7YqwOnt+W2RGvz
h4VCtDbWQ+QOSrDD7xMOF5EeS7eO+j6TyB33IxADjItBbGDNAKOPHJSOTsJP8U8WMW032zCV5YxM
xkQ/dFPfi/dM98d8SlY+dL4+YjRfEbpA6e6b+dE6Mbdbklugwpf2mNqE55JTfPg46my0CG0ph4gY
FyR1EJ4U/RTQMzOXR1DpjY6j50N4uUBYWOMPw3C9kUg+Lpf55nPXY6yTxXTlczv58K9UyZOIBoY6
cjbkRAnU9g4eek9BVV2ankegmp2wo1LDaO+vlDARn+esNbV3usB6mMawndBbTnkIsGDFnGnaHCOd
BwfWjo9Z76nQr+CARZHArgm6Xwvokva26gkIEogI+iB69JGJpkyWrXBXsRtb2CHPz2Rr96DsqJ44
t6QCJTSJybv1ZN/gfMYt+QSmMFCGXuaOsjOIRWnNjeJ8ogFFXIVn158Ha95ODh2xTtEOohCj1lzB
cN/chEyi8qUrL5C0U9aWAo2NoHwR5gI5dqgpHgMlIHvrFu/n+w7t/6/6Pxvq5xR8PCCzwqZ1puFC
yvjkfH+Lg8+8haj1ZSgAD1eLSqjm4nl7XfUlsFE42grd0DFzOXXJeeBdIawN8Q3aTwOZP+GxuxYN
y+4mJ+RXsG3YrwYReKFyrUAxofYfny+by+lZ8fNZ0v0SnjS40Skgo48DkrWwuJz9idbBkCNVgvwb
mJFJcyZdGxYsxJvTCi4VIVtJMYiIB0oIh7M5T5kDIJcFDHwODG1yYTvMvq/2FaVKrXsFm48cCDDe
ZhNkiDiAt+P9pua2zCWitxshi0exJkt7gRf2G8b2TQ/nBF43dZZ9qy79BmW8HB/T8qsB9SVxUDIy
km3MSezuUpJLF8H0GgpoaC8rF+tu0P1bTja/Xmo+TTpeG7lFIj8l8pAH/+WveFG9UpP4lzBQ5e3t
lrjccq1CxXv7AnJaSe9DJU5NERdnASOWQG5jk7gy13+HQzNgQ31J/IY7+YVNYqhsDXgLEdfcIYBC
B1eOJ9rk7gRRNW+95OBz9T3c0rthEPVWgx/l0MMPyXgyNUv+8fKxX7yn69s2TAbSFJv6sq9R/ccB
xbBP8TbOIp80Mj9T6KkJAFgVCyfo9dCF1+MLADhPoStOhnEspMK3vN7W+gqMT5G2O5Xhi1djKPgA
4KH+QG7+62n1IaKvN2C9tGai5FEx4oY4PJSBW0ofw0giTdTHfTtZClx84sX7TmiWYxWs1brqiZfh
MNSYmjsiU88PsIiFemiv74psJZ7o7ECUH6VA55nEjw7Xf1feLeAkpxoYnGbz6l7hwNqzPVSP8ZQI
XmHTdcdgOSqfRCH/s/K+dmaIpnIC0X1hHqM7Sx3mmyGBG8NXcleXypjepV+i1q5h8u/1Cj05UEaZ
SH6m6FOvA4jnQFyhH1xxuynTGBxSuK95zQYxxqOukKF/cPS7fFmT3rt5ULU0EJ39h4xqXUhJ9sIF
G8OEgdkOtWtLw1GUJVGQob1OGOsKPmjHqVUboi2J/twutLQzI7P3y3OWiJ9u+Z7AKt1iHrTkhVK2
wcmhGPp3QZMW7MSmOONYhzutccVb8Ezwl2Nmr7H3/Qf4Y3te71UK480p1ZRFzCNQqeY3BX5n38c6
hAnpWj7qQgzjBhrGdTaru3mLrUURlSoe+QZURVGt7eNzsltLpLcGCr22kWmRBnpyQH3D3HtBhPBG
N1FGITOhz95vMVQi9XAoWnlaPwFr65h+itl08B1lDo0opi8ecVSyO3pnAOqOWlwpnT/ziNxq0LCT
6o6L0OyWLxoiTPHmyRdxaZX7vmKrIOYtvKy7KJcnIFpRohsbF3E6G6fSN5hHeO+5oeXG1ib8Yl8K
RGWV8puAW5DXXNA77RAtjGiGgT1zuQT71Vt97F1EKwxzCB3AjC1kp7bWhZFLbGx2ovTjjYQ8ZUQh
eYeYyOJSAifaZwXcgmN8JeIF2zJOkrR5b+yA5U9nWicPHFLX+HBLQz5oJbstmIdiCisoOm9a9ytP
fx/D7TukSmeMa3XeOzq2qYvVPQ8/HMrfAMS+0IABy4nHcB42djw83iO+p30GxKCYAc2S5+O82c56
RwLpOeUOdUByz/1KgAr1zZiFmmg+YINyaHEul/ka8jMUiH81yoFmW2IbmrStZGZADgb4AlS/6MYc
jiI8vH7D+Lcsq+1g8tT3HK8eP8pAAKg6uqN4/2froxbN17h7qMCRs3Q5DEdBGheQZlt4Zzv8H+Hz
OYnr8m1Tufaf3H0Y6xpHPoubJKnS3wyRmcpITjGauGXBqo6n1h7C8XNj0U7Xh0Kb/Ap3om3lhgu0
5zVjOOjFBhzG3fvl9ALZFORVz9X7Vr/A/qUbjgsHpxM2fyo243i0yu2G031fguGT2xi8vR0cqpTI
tcfbE59wKuDlqloFgf5GvTPyyKOnjyuYYTUZS75UlbU9EkAF7FZmx3lxepIAt0GaSr34gl/QhN2d
KpkF9T3/XMQGJM3Aqpb+R3b0n8kWKkt98/XBdlpmqh9fmf/LTQq0Sai5ppyVP20A0om6GA7VaKON
uOPgs5tAg8YFJ6JcDF96g9Qb0iObowSYx2wgTpv+lSLnKKi5JKyRiLavQWTPphFWOSUyB9h0l1v1
jAZEwCuZvLbR+A2t26eCniqADGIPZYZIn7bnhyHHgm2vcD2Bheceiq8PxlvUWvIYlu4uYh+5Fvjf
H6d+cpyB44dE6OGLLxlc2P4ruOmogmbVc52UFXs5yuT59iONfd96BaV7vYvWOauHM28GT++JjJrt
XE09AamEXLDMKKP8oBhRRi2f/pCJXIex8ujTKCRBla0B2TouU3d0mNf/mDzYvpFHfyxyjvseyBuV
H2FG21xf7HZ7sHpzQab94PsXvE+OyhXWjGYqdufIgYCXm8COrGbLFA/aRSukWcx+XgWfgLKOqNcb
Jpud3+t34+oBsa0MWxHzsOE7WkzKIvIwqxSUodkwzfTGrOXn45JV5fjfkENOffZo3T1lOciyvXcP
xQf796ecgUdClvGslA7pqgv+RqmUp31SbEDd8Nvgr/Y3nvEZJI9xpaSm9N92iw9C4LDn+6PnOOyG
dUJzIl4fgWvozJgVUpBCgMR8NYeoye3i+0spEP6JW2AheGVE+PEcvTGrW7EH1bpKAUz/d3dRmBJO
1Lp+8m3T85p5GQ/bPnTjpypYMT6/GGEa+eDDZvz+zbfwIATH9r8CET78rGW+RabALJ0EV+wMBkIk
eORD//psixcVCxYyh3Xp3EsLR4ik7tONZa8bShUXp/7mEi+ceXd/+4K6+5FZN5SLKUFU1v513d0y
Ng7ygNOoPOp1dNy9N1ptZZRjFt6sxb/wWpp5QFF+ooeeVtDcAlNv6ptAL4sT9QsP+wzYpLHDXVL0
ErUQ1lYmJR7b5V/8LF3fRxOXnHLQMWPIeVcnNAS04peBSzN5bOf1I78FtlPVoiRkK2hY5PpX5DKx
8EhRI2vRPV63SE843Jv/GuyP5nKzMc2KPVz37i9qrvL6goOpC9j7mToCfE12Bfg/m2fuFm2qlAnu
WlM2IK4rWc1Z83gka2KS70dDyd+d2i8xJAwOYLIMZt9igrOCak4r+inAwTx0YqkNjRIRk0S5oWKt
OZ76I3f1PjURwMsj6EWzhmVWdiQUR1iFe2hiHbpPm6tiPhKJOsauYkb04TPBZjLu8KeBWvMgRsL4
ytZUANWguA/5aiZeO4cM5VnIX9FBqS7O2Pi9Q+hHIIp6tFL3Zy5r2cVqW4cSDeC6aq0VLvinRanJ
rE0p8z7S6oUTxlg+tIgASS19Uk3NBCRkxE/Zu+yzDL6ZhiZ53dwAQkNIR73FOSElax0eBdJ3M1fg
QpN2VHmBIxLJW9OBXkVIGkf1XCV2nVKfiy/HNH04vm11P0c/ZBfjiqzoa+Obe03Pb5+QYYevj50j
8m9FtKibEleuq3UO3J7lFk4TTOeJss1KKBicgDfiA0MjFY4fc1hYwRxHg2zjZbahC8TwszhYhKOC
iN65w/dQKv2/si+ELNQckctoWjVOD9jPjN4K5Z09ZPwzAY5pGBvePBAB+wYOzgbDs0xPVa7oY6tV
AreGdaOK93JD2Y8TDNUzMferytYjDVTvYfnh8xtuSPjhUjoA7o2S8CzyXUOoacBWCmikAr6nv9sV
crNDiOVCMrJaV2G/PmVgJCDtSAyTt181hIjF6Kdi+DE8roNgNP70C7ceu/VJ0QJssYrGZMBh2t9Q
R7pqeaOeFMKRHUsjFcnYayc6KuTpEsn1WTDFC1pcLm+YosynKNhleB29lwwduRAnOuRRdTTV9NAw
6/miBmSc70lY8/h5klVI0Fr11S1k17jtt5S3UmC004OReUhsd7VGxJzWINspfWOF7tiGOlwhQKFt
XmvrdO4In1rffnyYWYhobB//AogFiX6M1ML6DqEDDDYfdBf0jT2R+8cJxFhAmpc6L1wPQu3kgU8c
JW2mhcneb/upxnbxQK4mdqjwgpEXFs8lLN2XHR4+XBnwVK9UZx1nQz2JQjzP0Zou7DhK92NrHdi6
qkWCHlUwWjgAOBG9NaIKhWaDGMsuzNfGZ9iZKPdEte9EBcEevss5+EKs1y298NtNMU965gyJfsO3
phKVU2JAjArXb5fv3s+qi/XSID3oJPAWcmFncnR5JzdBIWA6vcxT6YB+Mzwe3NOJQxTsBO1zHQTH
rw5FfHQ6wvUqZND2MDBBUFUPkxcsWy7Mf2w/1eIXhPGBW1T5kJtuK4ignI8P8i/peLD/U8BljJxR
n9KMOIg6HP4sgKuVbzDerZyOt4qUsVGI1HW4rQOyDSjGDWII1S+fuQ5lI0FpJ2t3xGMk2aGLeH14
PXlMHhcZ0uw6T8JZl6dNGBEhFrvwo8S+9ppdsh3ZCJ6NAEwVqBhGTthcY4yRYjnRrlanK+BhIsHL
kl0ZFYjM3Hl4JpZjxKIMu2J0Xo9W7Z1kCITX9JEi75xLkYFZFkWjEJ1ExLc4KLlS9rwJSHinFKUv
h9FTvfR/WspstvAV32dIzvmqW/dvnAQEbS8aPgzXTy60Mtr7azO1p8Xk7uHSEKST+Siu8IHWx5r4
UTHODcUjEtdad0FrURL/e3DQhPNjFSPQ6Kg6JuE4C4MvbTlrvF6MmZBm3OgWfBE51uMO6NI406D7
tLATTmyA7aSro+HPjwf5kY8buX8R/vzrCWulCFb8wIb0jBewQbNp/zECkG9Odnm79he217lFKR5D
0aDx7Sgs5zNLggqsjYpMxtBP7TQYz7dOfj1p10NN07/VmvwAGcz8NMTcppxsiXN5IR523oSSB+c6
iX9nnLf33d7h6sW59oRqGO1DTo2RMYU6A9Elo3jP7f5o5kId5aMflXriBQcbdHbGtnwui1MCvXgE
ze92t3YodxKrXUVUhyBggOjNPTo/mh7yMtxhH1fuuPWJAXMcYxyi2ULULEfeRzhD63DGB7kag/aX
4+8SW1bHbD9ys3VDbag6GAPeXV2B7M5G9bRQW4plZHX8tfYsDpRTlIRV3mbgg4hy6nPiwvU/i4nM
IGRjzC0BXHef/Y/ILunsqKPjYe7kTtZGRA4B7BiHV1DIUByCfwnbSUlyy5aBJ4xPmrKxEDYHVyQk
mCjqT04eknEo878oXbh/L9YkWmbxn4QBoStX7ApBBC+7LnkupcE6fr8nC6OzDGyKbjMXWvNZ0lkF
BSRlXq4nMEmxHNFiF/16Dz/kBKCvbVUuNDqO86g6D5BatQMsCtjrgZdM28rfcZ/pteqchHZ2TAWC
HdJUax/x77DkLD6+UrB9SrClQChG4J71lsQkzHYVWYRKU1evjQ5lHScFMfR9s3XX7rIPTwSbWLYd
iGKUzA5BSiolkIcpDaC4NXUjJL6vD6Zai1Wr7tGcUV8ASOO+7/VpAvzgIjdVLui+C/L0XaiZYvg3
Bl+8ikXT4gYftBczf+jsL3c0eLuYEIbM7uiOhhgC7taIQvRxfsdXr53BJfStLa5oAvVsAmWVc8jH
plZUgoNBxDsX8/vUKBI+C8K6jlc9MAKtMjLSLaAE7i6Sl1MIZOdomClUVLS6jwGRZqDlHwbz5GpJ
jSLbfpCa0ZerJxA4guYyCss8QlDEqwG3PpOCriE5e04Zx/ilp63Lf9ijSIBl8aw9RWPnx6S3gvqd
OZiVheADvQCXFBCb3DeRKlVtgL/i9Ml8ZLSd6XoQbdo0LAuyYuMRYBuM5m7zQAsr6LsXt7U9BgPZ
F+Uc7BZlM69adT+wz67HbJIRAW53GPT0exaumKkcNvtZU1F5aI2hMNymYoPGDH7DRS/yguWYu5Oe
SiaaHz1kgIxvz+opVlg6Z5dr/2H4xirkH9dxPH0DpWDK9yYsqwKsc72KvWT210YZvU6AMzSHrzZm
slIIL5oVoNl4fEVSfwQetkVoT12YRbqc+NvobP7ZVZ2GLE1lJKP/B9e30/qg9GfvCtmRWVRt1aaP
KnrX/u3rFvD1IPf0ZYxq45AVOPpDiaVb4haZtZA0qJr1tL3K9kJ/be3n1Y+NJvjWAOQ+Ny6S1+QF
1INut2cmKPoV9ImM47p7ApoL+WKoK1uZVeyiP2dvV+LlBuTmgXx3Qnq804h/hXed6Nhm9BYstE1K
+q1+JBXqPpr0cyYrhFmbVFDAV14c2JD2O26kKTiQebSPKGhEjveL1vlts7FeCMmmITB/+ngBYPhO
nL5xP4Rf5tn64U3/v7phSdCwl4AXO8Rp325fbLP2VjP7HRQmR6vy75wYpn1JK9h3mPRlLF0cGqIA
JUG/RInHn8bOHuHUVw6cj4ZpofUyx2G3Yf3c5rQTezj7+/0ejP2zhDoG8pglmh/FvZveb9Nk+bdd
g1QB+s8+eslrjz8R933B+dv34NHJkt9vtpcyGhJ5Cn81NfG+uNGfEgiW51soS64SftM5k3og4bNn
DUUz/Uv76EKYxU682rZyVkzW1lOU35rXz+JSCkY/sN970Y2RT3FugtzzGKgwRxaujEEsc5B2QqCV
2SvYza+DWh6emOP9tB9lENiQtMTxM6rBQI2zpaQihYzin6h1HWS8ZNR3u2c0d4/G1WJbtCeY1eo/
HASRKQ6QfklcddJ/evtC9mNxDgYEPdinNW0RZW/t1yRyfVfpvBDrdamIfSXRbRWaY3neyCqdBXvL
CSuzoPAKppWIWIFhu+omq6f992mjLRYpSFrnZ4W2HOwfmDav8CPMZF751g6Y3SEHE3whpDtvKYkV
wpJLOv3Id7iJT54c6ccTTgyAJ0YAOKIWhhbzOaTDMEeEKRWnSWJ+y5ikLg3ICiXjO2VI2VutdWiI
2k/QUMnq/LXhTtg4Dp7v+OEhSyWxmXVgEGlVUOLso/fnIaKNddndcdQiViEf0JVhKeh4SwmBuXDC
lHu+WpYBZxDOSX7v1xMqOFRLVauyR8QH6hTBRyyeTBl+t4nkZ0hATp05YV1SJzGRyXiuWpwMkdcZ
uR6PXflAJByYXjPTZfoyi6QdAqkv18AsPc9ezAxtDe3T3ptUZi7CkXYvU8dVlr3I553Cp+gHBjGu
pr9eF7kVDyFnF5WZcR3uMmziKszkjAtnPTYJnMi2kmXMDlsHzn1nH6msIeDoF6moJkrCQyQHo84u
W5lNTXc1lgzdUn6bDiif2BudaIe5oMwjFS3wZl66il/sb/9XQj3qmFYrbNFvXG9/5MFp5iC/EmNb
/EluiOQIQm7HjuUCl4SVAfdrVNc3A/NC4yRcsi4lOKqX9DYLSDtB72cxeu7NsHvbXT08MxXwwvb8
Mafi9BFvAGk4yPEHtGkXLWRPDt9C8qNrkxLx+OIPPBss3ngkvN9rgJEHbwckXRSEpm5VTZ+PvWP/
Yh3hFnCXEQX1CZ7MywhRailfdKe12h/0NRXl/+ZCgaBCoz2wiguV4UTAT3qMBuONxBV1rOX7nnV0
OlEMmtCmn+1cDRfPk/OSNv1RQdJW8l7GLbcrula1bnjL1QDTcvrXoY1AkN59f2+xkT+7ivC7XEB6
fkv1ORhrbazNRosyOHvzWKQnZtNZylkPv4ajIhzNYb6DXKP6jhvHqie76rtmVbhKsz5iATNYHvBn
Wtl9+uPF54+t9SyLYzJgLJvQCN0ZoUsYrW6uC8x45RzZYuvQWsLwlE6P8PSVR7ijP0sOifTQ5Xco
wY14mGfr5SWcfR0YrWlAFJGPh4STlOxwix2NQjTb9rF3i2UXUly9wtS1ziSwe2yHQnt0LKDxioJN
JFF3d++Bo1E4dOf9mFMtyiclP1tYIlMYAiePDOpGFkNyYhQlw9MbOBbUJ8OJcCB8JynUQIKg/oAQ
4IDyNW8RhVW13Vi8p5MtZFcB1of+LseIY9l3AHpx7iAKNziIZ4tA6U/oNp3L2KP2gfriG3erujWH
TANo1SsI+L9f5oQARj3aS8FJWJ+xykqa2r0lM6dr6iX79mEiJJPNkxlW2eoQw8wbNsad0UK0uL33
dJdl2MT8FyoCzsVWucJXLHpsTWSxey27NsRjH1GE8AqdXq+P8gNRbVEGZvZnPTkgMGtfzx83jFyJ
X8hp6+9uw4gfHeSD00JUMeXSPGrOxOTzsw5kR107p4rv2NPt89Bf5yX9+bnsnvRhgYmj1j95OQS8
9YTXt9tKzKKcEF9AwakWaSZQury4rosEg/KpALIx43KwTAjcSHoV8ip9GJ8+V+/bP1kp92ot/s6Q
fQDFqqwEallbG7Ppbn1yzBQlqp+SH+/Yx0Yien5mgfSxwbt1PMBtdIQd/NOAW7fazeiwwaWphMSZ
6m6K89KhlkazVMEu1PYTWh59r+Ydz7NE3ptf/f7+cHZdyp85tUN8dbU/KE68Jzo2vL8nmMlkihWT
ibbc7QP6EhTI8vklR335QThMUuZLiw5xl1cbPuVITJftv4AMyN9f2OpxRHay19wlrvh8nHF8dA+F
smcVyD/MCy3nmBk9WkOO6ASEBCHB1s4GicfY8hlisA6T2pl9aXf5q16nUT18T8RnzYV2nysx/9+z
1YU2GKJlXaD9k9iFCdy0vmb7qQ7OlzvPCIrhXlyHbpWihsRWVj2c44HX9TGi2V+IGY6H2aXXuzkn
JLoNZsIEYqXNBQB9pxD93pu9w10zDV474R3TZVC60td7EHmEhweUrXaJr/zg45lvGpsuz4RZ/N0R
KzFYSt7QK46ob28N0V0hI6I3NrX3qzP7l1/1gu9dZ5by+fNurWERGKSAoE4AURcZ1e26heuEOI9C
E0ZEy5Vtm+JGrNbeRzz1M3r4zYK+SFJeY8m/x6fbDl8lVnpuQ4uX/TQe8h0uquPI4HB+fPEcVzln
fjitytq+cDj8vCl2giM8lIsBkqtN7M0VITFIvXACzmyqrbn9kYIwcD0pLDspuOiiJwQr+IZK08li
uYqS9Zc7lvnkJYwgiPBVp9VvVb8VL+6N2DZ5mDAlyq1ZA/KZRlu/BRPaOFOEi7oXnEDYZQNeSSOh
T42TPuhdhl8rh2wQ12I63McGXgRKbqn27pk0pF8VH4rSCIPsXbS3ppOFnaEFDREutuDVzrRtQnfZ
SnfryzEAEfjUT4bThX/1W1eRnXfGuFdqXw1z51d3MOyAIig+oDcPnm9qNLrmgUN0YM+dQ9xA2qnv
KszyuULJIgVJk4tb9Ijni7vb3llOZGjzJ2QVq2pdD0mRSBWkKCAPJEkxqeTF0eUc0MpZcytTmulv
M2YXgQodLbyus8ttC2oDrWcI7yZmI3Si4HKoBA4hqf3OwZpwc18T6HMrlTMNpuovrUWGnPLTNbar
PPW/c3yCuSRpvMeIM4nDAV02H/dLb7E3OWfsHU8abtMmqZXT39wlfJjqdOGws5xoJnkPvbqXdrVh
/l9FOSLnBVF+6NFLUf7vFEM87j0LxtKoh2v6hqyFeeQWZZBG1A9BLfPIi9skG3CwEepJrwAVYZ5c
eai1Unto4091zsHvDt5+4NsZSTBGK4ib/JoZFfd/JP3R5gBWgS3fk/FJ+W3y/LfK/4pLMmsDWnC0
ijRXCJobMw56yOLq0zYfdRbklZIGp5Yo9Gfpm6r1TsQofGMFRbe+Qk8pUSQbUxWQuLxXNTMWX2tR
p4SrU7KFN8WsQnD30kY9wR9NwbSA2oecnP1wPjF3cYzrsvI7Kr0Knx0RGtyv8SDb64rYq2VH9/8O
Bky704iw5J24DQBC045cV1jpDToz9fGbXyy8iadJMVENFlc26eFhxWL58Npr7/0qe6kDVjuEHRBX
kRjrjUg1UxQFmLxqc2G41ldvWPs3rWdmsq3pr+ibZCiLPQT2qznplwvjSB/hu63PP6ABfebo/h79
srKeh/kVxSWIdr+PlgvVVkwnfxjUfRrd5946nzLg45NjPlkOhY9F84P5GbAKskC5G1UkJel7TgDT
oi3RlR6KKmXM2bW4KYhEKZ8Af+hHiso9nEfgz8pd/ncp+2FDfPulAV2msEmnIm0AzzjV5RPH05+M
KTKZ2G9rEe2/cc/ik5emnnW1x2Ebecwpqit/qv2uF9DOEKmPRyuYLD7UaN1OhtgqmPSy/6tRuIiZ
BaZ2huxvhs+Urj1x4jeRcakqvqWSVEAH6fMzvX4OIIFOqaYmHgxMMXtRoXjyvUzZrBAdP0vXH9IG
SPO5oL5Q/sIWiR4whAmlZZBiOmQ6142vFzkLgYvWeX6awDnzdaEFJUcuVsXRdH8l35JAUFGbn0ep
8Fm9UKIkzPvaUN5ODhiy/B4IsxyZwvZc4BNQ1k2fyO1LpFigwO7gFCdEqU1f3lAU4PLtnrywjTw7
HqASKiTn//eQvaWxX/pN3vYIkyuP+W8rUsw0Nj7p1tHl1bq/osW00LHYgkwfdyTCNTKPaLyAupn/
+87TnoEyDKOxkkFIsoURqsjcyXSUpLf0ZKdey+R5j0vyf3Rzx68vDZTXYsukJg2qa+2xOWK9l+Ez
Y2G1u936QKv9kpFMXw+eAm6yeJHFMOhCJR0gfkjsNX3NTCZaxZAe4dolRBwNuL016bgpaSrMoAxz
sCMjYX7mG0PSugVRwm+GbErV4hBqo2cRlyFavFDVQyROukJFcl3BIV8QUC6GClhqN2aOFaSYZDVa
6FjFNdd1fPTdyu9JEbmU4143eFKDpCGEmPttxXRPFw7RyKdGhg5XV1dnj/+PnJJ6DSEWu3at3bkQ
c+WOPK8+2q0v2QRvsjo4h4SMUmffcZ8d7DCjAlXbRwRVinrtroLNLvGpT4Eb+FQpv2F7R99U1RYI
PRhVLT/W9ZyNKY49F6cI485T928nzpk3Ps7ScUQLRbyceRMpIKnc1nArZEI19qj6Y2M+s18iAyBX
+nm2QEwmnrvZHYyzUDQ68iwkzyKhwYuyfvNOWvZ2rP0VcBlLRorhNGkpBoZfqWfLhU8SDDaZ08P9
j2ewsrrsTaQM98ZoWF7ml2d36y68CkZVUV2N/JQzF2GWYzOexuVhGrdVz9r64rCZWOaL3G4UrCpv
EWdZmW5yGjrYGSJi7Q0R+8pu5NvmfxM3E4dVSV+638LnBDIqlgGIhIzC9AGzB9k/NZKHJvVratw6
MeACVXnh2k7+RPNDulK0u5XeRHPFpPwCAjJ9FippJC6ihOGrj4aWfnDGi9vH20KUjfsbG6Qo24IL
BmzUVw/FHubEUerkPGbKv4Ycmo0N8HbXSjCEWkgBZCUda8QfGGNPZ2nOqrOeXkb1KZRGDpWeHkOH
06QqDQajEtltY4aF3faVCl8SFkNHz62779B9BFuiaxY4kKGJzK2z6IIiiVG85AFivg6dkZ1ic3jB
cyq98lpfetGa9MsoQXTRT0fHlimn+41+BolQEE8BvewkMYchXE/UoKIZJ3TTO/PJGixeIRXLXpBo
jvhHhCfKL0y5rSmppUcu/6hKolNHUuiOMRuk/eQoWzBjewRZWTbNOEhYDoFhAgQttfAl0Hl/peJ6
Xe7l0jZ1uMOwFFqofh5WpVnwsy1f6qi36O/5yXljHrBCbvgGW+fncxB38NDzNRFHP376o1FKwJZI
dyJkSZvuYlBUG79tR3BpRFnNLtTKfrTw5UGY4YdAJRCmdyaYFhUE/Z2dcE83VofWbDL5jTGbFL5B
k1y/I1yzj3D9a6K+9gMr1KGbQOrajQs9igqWPVcQntRmHkiw3H3ylZPBKuQmr1CZa7dZMdwA35Yp
L69XHkrBve1as4pt3FvPMtRUr0SVsYQBnNIZgXCG6IsbTKhE8Rx3oNU1VMuEmkW61SnQZigUYAbA
ex0/PMHGhG5KHaJD9Q433J8IR1iNaa+ozozy3566cPIhPQOxAGUlUTYvHFcVU+wrnWWcLlAnS/0q
t67gwNYzGlWvzV7+GG3BC8WFObUPZ0EHwPXllMQezGt6+jkjRIfgWKiBFIStmacFw/y/kkH96plJ
oC1ZbAS/Av/iKhNRLRVpjgwVqb4NrbRPQKcVPJtx52INMCiZPQflG4c9io1TnB/00p1FHyLXoMvC
h5hOAygQ+J8zjFRz98H8AGLgMTUTMitr83PDqz90rGwmddmDcTU2+BpIBL4R1PD1xxvGTxzIbqH7
xVt6iO6xWbB84/vFSUhHPqOJsUvE1Hn+J1Uck8Jg6PUh6K8ECUJ6o39dJUC7r6EtwNkNG7Smb3jn
iaaeJrp/98qD13R0aH5HN2wxWDSxsLNfQNdPOXg7sEkYHJYgl2Bsz048qKiRXVUbu9nGlgBXZ+nC
SApYz9/q9KgPh/n5UUOoTnWAzf1zFFdLSD8m9zCfiqnf2HXHxupvUWafwJrjyRyX4Cbvuzx6f35s
1u9nzkiJfcNZsTsPkuakES6b4KRs3NoP0zvZtCoj1yOhKDSuKMkRhpAkeaJV+m5R6fL7GDXbb6Vn
DHAXukQ+Q2yRUO+eEEucuZYaPO+LipZVqAdzvK7yh7H56AGqMg0uM3DrPaRXZ5u0L1sNRcP3KR+z
1HDUnbPmtUxbgoChKa8GxnvxMF16MY4xgYJr7X9LLiDwYN7MX8rMktMoTezFzkDX31WvHEEmRBno
vby9fIUNDSYpoGa2rQVxoxVJTfDk4JuU4xQ0wKyuR8E/pf5xRWOWrbKU0MAv/Y2paL6vD1FN/vxl
Hnlo9alm54vPDbnNx2JyjqUy588SnepAH57XGUEXU6qUUR2D9mc3FZQJUCvCWgC1UA3nVj3wF+S7
oc9SbFO1gdevF5RgdvjBJHD7jZYBJ80ZUUvBknX111Plxyu8MBqGd0coVUjDenoumkWIO4MC/tC9
PFe1Dm4OZlR5yoezLPp2aJE13T0a8C85s5kH1YkjxYNLpPK7Ts0/VZGMNAZ6lYe/uRVvy7XizETc
U0A/eGRgG72mFLdm4zruNYwWpuMf5sO8vRR071vDsZTLVSQND85YhgkRSkykwWnBeR66na4ZIcWr
Rabx0R1+KGCw3nOlf246llRlhpcADf+T6gE/hxwFfgsZgc0l2NFt9exD7nUt/ry+aYHvFL7hPetG
d+/oS7vykAs4ZmGnK+J/Ecr9PTq+Ob+vhzLMF83De7ZIyhB/lY860PTz+nJ7CfW/MCKoKQ1NUQYk
1FhKdepJzIRf2f30VUdYI+QyH+bLFTUB2oEc5vNns4i/iUHjnfrIJK8UomXYfbaHpHefzUnTLGSO
uXW6Wnp9j2R7QsHJuBlLD46rOzncGcJmh95icYGM5Yh/sCTeyx4u0EPcYq/XSDHtqEVOcd6ifiNu
LdyljssryyFpZOYHa1r2hRnoDTMEaV0n2VDDaGUEc56EzWQpcFNNeoVUAlv+91vRprC1wtfEe6Bf
XgbLfDYJrIT86juRoWRR4YkI7lnklTIeNXt5ByNBmqdoW7+ulhdK/ygN9AtZbkFoOMwE4ZsHC3UL
um97IHiIC/pdJtM9at7XbxzycG+V/o3YDmSOCP4aXFojRy9+V7/wDVn/bCjIPRtcMclRqWwNSJTI
CMBSiUPJnlyiq9WtNLDv0VurDei5jrJdOUkG0fK0VMZ5qz6zkdsNcmEP+wDHhMm1eBtqrKEv8e97
pIDTIiau42yUmHh7Jvit+4kQDOgWPQWH3RthaVU5eThIp5bBcM7zEl69lFLMKB0MUFN6b6srvDWB
AFeKNVWpBFWzzeLNt8ZjHa7D+ikWn7yBYUKgSILWQYPKdEUt/mTK9GWNv9UfaQYOqJ2gAU+APC/K
F1nztdzRR7/yB85Lzpy2NmU8WGSrv5MrN7oOlGF5j49YBxvjozAWuJEUIt9agyeVkzideFjy2isD
9MyU7U/hshzdfJGER/fdwHfrmc9IUW8biXYe2sCZ/qoH/RGxMzYgRVrZzwUH12H8n4Uavk0xTIpC
aUGBahlE/31nh7Li41843ZZ43Hrces1QzdicL4UCjBCAMllo2jTSpN5QWSEtpZeMnGixVggaTf5i
pJ8HIvUsEDuosPr98vJU5H9RoJSuIyCN3uL09ulii7Y1Q2oyV6biS8Y1KMHBQ4sP3/nWIvkO1/xJ
4vwE15KSkGfKT8pmQjIPenW/m6gU9rTKxC8D42N5kwbibcDYXcvOqD17sDzpw4YTFnrvZbApJrEq
obPasyQyotkH2veQrUPhWeIsH0Kxvzpz5WpZNzClP4aH4i5VmbhvRHT7BLkXRLoW8Vko2IFsjZ9G
sUwew9q0ahWjUs29mGoBZbTbIIz2g5F52QRcLSXZF5PSLLQcwncK7B7o29TKZgynDb4S75hpZIkY
zxAjDEecp/7pejBEErSxr+GE+B2Rx4hmO9lfPMKLsHsDwEuKo9ZrbZSo1/aPsOnfkPyYbcQ+bqZl
ip7qxq1cysy0do+l/pm7pFM9XrYvvGuYrqzD/qnp2nCKIlByk9fbu6C7MtAk4n/xSd2BnVRJQz/3
fyuowngm5m1g+/bnZ5q6hxmfbkfueSrSgMUtoSoyzIoNFVwUh/dMB5kzw6XqfsHicW4N12W/S3dQ
7VAcd6bhTyrWeANX+Ld53H3vzBz07AGssVbnpgVtH+eLwv1zA405GAsFbbqpaEJCm/0cQ1zsk6fp
HV/HBYHrh8+oNg9AQqQE6gXpk81vIwuwNH3/0sqVCRscL44qI0PKbhW7iM2vac9a31nvcZ3mCGrM
WL0pmIOi0aReJuvEkOsGopkbmODFwL7ntPyRTWDAQaIqvfN64w1iPy0LA2zB6RwmnsmT4dj3C4/X
ZBAZjG8JB/AZjG3kzDez3v/Y1AphvUK/wwLX+R2WOCMeyyRJTGQBdinzq/VbZSxEKUWnPHCFDXXC
+u9NJV8H76gVP36NhDo7qDgQe602vNckH+NIXmXwVP3pIIY+kOeLIONN59ehDLnxnyRszC7bxK+c
s9uTP6Wkc2fxPLWLTJ2+sVUu7CgfhDT3l6FmGLejdGVwg1iywkBKpJ9ubdCiW4lU7S/dVwIUjNa3
nCGPVYjMxltYle/nky8fkTuRkaTFmeqqeXyTLvD+OZsRPkCMJMcDOdIPeP1gUYgGDfv9CMDjp3nz
8VIvvPK4WgJ5M+9oBBCNnxkv7nspVSEufOk+oxkCFbc3CFgeoIvorpD1YA5IQRSGXlc7uXnTbCn2
XlrEzs0w9g4t2rxbm2yP2Gauze/B/2UiBqFjlFudETj22MtDRc3aleh1pfhyWXq9ry5ngSO6zQqj
U4QtWXbVLMeS5n5GyjktMRWYdbK5niVm6TtSx2tZBPLVoEFC1ogzEJlKG+ciBewj847vp/Igj5JT
PYVVkNN6UUBDnWSahWLM+koqKs4Bb6n9tPKbLPl3vJlml+DDmlOHRuie62i+ACOtGnNq6PYGFsVA
mrP4FnnAdNeTAswossGicAwCeC7AeLDirHrRbGsxMyt40V7M7ZrpqSvbvVBBcuSD4kW6UkDqjAxy
zRJ+Y4fV/bB3ZI9F9CKriFNop+ABch+UVUl3CgCntiCPBCqfin2k/XLriwAfMR8M8cAvb22hK1EE
LUqGS7fvuhIr3AX1GNhE5bYxJ2CzeghoMwZNPc5pTetp8NYWRGQrOU9CJ0lusgGIT6rTQN/16QJT
7YxCB7dDHCHVw02jSwrdljR+juyjKO2bWdatOGVAE480y4vVGNhdRoRBCr44Zd+XN7BxoKFheAG0
Nmv6+9WSmgrjbB/4xfVQiZkuCgNAjcW6BrkEi2TPjl8Gu4pdaedPhBnOy7BgH5H2IvRoMD7GXH30
OpsGD5zutnUypTPficd2rZOAY6xKIB9TONrDXWjOrq51brDzBMO8YH9qPRWXaYi/FyZE2t6tnzLp
TyN1mslFzGEyRN346d7QK2NJxKbM4QGueVkP3GKKQPbvRFDiUtf6cGAnsbOsKX6T2tg4ZIaY/Qdy
YFiWns/2GOORsErW4PyO7Aq3tqBOzeqF7MJBnhuvspQGAsnu+1shuW+U7oSdNJ8jm4r9j1pZC7W1
6hnlZWOjoQGyvOCfq7KjYbLxPfAuxGUdHLTk84EISEOKmsJu9xJQM+UnHdqSj73wktTbRn6q3y/5
8BoMWnpNiQzaHR0cR/KvL18UG1Bel9wsOR0B0miZF0a7C3hYQMdB3JwlDeizlcfE70poT7gDbwIh
d7viDvpa0BlCKZWYKUMI+zuC75ivzUSx5jouyhcXhZo0Mje5eICmeJHW+1JYQAHcY2JGD8JSIb/a
yHkzQCwfQPNYxi+pgFcYD5N6apbRPOMIgPaRykEs76SAxeBwBTgJ1lA2ObmVZykzpZY/c+Dg1qzb
lHLOYRxXqaN+XTabix7w5lz5DywDmvAXt/vSsMJPYlg4s3/eN+X+rsgaHpSbK7v7O+zbAlu0GDtd
AwoTfn+o36V40S8Oz4oaj6Jef2FZFnG0yIWLIRn7HU71oeyiIFh0cBNWbBQZpjB+iEcCCaorsKcO
AV21lnb4aEI5k/KfMphutyy9h+qBlFBgqaabW+caZ7txjwUr5lfonBgRla4PPi+DzkLWlYLzb/3N
x/SwUW7LgIahjxZDYcbNINOUhXWG5y+V42O1AE9JOEsRT9FdM4N02FNyiykWuDRytkn2Ora6TnrS
+z9eaTCwGOVjiyc18Uqy3lAsYYNe3GKrFolL2a3tfoG/9fWK/TRk10fRkE3QcDnI25Z9AVYWo2DM
niv1RfCBC+LS6hCG5ORJBvCS3lFZ/jrkkDXZ8DynaDslN9otpwIUy7lPYMF/nIec+RGAi/wypFHj
yIgdJ7BG/BfMIuUXl85P4PtZjytK1w0hXKDwSDgHWN8Cy7tdTIts3oEr/na1t3yrGrs/8vwe9tlB
nKRYCPnJWjZIX+Tg+fV08TkC4u+aaSejLSzNZIp6wk2dgeDkYmwFkuzdKtM7/cEzt3fUb4z+7HMu
6Wv1dh6bVRotxqw9BCEkNcqO6o1B+TekjQ/E/Tz81tfgQ81uMYwmPVXQu9dPRgh/j7riUE8Q6VC0
0QhoVGJYTCOJc15ZEW75ITA+FOzAaur4vLPg37odVaM8m1TFapMpmTRMffihGW8ps5s9E6uwasb0
EuWcLiIUToPEePZZ/dBtNqYTqFEwm1YzSG2kPy2nmfXuR3XRR861Y5jdkLPG4uBx4Pn6YxCV4yWs
29O+0ChbTXZcUTrEHtGJsKNuC+aRjOxEnLdawSAi5mB6+F6xgMSP6fTPusKRyxC+zYgEamjhYzUH
Se905XqqXA1G/EKD3A/J0E0afFAtVNHs8As+HZMFhERRtHfaGrP+O7zj0HXfK1NoepmfiQ7TsC/S
jN01f5xhibkNdjEoK0q08K5CCKMPzN2K69GWLQh8xQ9i7gkjb5Y62lwmEz9Q2wMdFuUaU8sIuAR7
cMG5n8DooeT+tnG2D5LlbiFhXT/LycfFg4lnsJ7l+BT5FjY62BNgGdGeBfrav4ZVmD/ZGi3/eWnU
hKASLFFef0Ot6WjiRCTKn6KK/LaOsAsihYAQCjbRtH6w/SpPuFfLa1mCBcIJ9kkR3MrV2WnaIwkR
FAlBgbK0F3+oGlencNk/Qfx1bQKf8uoaYWP4tYjNI2CKFtgO8aTO9v3wnwZtJsqsuUgNC50tfp/z
42589gYWaLFkcIA+/8Xz9hq5E6b+lY5IvooEwFzfMDFjEfalDE6y2h0bbEfms2GLl1XZ4urVjitH
jqpiqKd5mrMgRmVHVAiY/e6Se7wAnwH51n5D+uWpJJi3L0mZjOdtZWb28ykiKbqyckztmjh/3yLD
0clw/o/PxIWeqYBs3AICitETUM9m7AR3FMQMzgD1ILBBTtPvLexTgXtmd+61PUEr+3PsAh491xht
UtkHLHXF4aE1TNwE4gfG18tqV9IZnqMwIcn2q8YyQdMKUSJ1ZETTaFSt1iiTnv5M/Ri7ya0MqBOj
4damdREPepqj2MWtMw4idN8/bBSHOqa7husgMvMLpsE1fqVUWn/JW9qdhr2iI4TbpH8Mlt14/xoo
x/YO58K4zA7+VsvBqRAKTOx728mS9MwU8VGGuPVAEY0ZGVMtneTlH4tk6EdV3f3Ps6rCPOm1Mn05
jDuo7472RHvJuhpOupydfLa5rXxKqzmDPr9vQNI0ztmywekbiwTb1bViKrNlYhzefiNt3O/lIMM5
i+e03/Zi6HrOIEv/vYcT3EijQ9HSOO+Q6yAvQtDr/z7MHBV2PkIDw+cq9n4xO0MNhU/i9w/AdR5D
seHPyLUoBKMcNDlTeaoUSP+EtyUOau/tSyuJDjxtQY6+b3J3pWLOFJtbRgIT9dKOg4gQHlK4Vn7u
1+GRIuPZxgKD+rOadl/wiTDWNVwb7yaHne8L3AHmfHGN08LsgZOSuykrYCGEDPzyM4esne1/NNsj
0C0r5TuVPtP2eL1klMnSGeOFrKUwhlJmR9/qGHw8+ONev0WZK1W0V+poF5jJvsR706FqxZqVGkzs
LJsN3sUJwU6vfL+x2FNa8PGWA3rcpR3fcLz25k3RULo2WLN8JxjdZAvZpavnnTSChkpkDe8ypSfB
dM9PCKPUXOdf3HyoA2GTBiZro+BDF3/tl+V2GurzmKqdkPrsog1uZ5IJV8HJObjib/iq+YVsTw9a
JDYBvg3jItrrPoYETkT+NUm+5TD6ApbK2cXcnKyG0dPruujS8lRsN3eSYch+lhrUaalSrApNPPsM
yZWeOQlfA8Be8orfOb7CKMcm1xzIKtep6Hglro6li1bRK9Im7idf6o3l+k7QT71b7zWUgwgdEFrr
ih5DiMAsd/Fic8QEN0SwfRZFQ3GboJMHp0kZ9VeWGiYilsXEoCVgtmXwu3FWAmALl3VIB4oOjB8K
ar8Ms2GIoWUVWABNscbSbHfWo8RMSENBh5YmEEkq6fnWozOyyouuYdsuwJBeDXHL64H9iqnrdfqL
MVVapdgIxINvcbMewxj867Ey6F0yjjBifZhARLQq35Ady57Or0is9Kh3X5l0x6PeYJ+tlABRKane
QD0TUZMu9luvzoH5wItZHUwr8Z/A3loNH/Nbr10jFNbneAn7BSh2U1OWNM1XUmqrT/b4i3FLr70K
jSp9KgK1nVphDJgsniImrFCNmzVF4cibfeSop+4Zye6JOgecXDD9pSG/rPjGlLJUGpAnTs2bpPKY
v3bFl/PY2+Q9hJHgeHHJ37M0fXYo/Dk+RXh4Z10lPtVjJRMs7ThO08Aw7hryQh82GHOQFffsEPbS
0ZzeGByGUjrZCWcZ474oceIGLQuLvpT1a92B/MpflnyaXQ/QnWagijJZqgAWNKqYVZQfOmooK/4p
+2CDtAY31oAuKUDRfiszBlG7ObrT4gvqQBTHU3qoNnSVP4MacGxeLIbx+Z5O8fjgxJoj4NYqebiX
f1CsRnlIREnBi25QqHS4mvPPaNOg8bl3GLkCzWETqZJkoTISocoS1YkPMkBiDs5FNQvyzRQrAjTk
mp79l7zkF7kklNrDueLCmPxaP/7vbGovKlZ7Qb/hWPQyVnDn5u7jGRSgjcckMDO3Qsfnnd5wu165
z9rIJVCgR7UqVOBWiw/rQvXKsoxHbiq4+t1fAt2R3N6PWA7nDCXcCDA9nqjrHhj2sHo5o45NnQAR
BejSosBEEHtvjXXDXYu3TIIirv6LcfwsAXoDK9oRUNwR3AO9zavldouHAekrMPYLm2vaLdiab1UY
GT/Pu/zdsXlcqKVG2AileBUkL59WBYFS+oZ0Vdh9LTtA7q/c7qEKFdew7sFn9SAzf7V8/USO81Hs
n/TMaZb+DKdSFWaYu93fvh740MO2rkSnqThpSV2jkcKa5r5W/gpbUgUawEG1CtOzgcto9YPjiuTX
Gfype90sDlD2cxWGL+VOqx53BrFxO6SWIqkRC/GqmqNOg1TwcQAz1thwaqMXMYYXUab0chlKFPDf
ZLGiGQfHJVXvK5qzlRH2GqwverK5ck+NPxqctUCTBB3Tfn1P+cMfVUyls0xcUJ/jvISpi9iSIpaL
cPSMDKzl1sW1Zie9qo8ahDKWO63WuL5Z8XZLVqlnkmqLKXvvNRAbY/N7Ab/myVhNmgNS2TaetEO+
99Ss6iThin0UbrhoDT2gBxGp9vzF/2JzQsh6eYN0OelreoZHg4TPy0ZU0KiwbU82U+CHKZm4Joun
XYUDzlvMI2SPxd7YS+f/5T+4E9FNu+6LSrd8NQ2LTwxK/UNXtS2V/4Ple7FF8rU6xT0zC7E1Imo0
5QdFywmzFnfQdeQCiCUhwW4PY60CHmvpO6eHm2A6z91M/rW7DIfqOVq5jl4v/FAwzNSDuLHktNb8
rc4K7sK2vtvFJ8R7kTDiY1/eV1XiWNhjbqch0k/Ml6VcYWBUmo1X+zymdfbgiYG64OZbxGHgf64c
KdEtX5tq4v25o69wP+gYpyzSMfATRWPCtQl+LI1s90HJCr+XK4/wGmM4FIiI1Kf7kDRWxpyncn2X
ShsOIqq8ysW0pzxv5zkdC+bk7rLGBcKnKVCjCXt5xJ5cYj9b5/FfhukYgl0P5iVGGmIjr4EwVlfO
6vIwMMZKSIKqwJbZ6XlulytAAS1N/wUxxBjATf09cRsCLeAEd6aXc2gPw701MHOhPnPnsFCaBn/9
PLVHXs92hSft45eDCEglchdq/Ei8lpajQQA7EHI3AoeV0XCmZXYkY1R48rLbwABGHe6Bw01eIrtC
iNN1MLjx1IqSe034AV1BL9bJRVdxCRzyDyGW9q1LM17OmVFSmpqtUKzEa4O/EV2ntq7N4XJyx8lb
s4E6U/+bailFGj8vor0kjfH7nh7Nbz4mIy42hncmrSuBJbYuhip1lsB20hL1ZgUzmj2LgOAF0HLB
yryMrXcP6BVNzbTw/PdyAOYBP9IusssJlOPPQ1tjNuF6LMq4ElHH2oAChEhZH2zc85BRXf9KAPIj
zvFJo9a2Q0/EeiFVw8H5NIUyDDasrW7lvZKL7TYg/SoRd9HvTBzLr8rzkzVCJ1WGOpkvwimXcwJB
oeal7zfWK0L0CFxcZssyq19oaKNLa6tNePcxxB+Ivsm46VBJwvleE4Cd35qgvOVw/xv1N9w7pt/j
7P5+yE3VX9jEp7vM92mBwGjZa/pU5LcOcoZfGzVC4Kgv2/LAChp6b+OLBAwyh4qPl8dfngGGl5Qp
n6Kv0/uhPaHBClAjhcQOppuCsloC/HcpzrNA5jzhlCcsRG3KJMVXZBPwxxYWraz9E2fdPf4rZg1P
bIP0umlLDTgCVHEc73uvpTs1ueFSYxJhrz+Ppxu1h4BPLZeGy8gLF+H+iYFZWLMbb+jrUXHPRI/5
Xd8syvZ7gDiJnV3dJEh3s5NKs3TPtx+KoNREk32ZKbZ8Vlfs0PSjVj9a0tVILwsvK1GmJzkCKUQV
rW7IwcwH/dSyw7GaiOd5mv/jyhcZER/8YzRncdoZx+vqR9QUG+DEIUTs4qlMHTnPEB+3lbio5egi
sMwxgHszEIO7JQXpY5hHzqe8Rl2EkB3bFeVx8ebwa/MH2gLuvdKnUkl8lpuK46URdqBr7Y69DCf8
yyaOxI6i76wFlJBXNpvw8XYVDsR9qWlavZ3Y45CdP853Ejp27uAIo11Q3K0VT9kFCXobcelKaD0I
EqHqWp0teWGYR+4Yy2/7k6+ihD/oGF2wPrwGT46z73Vs+VqNf2AHiQg8d4pkxbuVo/xYTRBrmK11
XjKkVgucmxKMrJAYoShieX0dbWLrWB+3U7qmBqy8z9lOFQM8wYK0Aw6hRjvLkSpWKxV/H/Bzq9e6
em8NCi96nPp+PbV7mecKATkdpB1QPBtektaGaBea8OfSdBjwyir2PIfomCZ1lPbyoL3zAMA0pkgs
Xo6p8Wjc4GWHR+aLPQNeJx8KjBvP0YVXt3kbTERiQxv/Czq0I9w3xy2cKOE1N2lhOaD8ZONt0YlB
f5MG4w+3i9glWigQ3B7w2LscP1Mid1FiwcjNd279TWDg7ugLE0hN/pnKqPVOF+obAOmZL1yGkvUV
4qkgxrPPuQ==
`protect end_protected
