../../../../../VHDL_Files/V3/RTM.vhd