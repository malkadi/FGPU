../../../../../RTL/gmem_cntrl_tag.vhd