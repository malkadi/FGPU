../../../../../RTL/loc_indcs_generator.vhd