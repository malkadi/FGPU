`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
BRBZ7522CivHLmvslhUhFYQoS567JwvGFzAncA2rwHIAIOoihCOXUBzaLTJDT5qPovHzDlW4yv7r
GP9s6lKwNw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
CGSFPehn4o5exPh9VqAEGC9Ban3a7ljD/wFVJ5Wiof4iJo3N7+ltj5Puk2trGNLyOVe/8cwCtokE
C3EHNPrzTVk2ekZYItDjGCLqFEdLTZk767UGKtc4+KFQ96gRMZEqc3w6niX15G8SK5RG7cenh0ZV
dIbp8Q4ZEYfKWH/MmRE=

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
G3aXPMgU2hkC/UtzRmAKroBoUkUE6cYbnGspL6n4cjlcyPs8H46gbwPbC2jNdTaMWd+WSerVIBKD
nvecP82xK8TcALyvl2FLWU2d/GuqCGUybrMythsQT8nDvb13Vy95OK4v7ajI+2gxF25l7rC0Qr/v
j7xd7PVR/ul0ChVSfvk=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
NIkZ8LYfCM+oWqDQDCOPVNn/5LpRuVnrhJyPER8R+9YWbLwNMtzqu081+IpI6nfE8jhuyqGOMJ+S
0oPzk7GaEseAdqBD+bUmcyr1JlQ8JjeaAU3lLDXNlgY6nO/8uHaEkpEe0mZmZs5zWgv8yzjxqkDo
AOPWrCo2lN+jFQJ/k2TNeH/vSSiVtB6HXA3nFY4e/eCw5rgRjeQzgfqYjdWqry8U0a8jgpzxwf9m
yRMRYo9Ios/T/zVLHR0JYSjOSgxXFB/c0Qdo07KpaAMFIi6+Z7C45rZyVouIxrApxHbtqoyaA/gO
swtvMWEQm4e279gQ7RfqtPd9BLx7hZK7ih78EA==

`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
GAuXN6U27R0wlFvl2eGHX9UJ+e0dvj1OGcZ6Yt/hA0Al5BRoN3D3aNOgAcR2uPo2k3Uq9uhn9eKx
XSf7G+8XNvMmZE+ysfGbox6tYuj374XWhhnQxLyXFsrfM56bRypB8jeFMn/hi4P37v6Vi/fACjMP
P67bfoFJ37LQpo42tvFOs5Wx1ZBmrrNk/BKiwMODg6GuBytm1amZ4nFTyHRDz5vjxqfKesH0nsgv
R9JwRuBOmNv1g4E5NoVCp2kemhpPGXtwndSfnPwKBwupzzD+hEtRvMChWzZ56nLBew+Sn54A8U7m
RtrqXnPXzdWyxurmuDufms+p1LJQGh4tzVbRcA==

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
maXpToiMo71Hl7B4N5vlvINvZp2Q7Ni4BiU+wD4RisruBbnDlOxB90knT3A1GldxApCQSDI55vfx
TiWWZRUX0LfkoLadGYU37/81cSuvFAURycbWadZzyN8qc2/SVUADxPU9Pj/VD85wLK3Jbm20/kZa
3/YA4HyakbaKe/aAuKYJ+VLUvhC2L0tbUKG2eMQub12Of4OOu4xVhEUteak/rtI8JGWOR5fJUl5Z
BUcXeiUvRWoCm87f7fKBm3yke5OrWuvQICjezRjnx+Ia/zFT/yoLW4EVzuJUKzo77dAwDDhcln5O
899M+jy8zQeHABRBQyGkYvtkXBAMoPIL2lERUA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 103440)
`protect data_block
kEU3Ty/RI+ZYnh4G6ri5OcgjA1Rj7COU7wXrJBNpuAwZPB9pV3KB6IA+mknW9bxnS+M9xwkRY9T6
IExOG1ZzJSUlHkC/W/fo0+KfI6N1enL+qAozSUA4QtrhOl0G1lnLbw+NDvtQknOMY94xWW8xJOWS
CgLvrqfDgak88UvC34FlBN9QBkj+6tzwURDQK1g583KeH5CmIUQMEIKaOSb04/4YbKpQg92d+VPD
7sYS22ZheFdCggUs1j/Xj9TL6lIO9fdjJEGVO/xnzJorVLVE9OS3DY+3dFH0kaQlr5V6omqB/orl
0jnPvgvCOAjIAIVtqiY8sckI6MeUy//d2+Q+y5jiTUHA3P5cYK4d9+9H9h6f/oCTQiupgIdYrGdB
zbTw3QBziKWSTFF/mK8CXXIgNzxySX7BiYI1MKW8fFuXse/zrg9bPlQE+HKQqbLj5vUuuz6VkBll
HL9leTC22RfiYSoClWHFp5y8hkKVnKpzLQPhvXafvKZpgdrmMvkOnhb0HU51nUm8g6uVpzE+jPUh
2mqqtGVGoX/KFxOw5I4yQi+Px3FLgx/hGylEVlMvZokNaBLLmt7+GYVfGD2qmKi6DMnpE0Zhxht7
LIRF5LajkCo1QJ0A7DvhjXcUiiOVVq6CelqyezUxjjMQQB5nURLOAuk4PKVkYXCEYxIMBH2BnU+R
Q8H5rJPqrTs7BV0D0SoeUB7J47wNSHuO2Oo0G++F5Iqn1ZgAFLyeX9Hb1LlX/yYPAKCXrzVfACAV
bfNNJF4H0dSA8VL5m/U9avrux1en3+bBXCym+iJgCGOgfCpyQSK87ggtCuKOa0Nk7w5/tEX4EnBs
HY6dBexA5u0SLlbtWmnQ9EBQehDIHALozU5EI4q/cLXA2o9MKfALm5kuPE0GtahwXwaoAbJwi6Ce
E4l//vENEqmeusnYoPfPPyan20oQjAGDGjejd//rUCB5+tkI+Vj/ImOtEjy/+w05BYBLsHmyCC54
IkxixAiyuLyOhdJr7uxZj3mewoo8yz8by/3ClhT+rlSv9YecCtL/t33m7lPzuEEft2ToklsnJdYd
XLqZSYbXCs6hy0bTXTHenxLoc7lOLJbDskI6vO1xeCF5Axamr4WMGw2giBgnIRwBH/gsH+BIXDHP
xcthzxPD6ipL0KeVbS3KmHXeSacXyhI7QVMIEc7M4UQOK3v0DgulHMh8wuUPK6oTEPC7nGFGsZS8
X7YAgypmG8EJp/VBCwEJMsLbEKfQrdi55lugci1Vm+Y5I3I6kTQSBzslpsPB/CmS1kdC6lJf9xvT
e0CBL6uDQhBmw3opSAaGH9yP5aYh6oymlsyLbhz0hhjlDayfFMDxq93vvrIC9rD6LHh0dOn6RhTb
gVsbnotAEwA+PbgbrqVS3PNr716wbShn2x1eg/Fk4Q2PyokuVY2h3VOUpNO64zsY3d1UQ8u241qG
d50iTJnJ1uXPHVvQ/QTpXPJrD2CiV2tXShW7SCbpxn8g+ruhVwkJWbUJ6hUrFqgyPn37C1TtP8Pq
xHcD9Yy10UDKFkT4LLDxmrf8zYVZ24a2ZILhVzcOlszTzwkV6nGacjDBGAtR26eWKEufDaRujqjy
oFpN9GY7oW5Nj05m/J9v+3OFkx4PcopBd1mEc+HAYMoeO8xhNz6B4bQdNGzckrPVIL4gC++8Y6rD
6XX7moZl0xlFrpzWkDkk8K5gqJH2xk1dRMo6mXH3HgAnldBjaYKb9GW4SFnvBMdnlzZprp2Lu2u+
ec3Vo7cmqyyHaqnJ2PhQ0QUeloMnS2NM0tMdJ6YHwYuQLB9Ll0dERkXKvS6mqLVmYyeHKKF1oTb7
Wa0qrX1DCCFQ3q0nX/XeFpe5j88iG8xKJ5cqiR33bZrNpdtar6mzCJ30BqUbWUsuf5PCAOchpEUS
UfQ+p2m+l63DHhdkTpNTxDxJVsNv6nyjY7FK3humdYf2rfeuS/ZlRrb+fqtwf1wdq+FVDLbYh/Qx
fgpyy+7n1U+x5B+Qx2zQu7PwWXZPODwhVa+0Hczvxrs560uVpBW5W/PjMDISowrt9dzAoDNVpHf0
vVD993XME1mmDIjK1oaLvdbcNOQbJAWzcUgz5RhHlJ8Dd9XHlPz0oSz6Y7wDQgZIEruOKf9G9hVa
jLvsNq7d1de6UDwHGQ+8rf2BnEI0lSghy8vryUR0oon6xxhEdDfPbeqhJS6v7BouGd4rwR5+qxit
ZhZw5ld4viL8coCQFOpZQd6poGtQ5MsXiwudstqr0bDdSbJMKOHPGFNGW800UQDsfARAbYUycXKo
WxCVVRSSrfWry3l4NEg3xRdLLL5MIseAcDT9PmC5HO3xB53w9TUipjONgGtm1gEnHMQ5gCNatQHM
6dsIyZgYksuKbl3Ei3Etb5dZGtYEZabs3cEG5JRYloTHefyi5OEQN5oFeiCsIsS2mkvqsVKjfg6z
SBprI8rDQnpqwtcPtdm/zOqSll1MD7jNUE303ifNVtZRx7VtXH7SYNgloISVLCEAEJdNYz3jrDZL
Lnv+0eB0D0i0AsXQiy6l53OqQUKaW7mTMp8RArCB0kLsj0NB/Xl9csAuZfCsg+YfVHBoViiD6RQ3
y3uZ8dbSQfT5bfBvhcqI2nEk3v7+BOdy4t8Jxr+5qWcHLehoywoB2vnu7EGkCTIORuQ4Cug7pzVC
wn+fybN8nqfQOB5LuUP5zeUDxf9viWMW5vtrV7vQXIzgQbPxjgBoE8Ko29Ugy5R7ItkBJ70efEXm
nnQPeP/QPzICmKT/O42hmyCQDzdcdL6qGukeg575e1kdUnN7KUhH5bJ3ozJ5z1IGPlWnrXK2OjLv
kj68xyrVj/TIPEBCiVH4K0NAQVhplMCWzz3NOpCaYbRorzfPE+5UH9m70C53kg9CwaAIooiq7drz
Vlw81zYi9iTiScMsWxzXgsxuYU9pRHcP0yjbIvXecKhaemSEUXCC5mJN0JsolU795viSAlR+FaQU
LAMnhirYE5LdObN+Zr4AHjyS/lAFn3Nyhy/fgoMXd1/XmvwV1zxuOXv3TqnrSpmx2/NBDaeCPkqb
JW4HhkwVTIyCKY7sRci/m0bcBhGMCbNr2Zlrdb4xyzmBKIw6F+OQh45g3ghN8SlrKjkzLeBe1fOv
DuD3IxucOQQQhTbBjqdxP47t80p+VfoT0EjLgBPBelPZJjyrJ2tKKLrsT3IGerq/veUBG95c0EmM
iMHeyhaK9dWitWCNc35//nOIpPvU7NuUp87z6oNgVUeC5CbnwuJqjyxYw1songnRdmUhon2NeyMm
BGyoS6riAs1HuLCAQxoFWxgwoDh4gT2+Hn2jJg6U5VTR28Af5itHJt8qndOvrw/Pv2uldOOM65T5
K7IouJGq/Hh8F1Fu6nUoaQ0QUqCyjrf2e/TTw2yG7inkyva4hs98HGlZYRmjDrvZu2+sLw0AR2tY
6hYWGSVAijKIEkAfcFve1zigdD7DBhfb+JolgfXqPKotBiWtzGYW2zKzHeB+89f+eqOZPvVDBp7M
QRwnZmY49eavzNCBKG0AgwcjseSmnjpymhIOJ6MncWKByhwXTwJPH64SyRmbhmJg93L2KlTJXYM6
djl5MEi5rTwbXcHWje0HuTLeVaWTwWrIY3dZIQQK+D+ZuuJ7ZlSCKbhSfE6txwGCp/QfHjbxELs4
2v99SOsYPjQ3GF5UXlexLGosAZ6Nqyj31C+6ExwaZtjZH59oa5f3+YPqV+5GWoGBgLkfYhmnkTul
93J4B42LXMvfUOYOGgEJLYsVK4M2gQU8S1rOcWEOWZNatMeF129wIARf3jXfFLZCDZs8pxMmJ5oA
QryzGu9gbbF24WkmYXQ+IyZsuaQjqBOtW9e0LNpSVP2F0dq0dsCx6J/wFP9UOdGOGe/gIfKaUjYK
/vd/ARM+HJ/JwHQAivN6rlsLH1o1+OkhBsqfCPZVfJ/zZBNOVvvwP9V8lXGvbZUQydQsbFWGEVFy
IKzCMuk1p3urj/MtQTH6pebFslIEnNpehP0vbHTHZUgl0G5/UwSdo6o+paBwiLNKcGvQTmP6Iawr
W5nEFj9a7SoXk86D8oahg7S2VIYiwdIRAQQR3ZZXq9uAbEpIv3qDGDID+3jjYYnctwRZOF17Wb4V
1n7Q0jau6OP39P9sv/K+J4jzo/3Jp4fO3pyIrEAAwHhZ2rDcqAWUGxFO+rtauQ8MerciHy2eKCf4
FqJjd9eRaTfqDWhnWcuLG4A08tldYpbKu6mR+VK9cRnNNN0c0vUKL07tWCovvopIAY/rnJK6YO6q
w/duU7LF42jYpLIIEX1JhTATDDoNP9L/KyGrOUXJMMy3PDnGPEZO4mnQXvVuHv6qIra92+iDejfp
6sukkWknO+08PGz3QCxYNbf0dir0SVun4sA9A/ljN4Y5MLoAVX2GbOMkuiDYki0LVPC3rgtCP1SF
tzKpkhW7bmK3qVfCFjD0Q6bo3Qik4ViwYd8+IVuhbUq27KD1YfVNr++nQbweTFgjKxL34PVsnHp2
LeJR4vpXUmFff0tlHb3CClQaq+fqByy/KgtEFx7NS26mTMVrMXGKrOFyQlVBAw7cfEE6cGjop2HG
P8MRbigbu2nJIw7pjYlgmn2cJNGCxpGAMPtSj4qdvwi0nBD8HywvqOej7CCnrBDrrTSSovdGvYYE
Z0C+MSbeie+4bwpIfO8UORVl/FGZKR8xfjmhywvf9rxariwIZhDtAL6qPfOdsbTq431JRL03KFR7
jnxf2xPI58amZLqZ/MwEY+YgYC+UN4HyaqzDvKISzNZCdRtIvGj6OKNyJllbO//v2U6OAaHLm+0y
GLoAqa3somXqRgh4vCR7gwHmVDpsB1flDOOdHIKL9LqbS25wla7xvqA+by40dAznUK7oyQGIAVQu
E3nlV7ypVNAP/QUjXkME5nb3sbCXniOwEZMgk3tplmYwCNYW7e0PbnVfZYbpZtiJdilG4HdXXVxK
a6+nFvRxyt+MzNchvMFHfqtT3PXec+n5DpVlBWst8SQjr3lmO95n17tHstJSafGPAqMIS0C918F8
DqcuY3xLXP2orsj+2fszwuDDaSUJVHtOZQJBaKiKNpCvO7ps55mEwH1rifLoLumKfZfMm29Lq9LZ
e8Jj90d4m5hkvad/AyfkkNS03ZS258vlPu9/ofptV1IeB2pM7Bwguxrzyecgl+g+UH6QB81b+Ugg
9MEoiJ6EFbjqIx6RwG1kiZqZ4QUovKq8OCLHVA/Y41zrMUYHNqu70tTKhCbGr0TC0BKJwHXPah6s
5fiThFDQoZGoWp/Kwu6PzaD5RDqbtiR06s6wobOydCGwRqzFdcA3IExxKfkqZNSm42VY0ZQUAH60
8TdOaqc2UQmg+5IEUP2v2tyHLvd3PT0sYdBxaunA0YLlyD0YXQMyS2EKH6Z8cJ2IajVCUAP3Ntfl
COL08fhitgppLyLyfxtToYFU0Rv9lYBPLZWYRKla2Y4p7xTbRVe2aNdeLpgMWL2VJt/48b33p+Oj
FrS7+Oziz8h8aQiN1ZqA/NMmNs/0fYXiwJ1ckKSp/ZmXMPp6U0MHDYIHeC2hnGffANjnCtigtEbE
HJPc1tR+unKT4FRMV+y6k0skbCUu9Kp6l7AhR8Ue38UtdJBMpFBU456Y6MlI59Vw1hQ8lcr6Vusn
bu19DXn7u+X0OFHAl/QaWVoaUBfbthuIdFpLp+X8Y96vvoKMXKeHSB+Ck/v+kUMCZrBwQfK2B3Di
1aS07lr3JNeTthaB4rD5Nqwnd31ZsPW9zlL0DGmOxS1BQp/4pcrXFjJ1AMiXxaqRBij+IZMwhLM3
thTXoK//iWPNtP8zv9mp35k9fvQ+1G7Ld/Gc7TO3OI/v7LKBPqXXyrGpRclyMA9dwsrwNwf6+Dxn
RdKuUVzFjDCpCLAE7jG7o1vaHp4GdgWPc8LNqinaZ7M7gejdYdNbQtsBXkeiWc3B07XiYjoA9ktR
Fam+YgfmYvv6qF4Hv0a/Ejrp461gTzLTqkvefbLMP4zz0wEmdWukUiOMw5VaZ1gobwnJkrq7PDpv
DTcYPHefSQBGnliUxUQTYarMCXgEN5Vq0tgaSsgd/Ik5w9RSwzHYLeMbs5TT/G7kYzjI8gozEZB8
bfMGc+xVdxSMKZjc8FM6I9t40KGL3p+0jdz1OZff9vdrFI7VLofVwqTtd8WeYehY6fzKHMS8QdiD
8ePq/7R13e2o1phF6/nnaaEkDFXl96z7FfRqdPP7X7KJC6yI7seca4URdr+v0XK175LJdLrctx+6
Lfzoetruq/02E/OnpP9CubipYJwON1CiJVA3t2hjmVt5pE2TNTkV8mavAHV8i9ZCflMHWI3Mz4vR
JNzPU4Cokf/t55f+6FJPh+Bgi9W2bqIji9aKN0JuvMmxWUCBv/4A4s548Z84wIhRLKZlyPhbpbBi
4QrylRzJQG52ZMQDVn7Ixpd/f3A5wbQbkHa1y+Di+dvui8JO/OGAC0tq0yZmN/IBJAJwYEYGoHf2
ZuTFzQTSLwZgkn4pW/XKrp0vtWvX5lqMCwc/vVXRfgAqGWxzXFZuIvIrje7XSI+74WWFLnJ4B42B
O/ClWo49Lnm+pnGUxe9gL4a95qcLwA121uoT3zcGbyyY8Mh7Shr4SGSl4BOn4myN+VfONvgCoQIq
LKzBvxBNCbKns8+GL4ruA/MAKLh0Cjpin6jOaKbF09kQnly30SFzHy+Q//279K0S3+5dFMTv/ZvO
NhQj82biy0x3bUxb1dLbCcu7eEkstZbY/t4pbpTLaO26/aImuawX3OqUsN+nAOYKlMx3kihjjhSv
YI9Xq9hq+Hr0R45J8mFrJsSywbqClOfgJ7aZEoN3FVsTjTnv8UAwX0uS4sfWl24FDU4i0121XR0e
D8kw4dIwERabve8AdAK7LORfQxYYiYvZeP3V3Wvc0foghGioqofO55eSGUrt23vEqwW70tP7UTcs
n/TwOAwy4nKY2aahQvanTQk/ZDdnQw1MW5zDMc/sF4In/j+USz3C71iqUVr5/PUi2iVDJz/eAvEd
rKRb4dxTMP1SeLUf6XLrmgOFG1DD+HKjjzU3HFOZpMOtP/cVA8BRYVQu7mYe8gIZyMwnTBCQLfue
T0XCuxMgudmb8iMdzLd5LGlOsteewjzpZHvqplxuhdT0uQF7thwtg9Ls8A8bOmFD9g+zBij+laHQ
3RhFujus0HbQYYkAgXCsjr/TjVpankQUZiAucW82XktH1MvmRAx2AIJpWjdHolcv4OD7PIWmxIPJ
NaTcGcC1Of0G8y9HMS3hpvTS18HoZxVu7S93GXakULWFi4LqZLQ6IDLJCwNfd/2cXmXZ4SLRzyhS
j0YMpKTSMo/B0ldCkvBpreP9j10A//eVuRuXSiXN2TaFVC3u/a8uXmogqgJup94PhAR+zlAygdL/
Seu7llt2JhhiqoPkWiaSp1HULrgvlliPYLJ3Stv8SkFPkiDbZSyGd0F8lCHqyEPMnQ/xtw+e29k1
PBSala9DdJyZC9WXhn4OWYoQ60h5xNwvoZo08NMlA8DpdY4tZ4lDdqOQNzLCKPG/V5kvBFKrf0+w
uRMCU+7WVsdEejMZRYw1W4oDByu3L9krIdtlugcNkNk9uil7QUxl8aFP4vBxQU1CQ++aYEnMFy41
pb1yTCEmllaEhWf6oQDe3s1y4wfSp2rNoQR8yTWrbgkLXJmS5/VB/vuXh+JWNxaaTtw69dLK+muf
wMTOKIUYZjmviK+MPAzY6GWUp424XX9EWup7d2jN730HDgxq7wgQIpst8qA8+k+EDsgeMDBWD/xo
Lg4PbpQclZ+WlveAMz7G+1E14eAfkDG8bebyaTnNolqAOgcOf/Y36sG0TxKBLXhbjrtINSQDeOhH
gRihofDWwvShIo2LCC8OZY/CKRn5ARD06MZerzc8cuHfCtrsOptNY11/IV/xn8FUCaqWRlvgJZrH
Of4TGT9J2D5xPgq1Zoodp2mZEN1PlOQWl4JUqIbXoufWtd3/WLfnS/MFFdUAi3toP7qeLGy2IO1t
ZeuONgaIgoxPiyG0SRNkU5Xw6VWg3If9LcOaZHV/ekXP5J0QOuTV9IJgO9Pxg9TvIz70KQHYsyHb
ThGWh7Y+vOBi0tUemFAdlSTmvif1WVS8M2DC/zIqDnojHsGxiCcJpQmIz5t86Xs6VtU1agj4ZcvS
iF4pIfv80ENDizs+yzBUEC3mZsiB703JKM7HsYdBGa2mmqdeow9HWQXLYM/vxHiRqAUqggjpgdR3
iXjdOdRN3+aadKabQHsZMx+pSMtBlQne5IY1jkuHuy9kJ4JRp5Dk0XVC9ZJ/F4O3oVRfDxyV5kaY
hcFZg00V8G5o8RGQ0J/yZ0YOKZrjZgo0XVf0YnZNd2agwjIlECQgEvfb7iSeGqYeJ+seeHAJInBA
L/G5U16HhcNCPllvIboJM1ZktvY7/ZuKz2rh60g81Y0mFeXspwVml3ysNNHhdW/qRe7Y8cU82BJq
2nhaNxZSmlZdo/HjDhVPueTw4LXym2mjqnsKTEXzUJ0EkDwj81Fll/dXczwNF90T4xnk3UIjQyXG
LbkSkaILufkiDs8l9egIbzNDEhbNTExbLUJhg0yRD38oFC00V2yipFyXVoZVxR6VRSS+eFNGR7TF
5Q43skjwqD7u3HLgIM96f8kCnNSJzehHdsuZSZ2UiZspLNW/PORLFvOeVb1SPS13x19cE1XRKqiq
yk6MTPiH+QIHeBOobonODVSit/jwGLKwRU3gSfhKUVBAe00TpnEd646/9TkAzjPC586un6S58mz6
BtB4xUxTNH2XJdILr2pulKhwwIFpEyl6mtTPt8/Phjnyqpg40p5YBvi+UlAOhlVsz/hRpZvbkLs9
X58HbSKarTXUV0IaxNhXD0x2Daq/l2eroPU58vs9LernHX8Xgy9+0KDXI2Lp5exMf6cRFJTA0I1N
meu8O/lZIvyDSa4DtiCl9Zu0AXn3QO2u0OhaLuEH3k+3oZ5HOoOL3dyJfOfblw5ZXBSOLs23icG2
pOiKkzVdck5B5lJ6nNjvA7aOBwJOQ7wE8+/omZjPrqmDaqR8W8ojha5y9ZS4xxLBTo0jZeHItSOJ
yddUJj81tpgcnGLOZph+9bb/X1z79gtv7YyRfqSqF0uH/3virrnVMD8HOSOKsCoFWexKP/66pJIE
Il2U314ce95gvOAC9zcsnAN+mlXSSyfiNWQo2XoABenv0uqZQUTfOfePmxkRQZbM9n6Ie5vIw8OH
EH2q8+WJYkFydDU+XUzeXPmIYRf4V229nO/WrFnuzLcIUuqJRgOdr6aQpgehxGyeEaE4TB0cSOCI
wApaaPqvwR4+D7LgE9vf2Kk/rPi7X96byo6aAOmttRgBav4H/5vCOlKzEj3pPgayXtPkXrVSRLKd
s+qFVBHuYERzihgYT3n6Bys8zseAPmPERlUc2LdU9QBgsol/AnE6RHkMeNaFphAjfylLk8sI9kJ5
qWYWgEnNLcJyZP1QnnFrPnh2RGvVHl935DKsWixfL+PTwyZnuRb7w4Bbh51wr162nJ9l1kAwve5p
qAz/cIHzmczY9FZlM2x6Y7lIrP7fmefD21QGK7rnk0IM5DU2SStJMrJ3Xy8ywXtaQB1QOT3GlQ/V
vdyj/76k/ez6+a+mQE7fmeTRBvUTDInJ2I4anAgLQ7pJM4QNw6O/WRqfTgz9xh3je75nDKIhJFLn
LbZ/Lb2v5tQbhfo5OdHPJnJ8jvscl4sJbHd0FfzTVPGfrPPVR4XSXwRJ/xRqATcS6LoCxow1Xy/y
AHrOHjqB8EQFfSSWSV2EFqIGkLJp1nfKOqU1LMQJY0XK0kO0zZg0Gd4oeuwDUslq6kgpzOcd7dYK
vcntpsCvMTuTXqD9XRqG0p+zPHyhdu18vOThy/NTKxL/Fjjr4S12eM/w8phw2fhGgTzcSnH8+Rfi
/L6aKP/c2AyBpJUQZA9BkKfI3nUeRukpFkohX/6wSVs1fywECIeRXZR3raPr8W0QFmUYOgx25A3+
e9RWGvC8Ib1mjl/sRDAaxFjf46AM8jmglRWPkdkgj0BAdwV29yGAKpX2FuIpeZmfBnlFHE1/7J9l
KMF0viNwq0Ar2U6lRml4Riha407MLM9VJzIYYFXVadAOKoqwXJ/DWuA4CVYt/OPD8GPMdCfhMV3I
dA3UE/kZP7wauPdd2FGuN9/gd02rgHORkyv/yxATZKacogKtLnr/30dEvShkKXn1fU+jDIFrU+gL
toZNwyzuGtU6iq+NI3ZXR/P9uQz4FDsYKAsFoi/b4fsS2VnYMIcGXwm582U+1bVwzGw55PAxnAQZ
AC2YI/pWg+4V6O8bxkpYP5KJiHBsY74ueTexP/ipdsmWeJxOroA02j5oyvU1iG4p94Q6m1Q8pXT0
QsVX9UuSNytc2m+41ltdJrdu2ByHMA5kkOAgBgbOr5+/u9hGlwGLzazynB7v4aNUXoCHqb7F6GCo
BCTj0zQQ4MtqABb+QbvrTFXh6bTk+h9UGiMAZnV0nEcT2Vjwhy4/d8RM8gzOPqkV4aqanYmeEvCE
FUcfnTLMn5+o2CuTZZ/g+EBLIKQw80NZFnctZFaYoDHyuGy4M9RZi61bEYST6+UsCw/Xb6Oj1WIN
bPZk2V/v1MVoK5Y+brA7kvLensNMY3hg9XLNySWmyLSvnA5tk9IRTgkCw3Ntgm0HRKz5QsQn1SUL
znb8LO3NP5qDKopLiFr+bST5ghd3KBusJVYv/jmuT/iRudp81hwX+3UoH2EyDPY9iqCbb2/wj2Ib
pr4lGWygPWA5bqX4vCRoIwKX18sbFw0QqpIJQJsAD0pR6QiW6mg543yQo7mkPYpRu5GlXOorhjU9
Lm+tBXOKwzDK/CG9Qm2s/Ez/HftFus+XMdwj6lW69eQ7PpKOveJ6317DFPir8UMw70j7rVEhGwR/
t7DHaHZ6eExjcVTXNrRTjErVuGdW9tJme/tiwBuJXqy62Ye+kbpMF3610syWD5zbMJgd80jbqEkp
BYKqfbWWs0GREjEwcSUKP5ZceWVVERwsVqNYd8v2DxcncTzFMNQ+zz9nEtwS9KH7HLqXw/HYYr2B
aO+R+hBpZBQt1wI//usSS7TtLUIgbr/DwtxIdQud8XDc2wMhMT1UxSHWVuQuvcbWiyDPfKrPRyOh
OXgJWimmiDBG5yhrJIbpXNCzx9Z2NaQbvg+4yy8QmKzRodxdzvsn+bPH1S2CM2EBTdmotvSXgIN4
tyA9epaJzaXQfBJuTf9shxY/1b5YMUyOi8AdvDPCFvAi9usnWEpmQ55kvE9Gs8PGXCI1f8tX+jwU
UnuOwmVlDdmomoMK43CuoWf6KzHfPAF6M8WvJXHPZhONal86xCRwrPRIa2VPtNM3947iqdP2QkL5
Etitif2lsqT9KewRFxTEEEJ7D59v9SYU26lRfvCGtnzSfSOFYNrPNeTU7m7LUgJzAcpVtbSpEVud
ZILCAf/Timqi3JLHPinjfsLVmWJW0ed99aWogxBBbfkOEpKAh1KAYfjBUqHiLAocjZQToMPLmkct
pxA4XcLsC4yaZxEVtn92B5gm7WjeVJZD6JHAkNQBUBNcUQIUiipXnr9Vw3fcCLoFZbR+WQt0Kgpb
Br+2c11nCRD/jpxYv5b6/0T3mnE7hyulQ0DYR4C5iU4gosozRc69QaZixtiSC6E/rH1T5GoxjHP/
A+gCgLOUnEl0xAtVT6VqOfB9b4tNuaHVX5y6GJcu8Fb3gdJZupus7mkiqSc6rVVRlQa0ZtvSUO8a
zN8A5X+MMoDVCGejeioFF5VslhYDtdxol0jsc91u6SdYVln21xhKbv/8GNfh1GbK5dYkuEWM9Jmo
vddH6py7fNUCTBEZBbVK84fu9Zs0w7JD9rTo4agt0heqYQ8fBGx5IlVhcNyicMGZpoxuZRzWyhFH
JBZdBfRQp3CzVBInI090GuU3hAJZ6tWX/Yt0I73dgfuGm+4iHwJRq/sAJYjWM/OfmdAYWvCVMkSw
Ssz/0YDm/yj1lgzLsWwwB/+MrGhXjjpskhNIP87wcWTf2lLrdi8J9ITxvoa9CzvmsJefWEKnGbx+
LMbJYe21d9LWmeewamHp3pO4w5qk9Z2vBXg9tNbhtVKDh4iWILHtCLiH/7EwGHnx6GYPUhafSz1D
q2dpRKQ894ZRMx5RTpEqAZWFxRrOl3aSKwnu/4QFR3UyzFzCXkFis8PbnSh6hvKZEWeQ47767TKJ
VhT2yWSyYxkEMh6aCHSTbRvM+hdSpi7CU7qXmIj2CDMtl06gimlZAt3JGuSiepro7fRuoUiH9Sbk
zDd9YjdDgXeFG0hlDX4fuNjkVp/8IOyz5iinsq7qv7NUxacNTLRwbBRUIgEOgKUagNp/WLLaJRCs
iBIdAcJdkz7FkVo+GMJZQmozAot0Zz3/habqeB0QzD4iUxZ5gjREOHURczkwFqU6HVMwRrr+o8uC
ekHw8RXSHyfS6hDjAfmXPjKoS94qF6XP2SSQ8s+1rcXJ8xto5lTno+lqdF4Kej7u/oxAF8qyekcK
Mf+4i+UNL5ldv6mO41lkahl9wSV9Gv81r3V4MB5CyIaQNOemVBaFl0dUvfFiGuF8oR1suP8uK42X
Qw4QX6HwLfAXJWpgmQZUs5sG293hpaboH3WdJ5s/DcAXPEUkHKYN6vKik/IfGRmKxB4Ce7F0NWNW
7U/y+k4mBj5KUS+PcM3dUZD003VSejtuefvZfNfh4uUmFYScakSHAZk0dKlwh9Zdl+lNNS1Cccbp
vLsjOlWsyC/Qs3hg8Sy9gDd4M80jb++X6tTD/YGP8/wij1S8pXgflrBokTKPdN1dBvviwoEPBmXL
omFv3J18o2NDzQW8vCBcRLSyCqPzUNrYkJOEP7GJecmoyMflQKN4usRF6u+QO4CI7qQFq/bszhhe
A3yaNf3mGzBrZ/jOJiK1hdRE93cQKXscRsElIukKFb7T8Ut8gcbpOTYIPlBY4gZCryWg3bj3zlwp
BmeZxmLmuIX5hHrNWio0/w+CXlfN5VT1eRjaCywREq+GM/mXYhJERbCpmBhfvRpONcmmN2+Z7h+K
2jzLyaYc+igrmZaJyCuCKG48XFcUepIhj4s/DC+z05laDr9uhPeEdIrY2f6YRjgp5hsMvaRkW/Z0
UpX8QX4yH49oIbColYHnFQN0GU60zjy4pU+nz+cVWTSPWDbIrT6GjpJUQsS65sNf3O2Arcq3aWCF
jvwzL4EYeA+tT0bOnb1N+DdfDvr8HGkCLNUv2AjPVHq/SMyTA3/9fnW207lCi6ouOsdnDnZYqIAQ
v6vJi+bKdmU+fs/1X6J4/dgGe6e/1gB7XDcjf+WlM8ojSHvagluMld9BWt+0uLnCBiz2cpZNO20B
x58ASIK9cTfuOwLcBtJUdsF4FXCsotguP5aF7EYWANW9aYRP+38JIING6LV5Mt9DddBf+0R+Co/O
a+UokfTzGYR82vNNZngnh8ioiju1uDghLLquezxaewopTxZK3cRxYSk0f1TTmdniyKNJu12aqOii
lVe851P9+HjeiOx67qnE1AM81h8NrecasjpoXC+M4ItGrQEqu8jg+Ohp23Nj73i/pSnW/st4kr/k
W/ntKXvvaDQcUv7P85cNRYcc8HctBA6TtW7UFDDC+noS7G57QWKHp0kwnx776ADkIQlRue5s2oI8
VN6rgJk4wC1DbNhxawy5jYbJ65A+Baz1V+urvST8dDTGylRDYi+kyRAjLNXm0C1Hrf1xnB1RqB+u
0pIbcTY2bHovSbt6vdiNYpHPKZZlxBhIVqD9F0A2mRbW8h67ur6wzGxAhzOm8+fVftI8JYtKFcHD
4+/VKWveYgHrzXJK9/FzsrST6zMi7o9EuvKokSzk3HKnszzeFqEw/NyP//EmPIkUQ7uD4iq55oS5
UGEvH9Syhf3RpzCbvyqE1T0yN7Ia+ruAeKHKnTHeOyKOhLm7BEOKB1KfNhDtjWGVvVe8xKvkwkbV
Z7u2gbdXqhKKWe9kztfikuIqsnOPhR48olXLWc1Hw+xySA2L/JJ/6eU7iHl0BQeZYhqm9cG0rtld
Tnh46pMn2Cdm2R+iK6+yLsp/Ci53P8z9tbfVkWkUFmxWiCh3fwOHCe2kONSyuv09XswQXg0gr3NB
WXzgTUtNyt3vm0dyTdgnbwLYZsnd1gEqSTIMWKNjkFDY8QnZdP7HzlHZokTKwUMLD/MkdUvHlv81
UlB6yF0HNzoiAg5waHdLOV6tlJ+uunJsJIUXyfhQmz/f0rUrzZyAHCRz1F3vZpedWTc6YN9gIIVW
/qcxp97ISjfYbgf1xFw8JrYdCSneV37sMIVaHRyuMNkYgBTS7lnKpI8/jYgMLUxffEsZK0MUVPy9
B/+Q6kZZfhbe70LiA1NMcigqDL9RP8HfGX3zBX8sBdxTU6Q6DTYwXp9oGwwWOOPSCEGTPLmXtwRv
Ht+7cZXj+96ichB1ENEOhYhAWLFRfXpGgxENKe5zvi/3K9AfkDNYxbChEi6WxJiIlLNZFSatPOKF
xkPQiRJEgYsCRzBCZ0cNvSHNMjBseWYc0TwnshCp2PwRNCaiXOgiktETYvuQcCDjRs4kUvWWR5FD
5TSVAd4A9YgcLrh1w8Fj+xW14u4UKBvCjS/HrTUatt0a7OcuPuwFSr88lqABMEnDbnMsW3rSY40Y
yrnR0EevIDaXsLGTcyzsS6bJZSbiXXgHVI06InioiRWHFWi097g5E/46xipKNdBEGDNSq+dcwhOB
X+FbcUs/agNvwHOzuLuIvxFKnHSTHM/txvgX1yiVZolDOPiMdUr0UOfm9SGBf80/jr+FByWNvtgv
+cHJJap+p9XsiEyOq+e1/46Loirksc8Whz773637RSAh1M7AH93SaK1T9hgRotv94ssFj71UkqUZ
iCKM6ryd4Mr2VsIGIfMFxS0Zapiy8t+ItAqDmpr1em4HPHSg0/1nfqTEkIlFsq1Q5OMaM4MBhz2v
6r/9XmqX2pP5avwTpS92wl0NEXSlpSGzbVjajzRMxSJcPRQuOv9duVkG1OBWj9kf1unVgvGSETMu
+Gi/0CL7gmZ9sQcXXHMHtriPsrokqwwiJdfao/kjrW6ExKXqVUdeVPbkwKtWyR2v25WmfjdTLmm2
jTmPR7lQfCohDSYo3WW9N4CDwJUX4pa4y4R0C9u8QzOjYBYOPyszR6vYolaKyklWhDYhhffZbYV7
Q4Chu1LIlZencbpyK980xbOw+zHA7ATu0sktvPyBMgBAiUinTAEvysVmOSVI0ldLBxSw1+ufnRBv
yryki2/zk9auir0CE2JaDQJk+sl2MQakYAXnTFvQzEoL09YchqDtGFC8Pcv/r1fSvexwkqzAwZX2
iwb67FXgbKSdo2r0PxpSCDNbYBS/i/rG+aL/216ha8Zd6sDFMHCVtjIRu7GyyfmmMMxW07l5mOLI
+haou2ohftMq7diOUIEsLQpzD+DohlYpf1MCpR4Zaboi+UMcUh7V0ztoaILM/GN/pH6QMXazhK2d
Qnq6xhc169YbZGYoxYCPrs2b4NrumKUBF0TtG2mLVbln19negP4BIUTpTjqlOACx9BcSkSPjNC5u
hdwXFlXYVjTxmYQCFOoZ/e+TGiJaV47a44UknM+vNI3CctDoH20LZ8N7NybSzcdcoXizgmAqRXQi
ctiSdJ+EpKBTf/nO55cxeDOGsZcyoIh12elmuGMiH+QD48ZT6DxeaQtqHkL9rixajmTm798g9Wpz
upmFVJ9a3ewUCALxp7gkP+3joP7ZSa0MQgG/bKGg2CY7b39Fa0bcfGJ3GX//tL0AYQD3u2UeE0CO
77sF2jIEIcolze2UeJC1l2n4mzF4ZQmOziG1FWKpSpGfv84VKfUrRYJ2evixs2b3QLMt85CYWt/W
8ss+Hf647IVVDOZg5XEu8T91SAoJVkFq29EUlNUtGKrsBsE60N+iaAtLeXhkszxcAYDMv4PlBd/I
goG4fdHkzW6YN+TsLmglBjKgcuqd539PgBbHzduLF0E+26vO2hdfTLg19vPMIzc2kROUjy4nU2rr
Gp9fbFJOL1dEmSq87wSTEnButHfU1fYM9jzoNsRxRiquQFG6Z74nD3HuaiXfU2EfzX7gBVAl+ftI
B7LY7nJbH62Ih4ZFk9xpfbSCUn/yF6Reuwe96OsdNuFTKJ/hd0CFkZFO0owc0xvSmaemKJTo5Hdj
u10MHmOW87DO8wSuF0JQkaOPaKOsPX98g3Xzf5QRNp1MqUzqgKg3jiyX16swJ+xrn8IwU4gFL01O
tKzaS/4yVisz3qnPnIKfBe3LUjGA6wz1DaEjkD1klhl2zEI51PKVcbtDT7BR3ShX/PdyZR0tsXR7
yQC4JJkEW/mbcdq3HPAaiVabio4sPRfN9ziS446lXfHGCecZByYNsOSjrkbMjnksjQznMnHZHPcI
Ehgkd4wck/1GzCb75V6WfUQBXOA7CSa99n/CSLDi99h+sC6G6jC57xeEqWKphkPEguOt431BE5Wr
YIBf9uX5aJ1SgT1rwLrJDQlRqcuTwgiAM9IiWuvLViOOpM8XnioIgKTgsLzDUJAv+f1jybocXMIU
Xw5DEQlbmiJ7uj7DdRDq0tGbXYEhylAJlZ6fNmRXDOsqZrk1LVlAZf0zXHUNgjh3Spgch+ZKWcMZ
vaSKr501iCNs4YtMeQVGjHmo/XdE3sRVu+Gk1NJrmICutJIbT3RImLY21SQs4CSYKHTuxUrYSDP2
nKG9u+/qm/nMp3q0dQ0k+ylAufP7W2mx5+Nh0ZgbesCZ+ICx0acR2Djgdzo4uYNI34GndavPmdI0
kw0rAefUemNDvSNFI75H9YRcZLCF/Ek5oKkgI+DqMqhfCr2erIYVNfytWn90Kpn81jNWwgUEO9LI
5y/CY3BiT7rxzH2C0IXh5wbKkJpm+nUqS4PRsd8QzCTmgM4KesxcRU2IL4HXNfPhTmSqLMrtyg18
6wdpMJGWtRH3zZPOOYRSvHNEBtmuhKVGYRAMDWk9J+pCDxH2KMH9mM/NkB1FUJbrjmrAEcArevaV
cEmkxmemzR3L/io4UdyjXABUsLELm2FFwxZZCq+nxbAOydXtqDst+Q6UBMdR17ARx/vCA+TiTXaP
Y0nXTpuj9+CXaYE7sfpP2VUSnLL++Tep7IuuCHI+3EAa+LK81tqCCCveStvCqpe8EglpJ45GUdMt
kxZD3Vjcg4GgJ4yKc7yEiDeny0J/yiqT5fSl7Z5eXdnwmIJsZ1gipfdo79URv3OXsKgbcI3Rablt
tS9B80Dp10wBJErl3yvnF82BhqlcE9OYo/cmBAOEeLHtMocr3jHv8pRMne91clfBUSzU6Bvoik//
/NXNRrL2nv6vDWdEr9Rp1130OfrS1MA8SbnMPpeJ7mpowDQEv++JPGXOJcasyWK68ZLOb2yCD8r1
EYSUKlhf8cQGUi6d94d26RLZNazaiFOkOzZxUKiNy2bl7V3xLxlgwmBCV5VEAuK4WSYEUs8CUZx/
hrK+hT9Jc8sgEOccdq655RQMtfFjQQw33HEsrY7QTCi2+W8D4saELMOI+lw7L4e2z9wZr5X+O5Ep
unkYL/2PlEUp4uHAXALwZtknx+k2NOQnw7VgOMARW8kFgBqiLKzUiuS6/uPw/wVeLcrUx9SFvN0b
oQgVVFwqyTkOy0WP0w37vhE0vo8+ENoP+nwjuE14I3WNwM2zOA6ml1+G4/agImY0Juuikw60XCVB
+kjXXkJ3/4H+kWN+06QNltqxvr0oAU5M/ibAgnqjWYxsC8Dwl2i7uwgHFnbrE7/1oB3FWPsbIPpy
V+P9k6iJ36du4GqHN7mmE1b5KhSJe+/cm+HF4P7w8axyrixPUiTlyxRLkNjxqmEiDxtGHbqPdbE6
ahdbLJvCKQ9tK0MJNaG/SELJgJQbWq7WIic8h8JHGH/4SGUCzavFYPLqBLqteb5LzwomBdtcVQ1k
/IRSuc964W3lKtC/JQSDUYZmG/Z+EFAk2ghKlVPc+NsLrnTWcnTfsbsCUddbhEcw/v+/GyNQPMen
Fx/bGqu6FuK72XkvDrHRcD6axE97+2r+RAH/pRzEFvtGnAgDpJsyWgiyKdM/kFHhdb7OfOuwzhi3
hJK3p+vCNnCdX0/3NnEy6cH7WgFf4A3pWWFECNatEQ5PJOhofqyjcE7PR0phzXi5/oSAW5rtgE+e
7BVGfyTOY++860OwF0AISZDpGF1bcFSkeuyCXIWNWpG95yJ2RgSGLoy9U3JKEJDfZlUbK1taXuJi
R+PTliSzSosLm7q1lnZw9KrQNitrTZYWG12msfyOfGJI0zlsyVGqfMufu8aBXOIbRa5+xJvEhRpN
EKBSZfyO7A/Uqk3VRtU62MxVJ9PCfyJkzX85rRAJ4wDjSvrSzX4zpK54VlWkRtUSTolnLIWpih1F
tXJe0/iw5DKKTg3C+Poywm2puYfk+/ibn/AKSi4/RY1vkvNePX17T7BEr+AfqXA37S9xYFtAoacD
vLwnrn4X3gmPwboq14ww+boS2Bci4Qcs9/cG0wb5aaKyiAIKZcvUHoFsH45whMcFcnBD1MNle8Ad
ZCUmzq/zsGVamS4G6kvkLjbrgz5CX/JcWmatWbiL6RGCtrjp9cEi8WoslQ4C1hsWa1SJoQOnjm8V
AzX67DIpTVn44w4iDaJrQjm5bDwTwapqec2dLDzkbI6viPfdhUp1L2m3E8Sn5may5QCdcIQPkaEO
MlzFuE+9QaxResQoFTp7zJUX8wqaAHOx2H5HcLLtQBhyASrv2jkte6GHyavqGLbvctffC4/W9ws0
VWvDavh0R8l0ZdSaF4LhHGD3LleSC5n88FEKbjRWstrlk2eXGnDUKvzpcB3NcGDRaV0PoJn6ZddT
kdP7z9g9pIl7n8UcJKlgyjD8tbL9iQXK7JlbN8MxtspcM99dczAXBw67Z8qefvp10SYa387iq4h3
7HdeOeSZG0kaF82z53R8UreM5YDyHeoM4OwHsfeOR6XZqJsl+eB3ueP4/cp7xGTJKheMcvR4pQPQ
kkXNNG3ljl2ip+f+0clhR5ICFldHGnenmxMCWU10GA03Q0vlLoziP5dWEuLuPiFapxg53YmsfItO
6d8mjryeKO0xwqOGD1oYv01A8S9xUDL4ukoZDg45NUYdFprooVq8tOZw8khLPFqbhtxTqi9djDkB
o/10hJVqeUonwg/JLyX1s1L0rM3yasjr5p0OW0ln+AqfNyLKYR9c8ViqUne7LPyIPUKH83cTFr6B
Kyms6vEGBgEsOG1bUgbGaA9WT74Sdd76gay337uq/Qe4ucr1YHLbV029pHi9ZoYAhCMiQNgGcvs5
gF/BaLQYYdZdTx7HBvFkd+fbuXG4v8e7llx7vgYRZ3pOGaP893PRKXBICZn+o87wxgzuKlP2uFog
wS0zk2iKDICuxW+WRaVPVhmsUzsJV44FCmawWjRxJyp5Fvoa0utDQwJN3JJJkauy0vcbt5cdmkhr
XQ9GlpTxqGSlmc77mGHcHZ/aAP5JO2eU/vkW8qI7ydSVSC1WcwAmq7+FoAQ0HMURL5jx23oDij5h
ZyW2LKzlziP4mk1+0ktlr5OfLCQwiiYFN8UHiTz2+3F9uPZAF+x7GY3saNSTsNjOXTgwXxniG+IO
Lf7gtQ3JnWAiR8PftC+uX67le/GOnykBcJ6UZDeE3SJgVHhtGNu2iuQsmo73AsOyeIxbIx15Py4u
N176jh8q8lVdICjNf2ZS7+bq/XZYyrGTFnZ6ppaj1JhhJJhJLmqlGHPljO3KDegGchYovgSMPqXE
VwmOmG1NL9f1UL2hrLdbEAC3SM98sGQlMe6TsIKrV0D0AUXHxKADnPOQIKfN8mKPpRIUQ9k/dB5E
DbB2FBlDa85ne2MdShvUEmkzNX+c3UUvSxd/EvWeqU6z+awxwfBs5xqVggFGGink1vdlvHDE1p/9
2MJzAjym+o8vgVkBG00VtDcHvwcs8uIOKHbmRvwvYbjK4QleR7tTOvmJqSJSPo5XhDNixOS6yAXr
vQJ77VRtqTREqHHpALvbMjAirlff1XXLr7tumcCEHII9/RtkUtCGcRHPy2XdxvqOk4Hg+uHOVtEj
3KjW0TBScMEIteqrtdFB4XRt57IdbzIuAU9+Q2nH1t8TCfC2MghAz5iOYWd0BEFy46KcRyfwDnlb
NUa0jnfLgRFu9KCry31+dd+aNNotgmUVk7VOB8ODX/1jbOKBhtNhjq0fS4p72TvA5dqtkH1WpUOo
hkZ/zLZrV+oBV8A+3iSirhBdCqE1fSBLMYcPW5x2gufx9JwfHoX2sLiOS+sOnHoV1NFxNzGP9RIs
EyFiT+ndXH0sXEWB/RvACZoRMF3exi9bdaW+gXUaN3qtsWyE11WyoRb0iF8CMgE4gj7cBNP+dF6F
IKA3PFAOj6Ya3mLCtAn8ppkqgXNTHjVHVyxQsxgnqpHBf5mzp1MulXHBJZSKtfpZy+PFdAfibOxI
z1yn9RLfvDgbo++0d6SivuQbxdZWdaTCzPlvpE9rO0qgKUfejnvQOPnacOf1Cj1LPRXmXtu/Y3VA
1X4m/A0JEnIkIq/0lKRqtBLtBo6fl2sb0lx/nYJeKIUtfqU90zApCbohrA/oirKVJSf5kq9bmdN/
tjqcTSHGm0YkEADh6DHOt9ghPiyrevNAd8boCuvss1J4jPnBUm+EEfvdVCj6Rjzb1MTUJTgBH3cn
NkTXuI1F8j9BhYVJnHrr5gcxTI+tLz0pbgwkIyIWJ2YVaQAOBX8sD9xS3mOd8HrPtZVOiRBDlPbs
/9i41Q3BNLfcYAjiBHg/fQFA6z1BaNdQrF0Jb5cDmOwJSFur69coRSQd+wfGxTfa3lPe46gPj/Ia
N8Z67iSc7ZV3bfD3rtmFL4nP6s6O7pT8lfWH2W57Ah3xUTSy/FbgdFwJ56y8QsvOnbD+XVcu+SHB
GbOxZeT9ymw1XVwaeGCgSyRv2PzsNlctORRiAb6qTQFV9ffV/NIha2YXUnU4joG/QXMN6jPWL9ic
UYEKVZqxb/adlshUBb5BsU4JgfXAA181ynVshFg3nZNmKdC0iQk1To3wqK5I1kB7W55UKjEiGk71
QNN9OZGuN1qXktARBl/JDzsY2qqNHP5zgf41raqfLm6KiWN3ZoAilcEiCdPjA35J6/uPmD0d/4PF
w3dSarT3cl9DXsW4fkLwm1yuvH+czzDoyUAp51hU+2MF3eR6jAwzGdYn4XBOCypTaN/U6pKKK5H9
BM4cGijqNi3IA82AqjVSKBToxGwiMvVjUBJ+cdjWqRNQLRrMmwY3yYvM4s1elUfkEHNUgMn7beWp
YtVGAyQcpnsQSg8jb1pB+RwRrLCQB6CpV9W6ON8BqQheGwL9+IFCQ28gRY46WvRttVu1iklaJojS
SqsyMeoXyiKPrBbdf/gdi0JL1oI/ZMGdo39f5IcOpslnq24M52pCf6/AO7Dbr10Xn/XgClPFWujN
kNW2/AiEyq+GK0hXFYa6Ng425W5Ce3aelg0iZhDS2QUWN2uGl9zmbpWCOeGwWgC1DHfM3Ei3VRK/
sfKOsQBWilvRqGhE7DFBPTT0mitmo4ZxJm0AMlLeWwVHTcWrT8Dy5DnPHgrOfUUdusY4GOlWzdap
0OADusmzw7qDWcZJ332ttCSPVMsEaPAqo0F/ecbMI0jt86PyvKfkSRsCvKqoN7rcKmK9RVWRZ9wA
iNoLd9pf0mk4g53/1gazLWlNOAippGpo4OPG6cJMBRfPhz5Ua3w6hSJDnhEXP9QpWrkv2EuRNB7N
J1mgjD4GQkw3GmFzHyX5S1+2pAAUdAPcBsJWgyFWxSp67U7XbRRBIO+AxGGkCfPpO6/eGdApX9Cb
IOQheK587BU637Fb8vdszV3IAceapeZfk46zbZFKayXuC7MEgdmeyC3VSyp1+269gu4uoG8T8cMk
Dcaf8n+ywlrmfNKlE7BhBsT/wNhSfMHYa8Tc9KXq0ydSZheQWgBUe7g1xAkSsSSC9S2jJ6e4QrUZ
IY7IjWMmmYx7Jd5HUw5egoq8WEyX4oIb08pfxmJhC1ciqZaKgV+JmvTo590vcjqGuycXQhW3KTIB
hhzNSj8oMEpcsxMFhQY5TWoOWnDIU7Yf5CwgnS6lLLmqYxsgw0L1Pq0kE19uYD22ilPDGRy9K1dS
mlfjOK5c0sEg02nFAvmyHAd4lIoY4hLLUmaE18VEhemiHGpKgWSiWpqCL2dt4erQd1LghdB8fyFL
/syE4fEKH4RLgxI55yBQ4ooiYiPqN8XMEZcr36cw+O/IYd62FIV+Lg+b7jeH1Oa9N9qLvMOOWEL/
J3zVdSy6pgBbTYxRMT/T6XPB6vkvsSQAUT0ougnBEQycmCNnB+sy/X0liQDmkm1UZUnaiI2/d9Re
CtrDEAkPt4UDLrHjBXZ8o9vtTvUDzYqMziFz64Ac93o9OuSiUOGAdAPE/KnshboHz/wlBJipW3yS
d7Fu+9lSaz6sIEazMRlr4ZD+J6X6KTxOJOTg256uND5JSULbfFEhpdgCmsDvc6gPEyDBZs4L6wTH
M6VHSrZzsAnvG+FiCYstKHroFS9yynaI146qnifzOrEP6zmTx48QLyWC7prAPRSpmnznbmtkFseh
sIhVTGrU3gArBP3F1ttfob6RQL93zNJUZU7fU3DBkgAtvzj53xDbszJkIjugAdsbNoVfe4IOj2tA
ViytNGHkwm1/Gb237zr1UhHwvT+y0kL0JK4JJZuDVc5sG+gfwSS9B14ONvu6wHFwQKBkgEcW1Dhb
Yw9mrl/tKPzyk/e2nrdJzT+QbeOAcyJXJyq4pP4BFuQj/QUZqHY6VthcGQvON7ACZuICmhTPUFZa
CltrPneOWhlDwAhzhArbQP8qPYJtwhVAV1z5HHmywM1nfppajFdaZSgE7BhUbyj44IEyyn/mHkz0
6ju3yrYROIXqSqvJWbW6u/4UNlEUNNxUiFfn0pat7zFXpkB7NPq63iJv+epAu8cyIyePPKg3a4L2
E1UyEkg8HdCvcviIMNQdUOu/ySGT4rNxW1jYs4wyujl/F4cmbFrDZXVizdrU2ti5hDESGPlAkV/H
yji1orJ9fhd5xSyUP1q+fadUcHnHyjurBCHwLiMBGhgQXbmRUjYnMb4xQhecYJSp9MDxOSXJZC5d
pVfZG4E6ogycRaJpzBS15qxS6nOqpcDsdnJ/5vqoQTgvF3HeObeR+5FEdUWb7xIS9YdjJQ149mPY
vBtSS3tEcCjkZ1kErWwEsTdy58RLrpW/vUxbnj1yqrjiTe1W8GOHJlHPk7z6S+3QYViIcU6hzbHF
4/elUZdRbowjHyXgLqYZVLL/qzJQ4DwQfsoivj935Q7aubn08J66BaJpHknVCdcAZOP3CeI5Y+Ib
DtIc7gKhu9dKAM151VDvDQ12TI3x54luDu25EVxGcVhwnct0+/rCQkymrd00A8F8K1NsyGcp9lem
NXSCqNsyblulK+cmiScbC+gweWJTPwQfBjVZiAJig/IHjZ0gPztXIjqMpE1yhOwV1wrKEJH3+eAy
23iO+qYCyM9P2bFo5Up/g6KWKrWLiB9FChRWY8eC/IfOwsPSFd18qmjtaQpFRLhwwL+Rdj1xoe/7
McLvjZVwp5zjtSwHXQoidAjQi5REENoEHa0zS0Y3sDaqEiEZqp+quA4baFw3z1dHE0XzxvL9m/j5
hb+8dFyj4d8H8rNk971bKo9h5tLJfyDncHfgtXDR0slifnaJ3Ujm4CXaVigbic8ag8JmRjpstJnK
F9bbDD+BIooMXIDAh/yLCstpUy7MVLL2Y//11+aU+mapC19rcYECuwha0KKj/QClaa/USiDPVcwT
ZeDQZ0iJsef63i53ws2QYVRcj/Sv/sR+UMz/FFYh73ioYvCmeUsOg89rgXPtD75ZVluZp4iei5DA
cZbpYmwJGyG/8MkWut2SwzrdFy1JPut12TFgQK2aX+iBtJoXas9MlLQSEOpFNx3poWgl6+/AUMHq
TKlu0l3o1I+ae62aXFmLJlqsj+vGISlsbWmozB/erQIaAa4/PFW7ziFPOSfm4VV5s+jb3b7lnA8o
uTw4Gri7R4EE+n7QxNPSAyI0IEBEYQ3XCjbgx22pMo9UHsGEvE4aHbsHaL0EzOh0JtZk0BOPsieu
c22IfgM687rs36VLUqo1j4JB7dFiF01omhRyXVjlbsFy8ecmZ5RQCZioxmkeZohrRYa3qP1OOv/i
1xRuGKcEIoiK/T+qzhF94/WWHD1UgR1PxZBn3ey2zrYSduym52vRggRQBFTFDXJP52Kz+h4YwEnZ
RxNWq8TAob4fHidLZ4jhvfaCU3nzWS5N9/WLNaD1KYNcyOM6WViZsb6kNHcXFeAVxD1IRAX53083
sdxxj7WtoIXdrbK57xTSwy/7qvZyyW9EWPncw8mHYuMoM8afehmY+nykIITM876jPbdhSb9vZkYa
6ZgO9QSHyrD/s0587wx/TpeueyGuNFyUU83sMNkCHYSepeO6DGSNOBNgkBLPeQ5Gcgd/h5dm7I/k
aWCuJ5nyO9gyQs8MMsoSFMlYHabOtPfxoq4sS3M09eAWrVDH2EHGAu/JmkgW/M0ZqDgLyJG7qcBO
n7jYzCHne1KrdqJWPE1qOsnNXnwbFeh4coYEYRZhggoz//8f9k+GOdFyl5FgU5/TIHcMPRnEMenL
LlmlJjiHzB9FkjVsPciGiTE+yDqxwAHPnDw4+NbeSsDnRGxeqmFn89jLd05VsBU54bhUHuc2wZ3s
5BXSHFwFF+NBAJtWL1AxlJI86Fo0nlkhf+qXa0l2vvBnxWROzaBj+wmdIWb/j0Ni83m6yO1d5zx8
2+y3KjPfn2V6cc+geJyttyTw36HZSy9yolsJMV2mk0ybz7zbSVLPAVXxt2TtPFeau+3yxtI6RYJr
DlEatYUe5n7YcYDlUIrMwTYPhjTwrzxUNDdgA+6yh/U2Dx9aGkdnUMdzyueUdCpsH7/kDM1vZXeE
TTlCyWno5zDPzANRYRoy/IIK1WkP1GEKuSzwdJoudkXjSTB6RlKOPr2rg112/v+vHpFAxEuV3HYv
SWSVH/2dOaXZ/T/N754HP5ZW8Mb2YHx2H+EJMnfYdy5sEo/Cj1FTa9qYC3u0QhLrqQyRoaLviVlK
FeVAVoCWwM/HFcUlMw1HO/94+St/3oLc39a+TyUr+gVobTqeY3jX8TZr8Hrz6q5Gm+Iko5n2u0w5
cMwFiOjp2A1Yhg3lRRz21p/y649FnoTNtFsn64FeETlCy7TfJb8caCNQFxZptBkcSsbyaEzSLOWd
8SqO5K2AcYpMtmO/zuRnzDxr6uFI1XGCzxfUPbnPXroIjmDjnwlSdLRzD3PWdFrDxa6FOZ7rgHRF
x0WnX8C7k40VwuCkyJOydzWaROrhkZLlXF9ulOKvfp63ALj7f4t+qND1RAbuWMxAUtsR/RB+5c2S
wvR4iYwM8zR6SoH4xfwISONtGdErtWJkgSkCTdfy5NaZZHBkkBQcvjJ7QJmRhITUVk1KQddY0pyx
jqqjhVumu8o+5e0ENNU4z22tCshJ/eAXfGNN6sH2maOXv2jnCTfgBDd1sM85B3K24ChpBes3/77z
dVUaR9dVETJynlyGD3QJPGkxVKRQfWb6NmIBtUc/q8swKZsMrR81uF+2z2GnkmUtIrZomCIVOtPa
/3UVb06q0TZt5HMDJvh+FsAzkzrRPd8iOKS7XvaI2kI3ZTeB10RyuXLblSsLK7hQlWRHpSgkYCbR
yueS0+NvYaARFZ8agcQBAyXs55tBme/EyW6Jb7JY/APfeWpKoxGDV6bf+1+rrGGazMpqZ4gcbfvp
kCh6zH0AJTBLHiWmzt5pVyA3diT0ejZfeEend9G0zXGPodHLVMw6bcn/WXVREw8/KGR023f6jC6o
jXm0n2WqYr2WWwaJGSJuy88RdidBrejZYQv5WefqpYCh32G1gtnC2baIgfchjdtdsBA/4cOfG6JN
18jjWpekdxSZeJ0ip0ss3cyD80oVXrAbuM0zJMoEeSUu7JYD9DFM93/RYQWJKjFXH9HvJQDp7frH
pu1+1jIC2QcgD+KYWYgmZ4GOUMqkeLn93u4+ujWGQm34LCjY/juB1pVigHoTkTsnrS9VyMcLfJM7
83Td/TWdPjHoolU9apqzDlD0wBsEQqTyz2MS9mpG46hfUSJ451lCi6RuuPYeXFmrDQDw7DSOiQIC
dzAYfjWnHTT3AP7L/E2HfRNRib60wpU6cHmpia4UdRXtT3499hXFdM9Jc5i1443q/pkTlrkx9xVb
SniIEuoKMB4A8fCkkkueacUeYTsnYKUQUplClrqDlTP7fqzQwQm27y1uAyufC17rNh9L6qztdemK
79Ra5cLGSWBzbA1zniTy3L9KvwgodyoUK8Qx6JATqN98jtQtYE15qnDM3JIpYLM1VrBKgDrQHb6z
XlQ0ukhCE9Q/AfuGiAA1i59TYn2If6smqnFmDq4QkaMMvRXGbVPE0cXek8uT4rGGQgLCTpdBeHx5
sVmWrg0Z99GQ+hjz/vgY5koY3nWw8kHv7JnTSLvyezTnyV+0arx+QW5JBVQYQZY2TSgeZQG+UqOH
WU95WiiI/guDmOxj9fCBdHO8phVTr7zLocJxzmYclKPTSj1tb8QmFGzu9fm2XPOWop8+kRrbcjL/
5MT6SV1XXcMfLCZKf3L4Jxnv1eB0JaKzWbSb1FqPwDXE3SJcmy4p/ldJKD6SpbGec3BQT1bFh4Hs
K4msmfxN5IyZA1JXMwnlyYGBvQ+xxbDRTNaeUT8T3AJj1hyEV8ip2itvfuvMXngfZzIBA0NGiTXn
M5J9nSGFjIdnyEqF+lQ8DcPeZ3uamhx3mrcewkomSQqpjP1jlwutbBQNEgFy3K1wsZB3DR2Z0q16
Z/fHJ5ht1N6CPQV0Neeo+wzNrxaoHDJQyrBd8I57O15oabJcae4aR/ERoQmlQwWSGqgaIAj141V8
1yYB/mdVpy3rB7WS52W2T9CzbbcNqiQ1/m0l+EmhILoepa2NCat6PUZyIuOmP5DeStLAr+NIrxBK
yOHWQGjwy5Y04S5UBnLDjXR2o5pjeSlrpLmIPE6zC7PkcFUPzNKQiHQIHy5+vPCGCfbjs2HefrjK
rtBs8wfaA+HaYlbXaAtZYbevkrI+xtl06FdAcD2zNw+Esh0B/PCpRjgKkx0eHpbFRVjcoaFjulvW
7l8nazwbPu1sWHUGl8ILq6XnCfGoGRTZez7sUs90fzvaT+crtF0G1UVPq/IBfrIHLtDNyOUzUrc0
i5lqAJOCxvfG1dd2jflbkktqKZxq6yUtgAXQmVhl7S+ZXpZX9Rz/HwVPtD6277wAnl2OIEQkBUiZ
SvI8mfcgePCGB6M7TdivyVpoxpnm1uefNmGSqjn1RC3wvT6ZAmpfIjZWTdH7mzXAoOVf409OBfnw
53nv7eq5uQ9ONK0gOfp5um6nRKo5UWD5s6qB/oH8rS9ehBnTVHt3dRNFy2bmvfL7fBINRRgEjA38
OCIKKvl8xIg7UCIA2XGZJEz6Cn5aniyxWZCr5z+oYXxd/macpAuwV3HuFlireP921IQIaUZV+oFB
3xDTVD/GjlIN97PT6SWfAj+PGNF0ZQ/DC8ApW86aEb7Gy6BUrOKbcGqxi1O2zku+18zTePgMU1s5
9hR58hzbp7E8FR5OzABsRgeOqf9iVgE5VooCPeQ1yKgLto6GOCUueHa7OD3uoDqmOT+yeskJY0Oh
tFt8yzxBVSjRnX27GPsDX79V+tmxt9M+PJmZI0jaUl0xIoASKMTYDiJ6lD437XDcsOex3yeTcubq
KT1ukUnI05UqgRf/FgAgFQFZDFQvCSz1kpaiiCBH7pwnfaQ0D/r+kPklgrDIxV6ZjEAJAq3NZjH9
jewio69auH4pvIUZQq8lIuVQ9Qn6EXe37bqWk841s7LeZgN44kx06FwGyb1LZgGFrsq/xhtbliws
GHQ4fqcwcE6xgFQKjuzNft3+LYyq3WpmM+6P181aR40kyWY+Lc8bm6FVw7eWqdZYg9PcgRMmS7y3
MXCDZkvJVKlQ6+aYJTbJzuqMaC6VbjWVj/ZDcj2gEMLeFGin4xt3uzXYIrcNOYWA9UMMSHkER2Eu
IMmr7taGWYqY5NBFMcUPjfnXgkpNUA+FfvsxFAZ40HdHbzj0uOEeujFVhF+ZvxFBw/uBw6TiUXN7
raDsQpAyaPO6tDljnX8JSIqVE6thM3TKOhwK8jH0pxYhxKeg7Pbkq2XBInWLm2m55d7/KFgoIXdU
HOyQA2UOoDKSPJmn1HwrGXN0wVoq4L0gcBBk4L+ozbbHIu4vpxl2fGORr31U7iNvTUr+ZdzbStVl
rL2n3p47aLFyZEnvqpzoE8cSkL+8nU66bCuOE5Ap74EUWsz3zqZcHWWd1ko5NE/U+S6rdFKw5IJe
BllX9iyjSDzuLJ74kTNvPi1ahSztmtzfYb1nT8a9LSjCZ40CWhd0MP8nQZUYWTsNzTz6rKKgUg21
IxTX7xfVINZ7J1WhdlwwirfOe+pRY9ISeHJMfu5jRap0r2Ms6eigZRrTqVidtMQEboNu8z1rn2zX
qnHjV4GVxDkqHoV7VdcTP1TY51r6aOTWpz1e0pV07corE7zCgp3/7ZNCCy3+PDGo5Y07cdzw3ABN
CslHWLbT/qR6/lMG1CE+ZXRxT8/WutmXuZ4OsQpelnmu60iTRHNFS0MvfGMUHYmGYmLeE2/x3Cu2
jP1JYPbXa4C+ZlV+AtLY85GyWH6PJgTJUdX9KnVKrnS9ZlBgGj8L6KJIaewsEywdbUwqLIOxnTO0
EIDyxV7+wMOP57hq0Ei3kKueDVBDw2i30RZ0VZUihilZ5hhsOQeHcHRK9I+rl7OTgPMaECqMnPP1
1/9ivkXFtBfvwwcOWGoSbKoyesAbAnd9Kq+c6RoNY1vsdTFS5GhYugvn7MB9x1AeA7eGiwSscyMf
jE3ttPOfL2vVzQqn49iMsHnnNrSsb3BOvr3RHQOuumQTGlqeHPvY2Xr8g0Pt5dKSpbQI8we1r6IQ
tDTfRZ2iQwJNokC1u93RQK9VMjO7i5UItDh4l30sH878xF0qzRtbf6a0DeoEOn9UnCItUF4Xos+6
S4rsq9ON3AbgAkARerjw8Az3FU65ZaB7V6c1Xh9ktuphVGlXx65jni+xS8HGpdUUoBdEl2l6l97X
N+bPXmjltWApICeVOTjGRWEw7h/XDkovzK+W1nveFoIP0YHy7V6DaI6bdPkK6cnSUwGpxW0iH+4g
XlZMV9RM1Tt87CQP4xuIePU8DKF+7LMINlYwRequ+Uf6M7CeDGhMmm00yTWSr97+t5bmPw5iwwGJ
0yGxuPtNhm1AIJJyY5RDQFERwIG1bnMwBtLg7BU/48F9/skUO6usHz+j+LoAalEOUbBTGsyLkiBh
g+6MIZwJDvny0Y8kiJVnuR1SSa8zP7aSP5VOHntYGnIeshbZl6HD8Y1zq6a8y4Cr54ZMXTNfJ3n2
hhlTXUjKWIxe/LZJoAIeUc1rAmu/cf6hmL/KIN0/mJsgVajN2B0mBtLXZzXwO3lb2EhwcJEr624J
0ErmTO5y1glmzkmzhGK50eVHpUxtJ8IOsVg2tH/PY2ggeA+yP9JOAbFJPVMnnG5Y+mLr9Fbx1Fjk
usmmuYThORn0xF7VdbU3aCGl/GQmp/9CmmqYZ1oP4Xgs8BQPWcw3Cog5Edkjv7D/DLEHwdS0do7w
ULZ3RENNVGqaqw576S+PS+48Z+I6DexUWMP1rS3ni/hN7c9/LVBGWbYTaO5s4dw5kDvjziYpXXES
to9pYs7TaIOq+/oXhkB1xmK+oelPTrrlVgLsxik+gu5sb3fd1urOqnlqm63dkN/ZAyO6cQvrSEcY
obyXzA7JegA2nsZecXLzQ7FKcY+SxjrzDYrj4yZn33zyzNmJ9QGD8xWanA9Mvfs0t1+uZ5h2p97o
4GObBoY62eC0iV9e3sWbMPrpHZzhpkebF8kJIbYoYh1zHBW9UU3NAMjzJ6Z3qrZvzQZSbDANmk4P
ALyBdCg0tstK/kmAvqYNUr7jWSmgoUrfZkywJuAR2+7GllCy0W+OTAomdWjfW/0wwaEJfPVJrSLK
mUKbvq3goGdin/ZD8DzBVABThhHp65KsBWHqj9EKEEKCzCmd/TMBRb41l6kOhvSpL6q/qxd7HN3O
0fV0f5GMvvdI27O9DumjynBJpl+FrtriUX6X4elrs40Msdul01LfpTFNxZoPwocs0ScndsMeelkk
u1RddjbW1PS5CyvIBXuj/qhqKiYwsfUhFDdyej2mc63LoHYuxJbxy5J7LyvRePGnTTm5i7daAp45
+zgl1xHtsztibzXyHZMVygknxawGe8wh0GlcD1lNWEvzqPLL9fj4c+mR7JtRqiYvYourypbSzKvH
uYFLsVB7Nz8sshG2ne6TOkcK4Idus26Dvs/ZprPtNi/ECo0/6Iw9IBCflt1KoeOmhm8hujuQCJcE
Z9biR6PyxUDA9PBUizfCZN4mwKFL0exXi1nyOdYezDDMcGkMX5AbR2T/yX/qOBPpEMflpgpzABqf
wwoLRfAVICzSzRF6GOWUzV6rWdXxLESBUl18kL0rAh/4zZOu8pTXfxVf0dvPRZE2jyptQE5CJsg1
sICmYUu5LkFJkno1kcUEEA3cBB+QDa7b+6k3mdTlMIEV5uAOCU0tu08NI+WcY3l/yjnJen3zWn5A
LYG+V+zAiRUT6wA1KYx1duIJzYztgjP5WfN0N+WEUT0C7d68I3MImB39Z4zWPrOb0cvO9myWywzn
p88uynsu/m1wT0Z9agxB63XHy57909Oc+23n58Z83uDI6B32NeCtxWaiFiygxnVLOUup/fgzyyC3
II5H6kA+xUG5rtL0FMK1urgPU550MN4qevLTsmOzAp3Aye+nK2YZdM9GCf2LcmPOY5ZbFSW3QE9C
iPwTnuQTxjYsjMoi6LbfPMIgjkJaMulU2t1bnMgkANc9g+cOBEJZiB86T2t4VUKw4v7tLjAL+3iF
sbw5KyZpoHCSnhy/JnVrMDnb13kIb5n6i32NIbc/Z7xwg3Z0oKLamuRl2ij9xiF//AAYR99BQ2E0
crewMQbJuWBQ3QcWkGYkD54uAL8xjSdueAYDWqHnZZnB3097qegIekklNDxuzymIGDUz9wsXa3k5
lL3go+mCmCYVQTBwwtQmmEtmoZBaejQQ8D8vphUM4FegWXHT18hVSKjLKkgoJ35nDwIgnVKiAgYj
eYpdn2Z13sGDlKN122QXtBiWAPxa1TD9jPzifuPMq0/BUV6vOWm/IiLk7rH2XeOPAr27AB03+SHd
9wenu1br1L4CGvpt8gUmL35p9PFHv/qCndWhxEMfwfyWopbGx1FWRrIkOh3eUQY+q87nEINHFQF7
ZPzSUwTDKgHcwKP+8QXSyMMN/twnnIPU15xXTqiDLvTl3UjmS7Z3KUtcIk1g58bB2V0cTF6c1a1+
d6e6puZnwTk9y/DSc3O3hxQ4FOEf9elrlPUPtQzr2yuvqstPTCavs+/QT8hXQdimKNwZWCVu5iCO
+VTn90w1JcDTq8fqhlBa6YGTJ9GDXMX7jsMxoWFePkNxx5SyqqNosBZksNJXH437LvbHWNHBe4OV
E7i7NiQbgdsUQQQ1JfmYaUPTuM4hC1zb5mP3pa3PFC7RdUa/NkEXPti6Ycop07q2aj+aJ7FjAgij
Gd9RbkQd24/1EJy9eyTg8wH2bk1TjKRZgza8z2FrkV9hIfBLxa1AaqAhvpfqiJgtVVXN86x7iqSH
rwtPEHEGBuFOA9XVkLMzPcxWBSOobRlLRfkrGVxJW9OAUrlHMpK3JeJmcfpd4PhaVANVFUT8z+jw
pt0Cc015C9SyqvzUV4UqdHmk+fvkpC61Jg4v6xnH1LcTCjKf4jSh0vwRSVnApemsvQFNZZ1citAI
SPfzW+kIe+Ml5Y1XY4BtQ8HPnzYizlTa2H9ZDEQvvqAvFPwF6Z2ZROgGaONn0CrweDgbrH0IAzmb
BHJMcBoqPuc0s8D37zTKTBS/etD4U2pY03tf+q7xs6PNhvWSeiH40lDTAEPIUX0Ae5ecrB0jFOdQ
nOi/gI5Yd4ypVg/4U+U4HlIPOyn06mOR0W+w2Wx6XgBRBuu1JloJII2D7J/VRKmLir80hJFr4J5B
64T+Ofodi3gID6r410aJE8QOhdq+Z6cnqt2YCo/uWUHW01i9cwttWwcqp5yVcIPVOJJEaB4SDpkD
AmjLmfMY+zjxI95tTqIova9a6KWyp/iaPnPxiUvhiMhkLletuVKsA2Wd4iah19MPheA/UEMLpyWZ
SBernZRfvt/gNPgrgWMIBGdufPUOi9mIdQ9riMQB2DRJb7WVOmWt3u5hoILgHD0CgWKUZ7FtJa7/
3AfKbY/BMK+AAtK3ufQWvqFkTp69zOJZIUXUK86Y1MzfL6G2tVgW9AKJlwUpO7jBX+TaJ4WcU9Bl
V+qbsW7LmFiOtYY7ljwIlx6cHn+QaUu/YrS7XO4BavWGZeFPJV3mnHFPPzoPsN0WChGSHv/ZJWvN
//eKtr4HJgj19aBfdxoeu4svA/W1VoEE02MglP6yrU4f+5SlIJ9F51A53wG2S7M28sRELJKXoLBt
f2NFHxuq17h2MNPuAJjXnWPPp6dna3b9fXd5XUSjFvo1JpZIB+dD04EW3bLKs44e0s/n6Nz8A2MG
7Q6IthtvL/1YApxr4tNeX1lCvPoX6QSVzGWjy9dGdWLqzM+hN12VmtvcIJVU7NiPEm/cCp5fMN2Q
EVlWzLuzDHF7Ln7vCXMPwD9CFBARfDW1xPI2+25BOqYaNi6KAqjPBln8+WPbAASwehtY9jubG59i
lg6gmV+Rky0Ns9mszIhqNYW79KrJo0jphql6IIG0ej2tucinUGo/n6rTT9SvhlvLqYcbqzrrTibG
gWXmC1XWNwGdljak5X757VYZ3Kki+g+4nFa0SzY19kqmQChv+Y5v8tCbp6kWNQkatJL6c5ndOV9p
IhK/s2rU1Kmvsu78YMoaGMLtdhdUoRsNKCEoiZBuhQiA0duL6yorDp2G2FxmdYhQitIAH+C0sLNy
bjiRcztcEipCAmwK/eLoUquhgn7fk1aCgftdDNj0ISntbgSDFaUCEimpJq7FMiZwIykSUV6YBbjH
Wi7WuGWx83yPD6r+Ga/kLXIHEv8qM0NmOwGZub/THy9E4tyxvC17IN7+j1Ye9962o+3r116++iXN
HwpahaHQRo5dmjwJB4v73WR98raB6CAJvRGyFZTRPNSKfc3mdEo8AWX+DmrvqPiPdr1BvNSbBCj1
+76j9KiJIzaxYC/BMvSri3AZtKou4Y2YVmXE375CDTHHLnOGN6dwXGBmOUoRdrvpQA3GZgaUdy5d
nsWirzHBobiDSoOqACRpyKp2ldWA4PIZKmsMU2bcoA5Pg4tWWXLxMri0VTHNbMFPPnkDeKby/I/X
OLHMAhDG9JJXUOEk57R2LRu6fM+QIF084NGrW0oAlHKgea4NsE80d5wkN6DRiUZOOaXeYrXLhh2C
LaJJgaOv9XTzjo26RbTO0l9ldnPpfDDVdzuMe5s9oktrRnKD6tORBKMeVvCix5RmvnyuTT082Hks
FOEcZJ8MS9QUHz6ax7JhN8cm0R3ZfdxmT30ItA3rEVPBvvekGHIxTsj0ICXXvivcCOtayXUkdF4+
mGQZlAT99GUKaqkn7NVaO85WXxmu6bq9Ok2UTLo8Hf1WysIaF+pEWxWVsg5V1PwI0LcaRDF2KsWq
ERMl69oZGzRHb7yz4umEVb0R1QWzxE1lQQxajqPzCassHVvhBcP0sCVNvaV4S3c8neEj41a5sdyn
Npke/AUwRjHZ84mDFPLA9P3PTLFROA51R2pqKx/fHvN0/XHLLaWGrtYn4JMgTFYh3j7SMG1O5ENT
z6HxGw+oyonXiMq/nTYr1lM9c0JKXS8hfx2KajUUKCj7fA7yvCj+tW73rmz6PTwktOvt+JxkutRb
ZUpdK+hLBVJV9l+6HnGOcwB80a1OMIZwicEAWRWHwOMSNNrFavwbGmweODmJG/MQWR7rKe+iuye6
AzX8okLA+fnINzlFcvy21tyA1sY3zILXiTBoCnierFZRO343vR8AKbCeNKtxDRiyth3IjF3Aq95I
EIG20UkQJqEIrnE07/QtJUARiq3DxNZKLlw0ewKwV/TVu9xb3cQQqSbuHHFVfbpoPDyiTwRxretr
lOmYreY5kcPVdjXk29jxAAYsfTPEXwFs4ATr6Q+uGkXXA1FECLIrCcJSk5E4Fdxy5YJUS/8ycQjR
QvBRqw/lKvhQVy0VjUAeVLYWB/PRtAxQQZcchseH+kyquc2toe1YoI4+P/MINMDpRekDgDLvIAHl
semV2QdWLOMOLts2y95D0nQ+PhVYGbzrJijjzDricopsjSK8ywOf14Qu0GPIkGUUtF5OCO3Ag1XH
3ln14LIjGcvpcdUwkcJz+i2QwYAVPAJHMNa1O9R4UeKqs2CtXgZnhQj4HGiPW4LLLycsIM+EshT/
2qlMcNrjiU74MS/WkBR2KHtEqHw9pmMcjRQmPfttkk8HvcTXpGwOM9guWpRQQUOZqJrZL0FZgveH
NUSLwKdM4NPQuKFKc9gmPIXkp0d8vgDdi33mJJl+KCyU1X0xvsiv9c/Nk4yHX1uiFyOB3SS4qpM9
/yAHZjX8qp0cJksR04DNFZJQAP39gyYtImS5VXkCE3dpfro2MyhQV+oLBsioI87p3s/5ZrqquDbl
7PVEJxHUjuHLXgdGGN3tGR/nHpWjtWMjCnaPS67DkBH1mC8a1Fg5y7U4ATu1pJ4GjbGeBw0jnQT7
+glv4vkqsgm5KwRzjAB1M2AvaYv9dkjngjXN0Sxxsiei5ic5qcO2xRVrVQy9CP/UAAgVMsEVQcL6
qbRrIxdyFyOSEoORxME1tN3m1mLV6Nf1fTNTsd4OovXUJ4OVzJ6d95WRcEcpPzHszK7lQmu4Tf85
Kq/Yvvq1kRWVU4UXA+SYqSL9zxJcWxxV0b8iskkDcSy4nFIADc4wDfwdu2bPZYz52uvhnN7+WeIE
+KnI/f9+2sefKRzHt+yPvj4tSqAhhpNVvBeZwPiUZAs97aidec9Tj7ova0xTqI7tOuBlwXsPXQHF
gZgdAzvivDSLS+wOH78ORq46cZC7ROUss9rd0jnLOtqzgz0eZOHj0dJ3O2sePvRxokAO07LzZ2oV
OnSB7MmP2CSULIkIob+n7UFc92WC68BNaqPvMu0i+ob2/M2r+N0zsvKUW3/PvqexpAGcsw/w6u/u
YMNI8+r/v1Lc0nRzyBJGNqGnpX9SQ2YY1lsnkt/RCcyo19cO2B48qtKdP8cuq97sQq7tO4/JSnBX
y82BeykPHAGIUTp06ElqhoCsG7DBoRrA8o5PQT6VmcapNMG/IKQ3/OAYQCDKYpB6cJsoS8rcK9IZ
KFxHnfpWYSvSM9Le8fW3FrNHKsbApmgpbsW588HOkL2W2zqNUVtgfd1XXIS7pTL1Aw1LO9/qKK8q
x3L3cdQx3zwOE9OVzZ4GZY23KReEpCgbmMOXLnjkc9f+bmuw0UJsEcCQG5teA9oZYi9cEgJzVITG
5zTOyJukzqKrtahZ9mOMPVX4xOIDFROUD3e+7f37F5xxjdx8vVMmeR4ra5OePlCj0B9PZbFmTdbH
W8hxg1p3bgKRwUEsWc3Stw5nKjk3OYJOoV3lynxT4WSvs+caqP6gn7kXRf7QX/YI9Mem4YwBt3Lj
rkPzAQNwDIH8pN2T6LTGbQXLZYZ1LkiENACF0ALk5HyMr0PR2nwkEkVvUPc16VFZrTa7j9g348nb
KDM0uXEjs3Z5iM70XF2SQP7YFFWHpNx8yajhVYiQyQn3w6PLwWER7ktyjIH0PlOwtfu32nsC+DXy
iOmf+p4zaEyGafY9f7fNEEJXMxeM4RpwiNgKTBEqmr5TqF5EiU6fFLK2NFMS1EIZQKM/cWV9ODRL
MmjWm6mouxhxFNFULyyzrsk7VqcEIGR5UxHBCIxDfwNkVNPb/QnWKerZ19zFVsEZODViGng1y+Ry
TqdIK+8Ek91cx8P/C8PpC+O+aSoRU/F3ISVinq/8X002uRGFR1seH+LRMJwPcdqKCL3OL6sMEfDc
Syt0bxgN/dAzOwZC43J4Vgk8KxRirVwFe/PizbJtWikg9GdbTD5RR4VnSykR1OR34YBLtca3q6pm
6nEXRIl1igTnROhzQuJvwUtnHF0OC9YV7lW8W0GkGm5tYIKHNMOC43MdAKRNjT+CAFwhMTC5uNka
bNiaSVrtfWVzlo159taU5bX92bkEVIT6vnPYhK5754gEw/h47PCc6IiTJB3AxRvUDTP1qWJW85bn
X6g4kTl/LUh0b02q2fBCmhsW5NgiLBHmHFFXvSOQRcTBtsGIKtPX9Lgx/PkGKUaB9zcPBwc3huqa
mhVZioQUIjhGGrXXUCCy1E6w782d/O6FcAD1t7/11DTyzP7V8Yz79ck7r3TkiHUKFVnIO0FfJTrP
Z/sg0r9gL1C8I/J8p6BJHKYyx0/ogPy9TrCK3Yp/IJ4IPzMDRDrwRmYe+eCRLga8c6RRZyrjKHqw
6XhXZXIrJvOr7eBk3zevU4CBOf/luGMZFylDNH8MEsbYeI3nGfkVb9OMQIhXFVvi40SqgpAAT1IT
Opxx+64BgRIN8L5KtQ7UJnQp7NafcvtgPAuTKuue50s2Mbbpzz/Iowq7dgT8Ym7Y/sYNxamahbvm
ynAvqP02mUnnaTdoqPd4RI+Uk23Rizf455TBh4BmGhrHEkbcT55N25D7PZVbGXpjwTswFb5z626/
N+5DHFkRLChlgyijpILKRf0QMiYyzBi2jGhf+bd0qmfQfY1QWX4xmtYX2RnY+IvWRgvcBeaPTvXD
EOTWSXAL+8phaOTJ0zBCpfQo+KKLXmN1+kFX1xEVIwGhWiSeFfK1lQaI3Gbl98SIBWIYFE2rBkLA
sYVvleXu65MP1hVm4BQcC78Qco/B3I8wlWsMl7uUy7gEonYFQ4sH0roumm8JI0O8EdMq6nxHVgOv
DyW8ZkrTstJhGIjCB7MFkdN212IzyofahMs+zO68hsSyjiGOqzXF2f39wszLgGge+KTQyTEGfanJ
lfS3Z1c/ShRwXhncDnxiRFKl3Lgx78tBHNul1LvKIScwuReAumRCWcj1v83oC8fiY6X5h/VYqz9I
WINhVBEt3cwrsDdgqxVTgxL7qsYICG23AThcGMtdTLQYGLtYVN3xBmrb+4vZCEVMHi1FGkm6gXI9
nUmspBNLkJKlwCq+8M1wycsnsFkMTfoASrwWk3VsXjjX4lMd5K/8owNZmFB193akNarAkIfH4eME
qpDopHW58Oz5coI1lCChoYDrz0XerW3Cn2Bk8Reba2k0TbNkKdToaEKMhoAJLLfsCOxVpDIDfEhv
Cc+aFoJE/9r85G4n05H8DgW3OUt/5HcIsv7GWxuIj/rYa1y6E6RXqpV5SzZcu8wMAfe/aY2ChjB/
mnX/5f8Ux0b07fgUjAEkFKQPk4/9t1peFWUg1Rg/vTYEEa/XC2GRLv5X3kU5n5MzSeEnpL89T8pL
6YIHJXqeUENz1a7JZozOINp/htNbllHWfGMxysYYHqxhQ8czy0cLEloqVRk4+joPmIHY1uhrEr9W
ZLMz+e7t4bG4YshFz3RdxiUATZPafOIpGm6xYzJAONtiEa8yVAo37wLBR4pgXmkg63c0jVD8f0/D
M/oV2szpuB1S4Dj/wdymvuGf+4Mv/luyiGiU7+hwJNzsi0WHnEwhRFeAAngd0OolGnYeWrBmJN4Y
eUx9Cf/hOZk3AhQEUa21PISeNP0d2WTXrMk1oJVBFWr8Ao8mEiLiQLyZZcEfdY+x/SFeSg9M3lYx
sYtQh6+iiwcavNikAYXwDcvZymNLoZwtilWKWnN6NB2GL+XV6FGYa9YTxfnLOOxLzu3V2HdyIgsk
cJ2B0hXVxdbgU7JLHQxO9B+e0+42m8IYHtRwFuFi3qBkf9RL1DV5KjEczew8aJT9Nm8QVXyrrVIW
azs2MRgwtjDos50NwIaMk26LKpl24Lk7MmnXuRIyIsyca/q4jEQCpTRyyF0Z/ngQQbs0XHRBk/zj
SmiZ519Gvpdsq2PLz5bVRrj1oi0a27AaK80GBLlrjqY4FhY9JXmYMmiDNxYwZlsmXIgBeo4vcY8n
nDBlblXDBGpz6CPJXgb0Fgvyp++lbjOAy1JS8+YkUFscVxUmtz6p1WSVG4NeZ4MTP6PRkN1ALRxf
l5AFTA6XlHFHEpH40XWBGgTGXc5jCe0HlUsgMSJchd0P8ENTmgx7QED63QA5VB7bfMp/ksQKUgoS
sFjEjtuCfItae2mA9aimhxIA13mE8tNKfgDW4gIZcgY500wSbNutA7nHH5mYvSd6ameOzHxtkw6i
lRU7l2fvrWML144y5GX8uR/eWZ3N/rQhEeNFM/fVuVAfYBRa8cuGvJktcjq9Id+Vn2zNCp9AT46X
Xo2rKeEEpwC7WsCC+ZYzOjvn5c6Jv1rizAXudpvyQXsPtLQj9eYCR2hRcWRShmpPR/UA1p/Uli3L
2yvoqIO53GS+FjJr4z5Yp06h8dmTZp6VbYsV/tKyDbPYoKZSZUFTZEFdFXT+N3QsEy80eGEjDI9w
AUvYNtDxf+3y81V0IjiF41h73mozHhjqoS16/f3704zpz+egDNv6mPxArfVT4LlDmHGM/auEeBrO
n4XtuIxQ94v2JgZmLTxCa1kHk3SbOaZMZGDDjBmfJDrD/9Ii16WD4oNzfoGRLeR1FQkoaOmTkc/j
iRSDs9L6jliYDGINo4zcR9uYcECNQS5Wn5EbOJHMZtJ07dnXOqgoP3dnCRGxnQoqBSWSMZNqeER/
Nzus9zPH6ogWgsyAuYyQ6Jn3yIUUWzdf3aZO9E++mWQdrftAfxo76tI/Qr0nZA+7QhWCzTMqR2lt
W4CiCr0GxNDYHAmnwmr1IIiLx+XLtADOicHODTIMFKP/csaDX+WqHNBN57b3IHNruG7bzLqjfmBR
UtLo+u40WC9yA/prwsZWEdx77ro7KXRT9pzY2Qb+AfsQrYssaiVqqygX4pNkedS9hDPzK8fhNRdu
XHB3akNnjNPxHyigqVdtOznqUHO6PG7wwpS6Z6R3gMFCh2yCPBdiYPCIQOphFwZdYi/pe1W5o/ER
N2MMZGMmnK1l94uDh6GQGjOF3o3tcUiGurd4ZzhEzBBUgl5Nq0MLnA861MnX85vR7mKVdFrHNYmg
0U//58BAS9qVM62dmWu7Jir4uc9L9VNckXwVPygBlkR8jFL1CEGuDTdB8gVzZlO96QGc/QdS9LSl
Up7ORJ+T3AKWTMhWHIpvgY1K5miSIU7hJFpHu0GcJmwUBD0Fs6biudglhcS4LGq4f+/jqBPH/vqF
ZGmfIupowwpNDPz6Q1fHB4kh3vS0ZY5YC5CM2VJ/lFQyh0oRanhCrRho6Phl6pYer9oIBVPNz+zb
8SysGGycEG+PsB/9uUNldql5XCsmP0WCQ8MSJ0NlTdrMdO+vTib1CL10gpBxnecgU2ixlkT4Crbz
Oryfrirp1gYD+87gtGXdqADWjAMtyjO7UzYX6lkDvNNrtreJAgtL/5Si0ypQOb5WZEQ8Z/oVN7iM
w8/pjrWdxs9la8o0O5TlsB4WAbKYNXXsxrpmiOuVSObXYefm/UYHdxEjfOqIxGIOwr4RaJ/twmzS
2zlTcUrCoP/gnvYIiCLdRj5f/I3qrPuBZSkubMFyvZg1sdZ4zUkMvAd9oodH5GTw8Z4LEL9FTsog
O6jPdOkSczbDCPwMzftOY4VioYwU18VbLVbfRV8ff/1HcX8a0x7p4Eod/dzYOnXwjkStue1AVOK9
W+kmnZZK2LRzZ1nAgHFUOndnjH+vrqaO0q2sUvrr9KiBQmSXOwFs29aeaJLoXq5b61tPdtQZPqzN
T+XZu5SvmJddJfNn6I9SC2zECHAP4IPDpbtgvzgKrxAMzES98g7DIwixEkZJMQQLxXP+Z6RjzNTZ
hrKfvtagntEYysgUwD9wfYpiJDi1FEn6nHLQhfjoHDJy5JQ/4wHg0P5t25pgTSvrVcHXKpa5j5EE
Lr6FnxwM7qJ9jiEtvLoWfBqFbhSMRRT5BXZyL3/eC0nw1UQnE4IzKHDybBhP7XZI64J+E0WNfHJX
KuCiFm4KLsXBOOgbsZER5CsAdU4vY+gLSfXO6mYlGejz5rAWw+I0ledbDAeo3kX9E5solTSU1rlF
cgXhDRcWrKc060didSLHLsJZJNwTk+NHgRFiVQ25BBWLVKiLkiuL0ETxaFVLKAdVlPLRCMPgJ7KT
OEXlSInv5fvlmFMWu4zAxebNrxdnKu44KO5hYuhH4TlBvUTI0k6XwFbDwyen5WnOwVoS/hvnRdxY
Q8qcLP63ofMb4WheL5t+FcVHqLmnXnls6dKapzk78YhPV8j41j4WoyTfuhKfxt+y+k/0y0Drdg8Q
zNlk4KF/gRXwiqopYj/yFmnlxpzfrLqlyeQSyha2AVZdo0J3uG5vhr+g+nH9T8aMPjhqI9guXHKJ
u6/3hSOMGOtfTOstCAohvZdZYTbOvzyiMqpHVtQi4K4uVv64Ny2ilUqKxz5d3i4vUot7cDOyU9rE
OL/jllgrQvbtW70qyzWs4HdeJ55DGUWpWPDD0DMTImLfjTYuHTeDAZpF6sKNs6Cki3CYjmtYr6HE
6T0zgYq1whzECHy9/Pn0DZjFUmKBOxzbimXQFjES3ObhZA2bG23XvV8BpVlQsJXfSX0r9AbZI7XT
/7kKyGnbnzJ/ixmduoE/w+FQbkAkXZF0IBrpOkVx58kUBgA/cPTOzGuikBe1ImLGUfvFSrzO7Kfg
0EwegW/QHZQAvkUZAHa0Gw+LFUCvoza0t1KnBoQRWWQFlrVENGDGSuygV4m0u5nWHmSV0rmnax4+
cLnofv0pG0oX2ZK1xVUFKFKQWOV6WTUN/8GNAfZD0z8nZX413aeLyIwe4sT+39MS8x7avSjHOupJ
rg5lEMfabxjKuYMZCmAKiPNIdqGZ9wtlLbzhjmw+i5NYvi/11TNQVclEt+wphCEYCGLGv2J2RBjV
arDv5Yh8Ls4pI1mo3I8j1cPj5E2f6WJk9qftjDBivFy/WF/hztgrYc+I4glYJZfXroZdj+Ze+8ST
LPmo30+EpUsY6HjiZvi7oQn035FrM+1CDzsK8WzCWoBCA/f7r6qtOfazGRqRU0mPEpQieBk2cjyu
b5F6NqoONAdiMTijkcKojKSEfEkIFKi4CdpDm5jn+IGOODh1YHR1SnDD+Cma9MDKsr0wSflGsZnD
3G6bM/QlXgAE0LaV7qZpRtTsnLorDsscvRhpEHs8IFTfIPR9zUQtNn+PjldPb6LwwoHD+PZnib73
au8WoEx96rxSci7chXMnCVw1er5L1+h5/jHEEi020hADQtWwbRxaClnowIF9m5iaEwubKi1yZX8H
SQPABqoOjMaloZk8o/jqtUMLvi6n41OXPecWgFCApQhrd3FP+/GEAXBBjXJ/VznjR8aKgugHspuu
a+QibymJWq6GFEw+cnE1hHLtWdWHdyWAMvSPy8bX7jnzTCvNcfl/u3DtChspIaU+QBiagxCPmzOi
nVzXyQfczhxvnQE/SlEA9FdlcIpay5fAm3e++wMpNXeTh8Mz7pAWxhO+aCxfa2xYaPpbZp//+CjC
qx8/1CR3BQ9nb/LP+eX0C3AQ6i16qANyWc6htbVmJ2qVU1LidYscDEoi3PX1G6Nh3m8vAkvppLhw
EW2XeYzMmNvNJF2Nw/EnijSV4Ocw66NVMnj1q04fHAK0+EfhG78Oi47/hbtMAxNdhoaveyfigMbw
IoSKCehZgfNld5iRNlz/jtfMa4qVrBvuoLcZtbt81aQ1/fqf1vZMR7FOYXJ89cc4nFIIl5hxiIuD
cU0E6aOHEqYpw1y8Kn0uypYaZK/V86CEVzgNEweY0qIXAkNysVT26JZ9ZyFTNC8hmOQK3J8e9RGN
M0fV1OOpRwyegohmNIRuGIvwSpy8S93PlqyOVfWDsUGIBy5vZYBakp9P+48k7kDL+4HW/heHGbmZ
QhD+ebLN16oMP+wem7UsvFUjOQJgFhWz66FY6jRQIx82n/aNJKD0ShYpMI4XbdyX51BzPsKOOuIj
hr31YzQKy3XtrA8rH7UqBEUxqJWCH64Zx1xX2Ud5gbERncraYcnjyz9+PWuByhD3Ol3iSdPQuLDO
4iWJJ/oXEfDTIaXpEEbae2Fcc8VXj7OK7Znb3J8hxKdShnVL+pPLUytFNe/YF1iTQv9vJxa9wHsQ
24Q0KlKM3qE8NOjzuF1h6ajRzMMiQGaOugERXwIxVqmyg21t6455QW1O5o4qGQKZlGmo5RKB4xB5
1N8ncS2mseLLOgCR3FX2WM/BenhFdKcliWM/iXwCMl9A+J9Uf1AowSyTlmb9339VosULlfzA0G1Z
vXEGAlIuqFJCGJfIQwLXKzetPgvTzvLIr4GmNacxWJgOLf+NBwUr2c/xojZ7suMitL9TleElc4GZ
+d5Vzeq4j1rcK7DRnzGJ1OfQ3+99dGxlGS6ZYrlWH15sIQyjJ42p/EF4melbsNkV7Nm/k7jiw97L
ESXf7ghM2B1+pkmPxoDSA+wC+wbVWmzlCnUuey2Nn3ZqwKCe35x45i7Ur9o21AwV4mGJPse0Je32
tBTQaRiljRhF+OIr7YSSE7AYe7VnoEYRtTynOz6VmSQiCTDZE76mmxOGS0PKD9zvuOLtauWk5iKi
Nm1N/i1iaUJE2YkBKzW6d3cNtAJvBz9BSVOWveH2m0vSZPblJqJZiUMnPokxcBbC/Pmu/9qaLwDa
+LCBfF4eBpdVExMlkABg2IFcmdcXtnEiGkSfltCSOaokAaDt/MaNwfIP/nxTikxl19a1AuBSOZ5W
Mp+WeuJOI6V8UhcqbpObXn/2w/XZby4Lhkn7IojjsNOr4uEouJjjNpRi2m+WhK4ZU4Z1ZENEMcV4
b8+0lTPX5BMbH2Q6gpa6W1huLTBdX0/MuktVL3rb9/5TiMQOB2MmLikqeth/3zzXRSGhT6wM6Jap
usoMgvhUyx+KPiceIJuiwsl2oG7vK85ojk3SKeZELMTQDc5LG+sVch+53617g42q5Aak3PzHeitb
4+Gj3MWQPvMOl1tRwWL5Fh1swAZQTxtI3fRLxuLhJofm3qO9rXLZcc/RxDunin2vFxmA1VzwK6zr
qXv6PPGE3B+fcn67wF4sR69XuCBR7to9JUuY8cD37yh8Qv1eNjVGqk+OiALvh6PimFTZ9xvnKGb1
jgHWakpYZlFxS4JlILoE3D6MtqvMgUkDk2NjGLCnLG5UVz4K2++mKONpyfV+9E7gbQRhYmGxaag6
8JvGu0hFnipydYq6xIqA7J/px/Pgk6P9YQFYYawtyxTEYhexfXsdvKAJL1oljXCJdzhZcsS1bWEj
i9eBW2oO9wqLpNntOjyN04pAIiRHsxJMs/meme326bLTYk7vBkn1FGJRBk6FGj9e8TlefS5uvpb6
mkmHBplp8Ck+eco/wpjJCL6+iDA998NSNd873311+bDuvpNhrZnXx6ECGPGGL5fpkMgcNoCJjPAk
SXu0l7GztA2scT4T3YxQHNZyburIpfCrMyPwECVSzUmPLk4/xfID9s9TrioZInBufuFHPHifvjwu
AdduQJr3XfXNwo1tOFqp+an1Y6TblV5n9hYfNLK2pxxy9g80I6vS/Q4nxh3r9AT6TduI28ugOrHX
HYSpUyiV28qa5Vwtuc4PgPoJK5+bmjC152EmzPKpnKRJuGI3zpKt0qC58EIRB4baGwhMfhy1PJxP
dDApik7wTUJP/3+PZoWqADhlPlceAHmXS4JTUFF5B00EesI7m8oqUxpKfnuCjO8Onsv36avi8xqv
DlgvIjBAoY4zhqVlvIliT8mxyeF5pHnAsSxU+ZadI22duCuoKzM3a4KthXF8kWmFgqs5LKq+sN13
Z4aBGYecIAp0ELf84uhg+cYk1NVgGUR+xwXbI3MPRrpukhOMYaZBYYR4Mw5051sJh7EX/ymTyBZc
JjPfgwi87YVPX3X9RnTnkpGDg8OoDc8qxuklImosLLhBBF4T/Bm//NOLXpXQwu+ol+Cos+Bt2s8R
0DH79IY8zXt4bJvtH8b+p0RP3kmOHCCQiZaAJHk2737vpfSox79+la88RNnHP47iC82BrKs2jude
jyQ79JaSZZdUeahNyC1Z8AQzzLZG9vRMaBHxR4iZjbgZfkqoyXRe37RxiYrczkI6er9aaNI1nyjG
gtlQRffS1XyltnKyMPDZ1vUvT1+97K5ZOdCSgfVxEbjzQgvA9WqNto2z7c/nv9i8P3rfXnceJhb9
mawTewdLxgX4XKEOXVK7hWFJLHIOEEzyneClhu1CzshDvhxcMC4P+GeevizBkB9vXlDUTSFYfMY1
op8htQrfLQTYDL5FgvqENeivVgCFI+epKi8VDB4kk1YgdidSH0nEvWh7X9GN7G318gDD4tuFCNhE
kTykXcDkXV7BYjnz4yZ0mtVswCnth6hOiCmIx3/bbQG6/EQOFUXg6ft8ZQZI7HfIr2GxyvjWIXOQ
MjwLnU7PFuBxG1BNDYwEJVC/4fAbT4FpIVagCDXrYEjQp2JkLAVss1sCDzdG7ekaT0vP7gbVUKq7
vjbQVAiVeAYVOujxVtRgwjGuIqylTgbBeYlMxHGTN1c+BF9K2ZjJu7LHe41L0+S+A+/AyfaUR0IF
Y75188leoARH1IY9bh0OjQEAuCkAqx5feZcWoOu5lnNaNtP7Zc8N86K/IpZYf3kC+/jsx2/L6Dwp
tDaM29uNFSLpQcv8QHaPRS5E/1YEDLZzxprrs7xDTv6kClWz/V6LM/R22l5JkUQ/QMdaJHy+J51+
141ISEEI910L0PWdRpSPEeScKkfnPCSkNwVDLoERw7ivuC0kAlXGwDfdHHqAw7m1NjSTq2m9tYg6
OJfiQyMlp8uAvWRBGC98BlWFzd5Oe3lYpqSSejq5SW7e2WFXgyOmB0z8Gxg8rV+PmWVJ4NhzQzPM
xqszEhhCTpjY1ba0I2vlxFJkE71zIEsQftfAYadm4POizWptnfTU7Um4NhG1+3UWKAmf4vj4ztLA
SIsTR/n0PxTI0iI69M+siUGUYSBNg2tEMe3FEdlXXp1pwL+RMkZ/plO2AdE6y6QgT5PkAJQeYtSF
hIXuLuDTOmDJCrNkxisI203xuZPpf1yCDYBVkla8h2yQN20JJ0YHDJN5bV06fm5rdeblqj8cKyA/
I3AYWn2+N8H/EwLb2MuTnpGpVGwUJp6LHneHRuxMrEPkU5GP8uOPaBa5OcS9rOf5m3xEW3jKWtHy
u7YABqgaznxtVSD+EYwNp2q0bKkE+gJPgI+j0BYBanp3XEpAr/zeTLKjTS73HHD1DpvaUotm1JE4
EGldL3gmbYG/BLk2zH9n6bCNMlUSras55qscBmEK8cFQS+S16gqzAoQl7LG7XqYMVKxDqa+sc3f3
g1PuJ3seg5TI0yyQdOyg5fYJsDBA0DlIoiDQ6mJ3KYhn+Q0cpTZOsrr2XcBX4ssTeeQOuKV+Qyrd
lILlzI4ou3UtMLJXGdQVI/wCDqStV/1KrPboCNigau287Gboo8wNbUrwjBSTWIeQOGBXrKHqzRz2
AqO7jzlVyIEx3tAZTkLqb/HTfOGBCnwSMsRFoum+/txzKk3o+LdzpTz5FtgQYlJuBw65McF8wmYO
gVkLN/j4nJa1V3Dq6D+YQpGmVGdv+4jHg6S9KIVAdUjeiWgKwEzmYfr0yUoEG75js8+VUbyayTfK
EYQPGrfQYttFF7M4TU60t0HXQtrId4MNBRCUDxS7AXzG5PpCPkcjGlLnQaQ5Y3qTRccfZuflYRvO
R+YDMqv/SzthE0g2Xgr4ByllnFWYScm+u6W63aLUeIQGsF1Vo6hgILDcCpceh5bYFPT4q7CMviiQ
IlR8BDGxrvzD6u0I40hxRvl3CNXRjinPicTTYKtdBNZJhSCpxTQ6oGiwRYqW6kK26i1bOoAD4xh/
SWf9jgSTqKuOlCiyeJVT3oJoUXk79wlW4wTmxpRwTStQE6FXBnpqIY5mHzjnm8q7NtU+kTvuMnJx
POM8G9f0TfT/lUISVhegoopsrGsKVJi824+lxxw87snw0R6hi3wdHceAC06YMHthp7k8YNfNjVpQ
AhfQ1353NZgfCGouwzVu+mz9tcabRVWhOv2FMwdz9VsM5MlHrzdRI6o+Vo+ED5f2Ex45+XEM08pW
84m/1JTRdeiqeVVZfwN+8N0+YvX+59ZFTZ8o61vbASgXr3DRZnjgYv/w4v+wyEiPq4OuZDOGmNsU
S21xjMiJ6Jfh6bgymxDk4Nn1wNBPWRtSnP3X3Etkh3xQXbuB6xtuBCfkBct26ySLvgJpFljmeYlv
uYprGkPz4VAeIYxCAS39zNuHT+VtnS1+qlyvoMzASeBWgKx0pPohHUWIH/hJIAEMd9JfMBIjHrDo
Pux8yCFNO8BK3mikqedqSm2Yf3COTcP0GXMzWtKQrMNt1wcGtEZ/8mZs/0Q7Ze+rqZ8e4Hfr5lJ2
bcumgkN24nnBg4h4bpq9t6T1COM7236oe+90l5gsbLY6jmbo6phMuEBgokBgnALABoS0OGyirB/q
k2jz1dHGejfEnf011x69K+VZNw8kxxnUiHjBawziopaoqBrcmcGQsCgJfoR/wIi9IEV82b4xc+uk
ke55UKF9Kfv4z+vsiypuWVv1WwM60VEugoz0Q8r9wACVMepjBCPeGUbDVeweJvNlZVs3ueY4//9b
7kk8Ej7CYwN7mAkanGaSjB8RTodDJSJ5zZLeSBICy1wS3hxzOIDfNCpuc7nNTvfmULVYJJGS1JS9
ZmyhmStIqKQbFcn1yauy1K7ZF9qtHwWfySt2UJ2TzyvelVttaJQu1tefcfq7s4MOcmh7SMf6QEhA
/4zfk8h5HWLr+azOyESZVTa1a+hjqz8KeNfh7y5obMDtXPi5LEPWbFMo98Iv6Ys6juMXmgiugeaZ
gdHhneRemmAqdX0Uvk+soGmRLMFv4zgN2VpV8SFfqBFMvJVZVl1iiQTVgMuBSP+s5yMfqER+GNXz
GGr2sYRAaHaOD/u5zOW1lSlXTpkupgReEitRkDhfx1Z6lt03U8efNPIItpy+FCiJqnIzT72XBv6D
8TkrnlqEQbM61F41IbdDLSoDRbs56816kEL4g+ycot1mkltROfXXzyEgwYRRWbOaLxyRtDzZYwN9
Y/5ihQR2tfqtOvioYI60/77xzX+WOl9ZLef7kz7TO+FK7zn93wHi7e/9x9RNmyezKIJ5ZZYfQD1B
QLE4SmL9fbHFaJTcYWACufRyoin4Fd0KVt8SnaI0tqwyT/OaP8e9ISpB2HrBdsQ8a2OrGNZTJJb8
lSPXJA3fN5GpHXIDgP5i9dATPi+sZldVwsvw35qk5Iznw8Ek+CibzHiKWWRdugxSNTzi8nCxPoai
1YyjVn7KzUhhafaFbyOCDr1YyGjrJuMAwEjHlATJ1bB75edIRqwNCYrvgbOfB42jI5mCuBHmjgzr
SOHC75dJtEO133YxeZii3zxaF+6QhD7XAPKNsL/tT8UfQ9eevW+hmpGoYcXB8f5XQlnmYAgjz1+O
pM1cqlvpgXqqYoof6qmHBOI7bp2INdO1qjhJMGgRrTLPL+pScglYw9OEHsowgUQKrlN61qobS64k
hLvhBEbffBmLi2DUSVGIH+NL4eOxSKCd8BsVPRCmHTlFkA0QOJW8Mm84u2R2VlXfk+3dvMG3zIQq
0yfrYSzWAMIUZfLjVAF+B1iluMifR7SO942nU6kU/FJVXns8Dvf/wToFsvePie+/PcCgyIa/u+b/
lVwXgLhFHypMfgoeFtRsmto5x24aY/9bMqH43cNwmMA+Q025cDpI+dTNmWeDR5Gm/kGKfyGZJ6t6
mZ7L06TvD9sobuZvnjbt+xQkLShLOPpfBCdkXmc2D1p5o7cSFbgiVNxKqeqkKoR6qIVGCQ/Yq+Hm
/1hJRhDNE5xFhiG/yfvhZ7kAqky1L5RHmNPzamfwrf9FJVMUtz5dOgcDGcnPB7QreBxUMoWPgTBK
V+rUPLKR+uah5YevxhusS0DXWXMHf6j4+o8o1O4RxQDoy5xxyeMHPZ0PSodQ26zZAgGd00bnxzTx
wWacb6wFVgbePgOh+NnG7tVSGhW7/fx9oZZi4kYdS0czud+TYQRdYqGY0NfdHz6fQUDHKDCz2bfx
jm1rodCAqYt0KRcJAXZ1M+Fiw7WBsgxf0tNMOnEIDUfxcINVdZUQe2cPz6ahLXVw/FIDdDdHnrrF
Be3MvUTXnubY59zaQWZHcc54uo2AfC4tWj11fdwwlPvrha8Lu3tzP4iZ0nB6letq5qyb0rIoHpKi
CGVjSi0sTqyWtPLkiDw9ZOLGL40OYFSdK7JOruG9JJZHkrfhIR52gqzdtyVrq0jSdGa3znzJZWIh
p0bVO3B/SzkR7xSHH+R96fFW9zq2mA60pMQtDyH/yvb1rw7rHQs3CzAW+ZrSNbWHzaaWgjk89eES
R9NRFkFRpzrY4QGAvGybPuKV5YLuDHCWrGziiO8+T2MDAG6e/eS22l9hOuIamdpmvIUxfhHmSvMQ
oevnyvzxoO6FjrEI6Q8G63RDGOZVqZ6eHgN+NLdpSDIdtTpoEZz9OlPnOml+fu9qDVV2dm8mdoJl
VJFasV5sQYgRbVXJsc9FVV151OR7JjRVkPW0AHX8Mtakz446Uvjek8auJz71UKdX7HZJJT3gDpDG
gndRvlLdIqgyv5eTW+iVL6qeUx4Uau/4WpLwSMhfAH+X8OUrsYd2t89uNOezZjorY+bkSkdnV8Pj
LYGjhgj9yO9Iv/fQ0j7XJ2YvhqjqdrYe7JzzpC5tLrBVD35IQZACuq971WIwk+3TyHGEjQmV9wwL
4kRPYdgISsIChLxqjCmpOJkFUJVjiGPGISm5bCn1BCFZ5cc+W0Jrbe3xGBaxkn5x0U8TtJRmuF+T
Hyj/qR8/3uIYy5KljVhjoMqpM1lgL7j2AQD3xK5j02+l89mfqyWMk98FO8BTItEWqfJyooQLZEP2
bEV+7Nd3XtMfhnFzbOmNPG90fC4Rh6O9BGbPR2iSO5lrIG0E3z3iloq8RSNtrl/EY0dia4TKjgOh
hMEv9gDLscrhS71rs0zaMnGFeLu9FnHtcIB9bNWGWpM+iT18/KuJak7SmdHCoa4Xsw75XLyPvP9W
dHYfQuBuUQxdfgTuHdpumYKqd4Dnfs1mVeintEHXeLEuzwq61PGSrJ+qzW5GLpIF1oAFMF7pfauZ
kfX2XejF2/W5plYimSijPSV4OLIsfOVetlg/hXeUKe+z0f8X6unxJiqL7ZrtIbxvO7P2oGm651Y4
TPMK28V+fiw2ZBIKK/FYM4Uyjca2MdACXJEgJQptfuEtosUvGCgNgtD+77LiXzbzVQoPrwF/w8sP
Ajg8DphANibpGfUOC3VjGkvrcrFblB+6oPIB9Is0wBkAyFEwNCEbRym3FMOA+ihyl0tH2QAiEoim
nik+vqR9whY0C5dSqxGPy6rtIevGQTw31hdfRxgJII+zozemRuD5zq2kELwFM+qEnKYiux2ueStM
oJnoHDWA+Vds7B1y9viROO7AlYdm2oI2wFOonTT+iXprm9kJXdjlyxV9L51xEGRlOKuuY0ldPvVm
y2pkk4tTulJHxraminZZkgE4EIrtzv9B40mJ//qtPW8vAYM3jeqSRjWCMHDeE6AlSpH1ngD9RlSH
HkiGMwo83ktdUKJfo9swgJ3bvgPlZyQzw9/V6ByHtxomOOPPYJS/qqtpVDHrbDwraEguTP9BYW0c
x4IZH5zBzXTpdFHjOa61jgqZ7jUpSegBiubg56aa9uQG8xAVhauFyvyS+31PFF6PfDquPW33zpWK
wbFfJKm/MVbCmLxoAt0cqkMfRFYWWFObwrukRFKvuNfD6lnvZK4TdWF90lNe9yl06cBwTCO/B6lm
cqD6ftJQqFkI51dMJxb4AKgCfwHSiMG2nRDjlwRHjUf+onitFc4FvWSxrUCs2RMr/vqEXVrA0Sag
S35BVn+MkkHC2sHGya0ZThNqdt1InUpHFUtGATyYeYqLgyaTui3qbpu/c3s7nUXPKwH+JwkM/z2Q
7jmgx/6Lc5MSkVADmgOI3gLS8Xyp/0WKCG10BzuyF8HOWYriPHSmkmNr/b8OYxuty9695OQlLOFF
1Skvt72EA+wECakyXmUArCXAoqtjEItQZy7XajaL6n8BYy+r03ZwY30sdLRe1SuzafJ0Ju97ibLd
5iDL54rMdtGeY5/iOpCxuwmDqp3NrKz6DFvE96K2Nq6VVELGF/olrQGTZEfLpLtTVvBBDxCxfR01
4sTKENDLel1bOSTlQZvHcEwcYIzp7K5eHNcI8gmbJsSPbcIrDsFSc2AR4wM/OE6kWB5biS7M4+hP
+ZIk42pAaAp0n8iqqX6xPmNbC4QhisOYDnm1HNLa3nhVNhk//h5G2j7ooboUs2NnQ5BUjyq0A/1f
WmYX3yjy8u2RVZyd2K6Gat+6ZD094hrezWeojA6KLQYNln9tFmFTPaCGIYGVh4cEMzT65e1nAQ3F
/4QkSEA1a2NXG4Y3mmZErB9Z2XA1cWaM7Q5LWP12qtxMF4O6ITxah9Iap5gn7MeVjsv7mkf/q11M
zoiSuD6g0WmGOV13doWMDfWpilEe+VIjmbw6pF2+4TWNihgwG6k+1bw/R0hpPo4BvOjx2tOqlJJp
Lki5KXQmiRbXK0jZ2rj3Zm7hVQFtDgdbT6ngn7uiRy23rXx39QGHHr8RmCidYFCwc5GlpOlNwd3O
LeWyu4oY9cRP3NcuD6sNxME4DiEDzwuPaajUhDZGFhHPgzE+BBwKIZlR6YGGwtFArM73yiBZzH1Z
rWr17VQuhgB+FaMU3PlSX76tNhnmGb1qXL7PD3zIhLIxS0OHC1FCCvinZqPWE8s7ou2s52GZmHVM
U/lVaeOfv22yNClCDZXdmgMft9j+IUHr9IJjCCBTpioN9oAvOZbVydylOWUEXH0CDR+rrH4sGyfq
wdUly1mRPnGQWOYr6Bh8za89+mMXCVVNDT8r1RWs76e2VIK+gPkzwBZPm5C2NjUpHFxldhWHngMv
Bm2t5lddamzaRZ3dkdC46bEdTM41fyf4HSlS4Xdeim3AT5Vi2uz634+/PcHmfNtqcCyX0uItCU7J
9O7J10daF8VrEfJXaPOCxNgBeA9iCK9QHk75KAiV72F3IgLO6Il+huBdXO+W+xfggZ14wAzCLkRg
5O+4lAh2OnT7A9yH1C/AU9lchaqCqp8TJOtYtVOeaYIdokGz8Bzjtks1UEyL3ftonnwgkOcI6n5I
KCMR5g8V7nrFz7EdYM574INDV/u6Z/8kkKOElKNRzTvhKmORD+z8CILbWo2Uc8Dupni444XYthBz
OObCKqI3FF0NYmMZwPr6uQEEk15cvAHsyCmV/cNazRoxppnn8YqVSf7xHF2YcnohegkmYJFGQ5US
EaWJCCaXREZtvUz77gJkQI4blKQm/7Yu0Fnm0M/FELOam0nNc3feKLmNIkdP/JIYHz1nX3obQG/l
7oFQ+3iTbonN0XTXC+gfg8cA7378HW7LvTbbjmbQmff8bAHKMxw4xX+mxFh3ZHTQopa8FNVANTKA
UTLtyQq7VVvb9pB17epoTc60znzUJwR/pfRQ9xDG3ueKoXdLQhW3HyCJ1U3dZIcOEf4R5vZn/lI3
okqmK3YYfKD9BNSyrQXgRGIYtcqdxUHZ5I/4ygen/aG4OZDbJC02RTIaqj3O0CQ/gPMhpFMoZOOZ
UxxzzNY27YYux/fBMNb8le68Zn0KAk9n9Yoh1QLUiP73Yas5WQL0X31fUSL/Adv+2AyUs2IM0sAf
OWtRZ0CrS3ldhQfkFzrWjaiKhDjHEmRGRqwMts6WkuitIUGAtrTJzwatGlgPxJm3P46+rWAp7BSD
1NapSNGZrhCeyyTuZxzBxGwnSyh//E00fhm+alk/QQmcwJSq50VdIiHaEp/BUEaxidDDIOmJiSXx
snYWeXMnT4sRTYAtJi+N2lvNPHjvDyRfy2umiZrz4qkN2tJ61uyAB0JJffbnu6WOOovIBA5iQ3rR
vHJWKroVhd2EMMIyoLMJG0z25TVXhuso0JkGCVW4hK32lXQQAqjUbfMrKW04ng4TrZ2vaaXNHFp3
ccUZKg8I9NC6CzoXfNwENdZmu8unIsEtL96/ILbdGJYgpOdIQDn2K1EsSsPuTJjjuZ0HwbQ3wDn0
8StcM5bMIiagfai8l1a+5DsuzRSDtdV4aA1dNfmyOG/wse8wjohlCCortKrozIua8DF1pbtFgbyn
q13ypila0LmTyDBLsqXeQqPZ1uQUijuVFHnGEMhB43S1Uh/xRNvrjIpVSPXKBGS4Wbi8zpqhPERz
efrBzKxzj8sMLqfuRPv2sVLfxcVSn5oM9mfnCZIBYBAbARQ8DgHcsHbcoCDBz3QsHA1Qybs+6pRI
yOIo82DLwv3OAMqbrdWSxbrFqcVHlKxz3u8CO/KH006jtR9RrEU4bQGMkcWlJlBqp0unbXjAstLG
pqVTMSeOLyTemZwUVGFK2I5Cf7yM5NTv66z7o74Gp55ffofHZ/j8i8l1nJGrwvEpA7W79Vc76U/N
Feiesk8nxmVYly+3P3nkKf5dgEZSjW+Kx1d4rrk5eOXB1378u7igqlyCeT84pzpa23oFW2yJ7uyT
5X6+u88BMR/kWgF2PQ0Qub3SalHNf9vuRk4GXJ8Wug4qT7JMR4sKsM2o6HQFBzacY+tYpBSeu+vj
cU3lH1CXrNrK3TJzdvFCHvbOaZeC6n91dXkNRJJ41JkLWREbCh7+SmA/sldOY0rTqFxzWZZ76x9x
jVnAuTBDSXcAFrQu/JXXyenuwfHGSXAC3C/6UNpw9b6Ed6CNS0BYIzKlcOnpRFICk5vVXv+tiqA1
xVl5sVv27SkHFvs3eT96C5UN32vG2y5BNpx6nUZb2FtXYDy6SK/PkEDaBRRPZ25mOGNu7BoZUHt5
PhoT5jV6CQ8g3++bLInE5Wb/RLiErUBad+jk9GnbGB4us2AgTgSeLIfUq4HGXywR2Hj8wH2i3wPs
cVNfRfIHF5am793mmkSx/k6Yj1vtEjxZa/D6yxkc/Cj3VkOV7z18SMMR3WCxAl0VKjLe1kaykhn1
Nf4N0dpsJNv1Xlo8+sICbXPt6MREKScczf7Rs0hS4/+qv1RlEb6Gqj/mL0fyMLVHsBgzRLO+Yv0r
ivcuQ1JWvcOoy/BxGLtLqFCHZI/BaphZ97g0JR/P6sAfBp0vkwyYk8cMysIBF1TyKPX0Pq8Z7fye
lJTeynX8ugkBXH1jWCEzosqBwEkH8R8vvcX3QP1UiVvUMDodHWhGuKeiEsv9nu9pTgdHkd8+Ouu3
RvScig76CwC+bZ/2vww2i5ahfCWxWtE2btk6Ck4y9hXiEETGWjt0HZTA9BfCOsyM9/IPzdwiD4Of
KmiU669qrav0DgXCWfgB4XdBIkNuE18ZpXw12qJA+X8Zeb0huPQ8aGye/9801fkrHnjlZicL2NJ8
IecszoWhbtWblXGZo5qIO/K4PFUi8Ss6FtKwl9d5I2lcWqj7OQU1sTxFomsrYipbe4WRPNdiTVnz
dMy1hrDpgFxjRcZa4qRmolXjt3Pu6E+QrgAYLosxo/luYHdrABjziyeUL3765elP/ymBzPNU9q5v
heAiIQkGeys0L0ixw1q8ySUFP0emP+l6ZfAqUbr0TGODoGP0x2zJCz0aJgEMgLNZkMvBV605tfXt
/pjDtMrI1MNJkAvjU6forr/puiA+5i8YPTdG3KcT7XAVlx/zjEFQB8xm4Y+hpv0FJvfdwjHQryu1
6oDTmJIYq62DEn3HmGeOzdDJ0tLAIykJp3f5PPMEsQHhQejFfL4UttUdJxnITulMiTyLsvobzBCc
DxiQbxXXu5P9h6/vESJUMDoS9CHBf/GzGpp7jiOC2L/sxWmshtyMC/3dYlsRBDI9fgRkWnGTRU9j
1rOtoNJX9xMUexCKIXMntmN+jx2wob1x03Yyem9p8/32cAQ+3zDooHYHcDDkh/sVVLmmRzPIbAiN
PbwJJaiiokrmmjVwBs6IxVnTdTwKC+TfEZiyW9VfMV90SV1m93uBD6lM/SWZ5Q+C0VHUwZBzwl+Z
S4m94g4FykYMUKm6tA/CrAp4/XuPM1wIoaysyvAx/CLgQuH9BFZ9Dcmp/l7LLT0xdkayTskBaRQx
BZMUM7KPFYYhHWrzC8k4GzCmsQn8u0VDW2vpRyTC4ynY3yAvT/OaOLYMbj95FsDeUiBoDBjqq1Bn
wWP1pyUkWm1ZMEDHhj3G6YlK8UcQpHSkl5/SuNaGWOU9BJXXXZPU97VME5uuGO+nitcCpN8tdu69
aa2kuFbzwPRLDJZXd78XFsT7jbRNzLc/gR71m+9UokiwmE1pO9X/hBmvGC6OT2DuWYnQIWunY0jn
95EBiyi+/ZHlEq4cRY+32BxfPkfvTtXDm0t28fc9SN8C/QhX203vFHbPftbDrQRf33DdqV6vfiUZ
054pVPG2IEFj9iyi3XPr8RXNLH5Nc6nuqjjuXImjgeeq7BUmhUI8AFFn1sBX7QYsR+m69tJiLN42
MFH5KmUURl2hXVSnYEeynQ+k/Y7GvmyLlqrlsxU2rz6ZpOfBhSP1Pe7UY1rmUAQyQpLumj6aJ+Oy
6dDmCZvBharqp3yoPoxofHxXmth8DzO1a2jnbPfFklud47BovBu1XQnpkqV/8QY6gr0OqT4WLOgj
pttkm+jIT0rLqxpBesj1ic4R9czZpL8GvfhLgUC83IWBgtrj1UfFs3F4r04LBBpuVkCwXxxqjsFl
NjvvviO4VkXASZmLsUu92SDvtNthMDR1OfaU9vLVjzJvyND189MzadIcB17O27Yd+sp9fABjSjCl
cXYFHrkDQ/eYfpwAqJs15s+81H/znvPfOtvZeszP9ev7NsnAIpIKkPKF+uS2MZmIAewfFcQmdAms
aIAYW1N7uazdUQgnrQKWhPc+uGBNv6ZuJ38AYO33OC/6C+rA3y1B/AbxQ8qSVAAFgVIdXs7HHGye
e233cKIOrRUCJt/3yb96FyIvQdPIqpD6SX+AEImjwuy/+9D8CEZpCCcooTA8/Zko+PjJuzInQPzk
hlKUHO+qkNsPEFX6t+FC7JZv2wrJvDVuIZn8e3b/5unVYm4JphXmKsb4TT1FVFTTc4pAyW/nRDBD
nsBvLcXGg2PQhLMns+HLGGFW7fBnXgtf/QW6B2UrqdCHXa/wxioZwxzR97kqTnEpCUCmO8iMi/5v
+CLqOg8oDOrEh36ZVFx6sVgB5p19TCZ8mfbq9+S3/r6/wfS2keQASM/nXhImrvNp+394sMsbbGlN
VgtYGDuzgFEpDU1rk+jlHx6+yGXxTNESxvmrq8144W0w8Ufh7BNYrI95MHJ4HDmws2KIqrrBewGh
cZJ668FzK27qJm38QfoH+b3/vIfyt3KLJsXIdj6BDvWQ2RiyPio1NIToqi14e4RuQXMvscVVdIVf
SHpeiACoeYit5livHna3e1N+4iJIbh0QxATRb39+UdQnmM+AS7X8yGJl7pBLfqDLfXfp6Gd3MZLH
/wjIZW6DXAB/f7U7ZPSSJgW7xTnk/LLsXXdJIRV87qDpH7sQvVl/YDcvbSQo8vlQ49DoB6fYXy33
RUg/9nUgXZfSUHnX9QgDtGJrTdI1Wik3PwgrIXvoGre1sB7b5Uu4QQGswj1ZoQrOJdAyuvCorVdv
8xCrAxhD7K1taRkuNUQNRjCi68Kd79HawWKkXGTSwZXEhQGWsH/LSEP/DV9PULcWlMOInQ56xjDl
fn6vFSxK/yYBtR/mzR2OvpfsinwUwA4+ZiGkTxwIb2228DtQWs/QEce4uFafsxKazV3qJBiRwTO4
htZdaxOQCUZ1O5S2mDAJ9jrt9UNglnywPNCFy/jRf08M8d6SWDaGHpp0TS3+idPmgKMkZ6rq/AKg
npStQDFx7aBFBB0Hs/bg4uqxjwVKa5GwLE9iLSJYAakp2iQt9EK6wiCmhZW0lJROlu6U0pizSpIw
rDHnLKsF6O8aX2goI6yfplvLEAtohnFIcSgip4dp5JcoiTtG8uYxewiZCWu1aYA0RgR+0WglUsWe
OMN+/EN39dKQ/ZHutpRajE7qjnFyxdH2+vTDYf1EfoA9yY5U9qjbKxm90Fv1ZjihNXiy3XZUO8e1
BP7S7iwapBHa6fDe5sUl6xr+vXG81hAcDwwfKSVF6FpL4qapIHnicWqifvxd/edoBhNMfNmtw5q/
8Ld7HQB3wzRQKARW2FKtPYZ6rE6+jJi4MKGwTaZKr1jYosi8XKe3yr3rti5hE/RL+VhEopmgeIz5
l1ZPd1p5PhBu+/WOi9fDXv5pLE9Lh2X7YJudbPETg47L5mKb7r9w0tByjO0yEQjIV0C3zlX68/cS
KYlQxUZj/yHgY+TLMiJk1Qfo1P2W/Gurdssl7IC2MZdwVad4Syoo1j6E2p1FSatgQHbP4gXxcXsI
uxngQXgfP+ngZgxNT9WeBetaOQseuypFhGkWJr04fRfCUEOp8Fh01r2QigelA84zBH6F2Unve9J2
1zECdZzeb3uXerYpSlvWTlhfbcfwSmtE4SHW9mEbiQcTf53eZLMBOhY2/UQ0FTuYvbRFI4InZCwv
VjqG52x/KuylKFeJOgSNhDFejdnGzG1BWszOX1hv7Hvxmwl9ZWit/xGarqOWzuiZ09LvYgx4KkVw
hAheaCP/NTPLeOYklJIsIUTXeDL6gS4grzsJ7JrBI92SPFixOe24ysk/vK1eriJbIURVR7M6F2Jq
EARa8JtjyB/myCQlSZ25PWcm3AQzT6bQh+HDiq/4AxTdxUPAACnE69UnQh0Q2NUq3vxyGdK5c0JC
c+I2lVWi5LQ1h/rbbqFLKGVhnczAhh/57ElSkjYBzY6RSRZzwYRVIHxV6/NPoLBS9rdDcpWeWwHJ
zKDUnVfdwMBUsfER7GwTKmzL1GdL2VF2aCAQtTXbNpgT8cS3RtZd+jZtJDE/Us5bg4ZT8SU0G77K
uoi7NB17cEKJZK5XjeTirEVmCWT+cjGIIcQBj8GrEN912INbHrOh4zHOKRnQHsfdksoeiqxHIvDS
KR9g2TMo9z01f9a5o9AUtNKcbPl96tYoOd5mdNmNQWCgrME7bZ0BLrD6CQ8E6Cn4iw+hIpNirFp1
9pjOBtGPgbKnGyfR1glOG7f/cqAiHonHhwGAp/IKq93STZhvzxfT4MslttzBTYl6Jr+V24+uXXPU
UqzMuqUhtVI45L9hD6+Z0+CzhhRjac+na8W56wOAk+u5F6zfzqgoIscKFAol0vqEt71USkT2vSM4
1HuwgQDZNdb+kISR7ifR0OVFLjTikbaTGOi2TF8vVcYDQC5p4iee8Mikoqt3WGTehyaAJOy8MkT4
lJe97yPNfQ7QWTQpzB6zNOCrzwLwJgYUYDO2Ume/HzfWcgXOp8W0Tg3b2v4n0Ea0U4wVySw8CVlG
vDU1oG1c1ndSI1NuGo2eJh+DZ+vUFdJkCas5aM/uRzzM5CkUkEnQL2pAi3jYqgWE9kr7fHcQXPWE
+8DO+9qhOU8BXp5FiL+6+lRUapLIYsG0b+bS7kBO/DEzb4aFw+MLWW6TKBFKA0RKCpQ7D+ROTHa4
Jbe/ERBVhLgBQLOx0gZ7W0swnxPd4t0UtbHdjFDCAPDnY9ZCoCl+pIf93Kd6ObnP6g0pENn8u9Gs
yshUkARAws1yLfy/+M9W31qQu0mR3rXjz+Pg2cxCD392EwWXvPGnemDijJheiQoQzn4xd9RShoan
OBth/1rxyJNRdOghbkzbEnxOyZP18hwTHxDdZYjQxlEhOZzxIPiiFcJ5xE7xi69oSy+2Og8IHUUb
hm8uhVsn1mEJAaHv5O9ltclgDZ7bt4Ym/vOMrqzPJ/NZLVzBcmpEuqITSXbJwlMDinhn93f1ZmXL
LjycWAa4HYO8sup1vRdCFYFRtybQD+pY/KJrmIQnwCSqbTewBUvEK3EDxhol73P/YcN0/OoCXTqu
M0xxXlOwSBQRk8C6ycW6yELiyNcSpk01BaKs/TdmgUnKEJNgJiDpESejF2xoCur4hyqz8g6CoOLc
YXjwC240iEr+fAn/1f13anwJdLDgxwDSRFTkr1LFdxuk3cJ+5uJVxrpqB3lOBxF2xV/shPFHd3pZ
pyQNPBW0ORqblMhJKKb1gq7vIRRzu4kwkhuyAeetHCN2YFPp2zXZzYuO/jWQddUdVKXtX9JAN8TH
WT/FDEzpIq8nuRkbagYINLzdJ505GhYN1FNrfuAQ8yThnBF4JPZIVivrWNkrUUD7CcvoYC/TE3z2
Uvx0Jo/Xdp1Icylicp93BTOLDtZKylc+wbsboMbw+BY6Wpp0QWU2jiubNAjibHwck5njJ5WJqtUc
o/o0FGnM7MsT/x7h7eDHwCSKtWkegJ0pd9/jHmjKZe4H9lY6Mvax4nZ6tkc4ZD4XjVrSIKd8Butc
FQ3BHyUkxojHWQjhEUSlp89RU0c9/zZl3FCL6aODio6YoqGdInIqJw2tr+TqvQVwYFLqSk4KXAc8
/kEjZC4KMM+jjC5cqFFC8KLVdRvOfBYDjjGCS8dBY6wsCEX3A4JcaSW/BlBD5J8cveK2RtBhO4vo
SRPipwNQMLf2TOelC4le80iY1db7s0TcolobcHfVsoAxNxywIYKJxELzl+S35US0rgvZsTIAyPnn
Cq7v4ZcrImoo7tknb6olfBlZ88R13VQcJ72tKVIFLQhBv2zPN4+8pi+595R8atP2pkdrUvx3CYK3
tvgXu4KzWsFusG/N15q5m/omRPtR5ZnRF1iN45PsxhVUzvEqSvg/y7SU+m35VFzomNHpKtm6BUQR
I7DaTBfhD1lp5nmVhcz++2QsdFZmKa7piQx4BoiHGKVYQ6DjZdS4dSnnsw6C04nnF3+r4wbWS4Go
+mmnqtdmfKCTMWPaLDAxJDWxdTMHMs7UbabxbROH2eL7H3bnRFLCmCl+ZTL2kLlMeP/kh0YCR/u+
HT9Rlj040wtrhMwY52tDWcxWkxltYWNOcQa63/BbpeXp5CEY5MkHEbvLwSraMq4GP6LQ+Upwcfir
7qFRYjPZjHmQVEjz7vRpjQkkRNrd9CsbIexhgRyzUZsIMlY3TxkcJAl4h5kbBMbgWO3qDTHokB21
octLW0FZoNliiBRD20DZsucD4FqaplEvWDu7gabdZqV6U+L/qz9n6FebGRVs+jlCwhzZRvqg6A4T
JPfO7yYO7ZBffIYIyHUKF0gOqmhPrk11lCSsOVn3tiZp+qNkcOXp35Uq0i1OR4UsYzWMEGeGU61q
IAJnb0ITRZOI/NTfPxXU6QWIFY6eJEqW9B824ESRWmCU7NN0aX6QrPgHbh0P/U/tvgMO1s7mIpCq
tP1MntzbqCUI6mLH0oxFMQSn6lq2Nc1JRUAoOM5HC3YtPAXY7X75MRgUEQ89VW5ZV1sNmWiOADCV
HB2wC7754BSGDP1XiPmBJcKJLrBaxK3xQPJwb+qHLyLKHE8ewAIZ9+hSzHLzvFMunK6JQsO7Tv+Y
/M1YyJ6Jzh2tvuYsQ79imlAegLRKraQQOPWAM6ePshlCwx0qXukIfWglvb7sGFwl+h4lJumeIy/V
lOTr8RqF95yXIcXFHpj+BwZ0E5R9vhopg5+TM7TgD/ECiGym7ZqGopefHiIPBiYa5E6w2woNSN1V
mWtqhzfP6Mf53nPB/sv/kvMyt3CoYO2y1kbeKZ9tEpwi0G1W5i7mTiBuMYxt2golYqjYT4eKkRHF
9gLsk+b7OfEwNxsUeGwxMS1QSDJjmRSdZmsQ+2OS2n/x2+tkPMbIg71v04SrRx6wSu0Xop2nR7TF
5dAVgNQbcFveNmX6tOm6JNTQQgDl0B4jIY2u0goZS+6sae53oTnNGw1t9wginaNYkd6Ev2KqRE1o
NjD0IgO02WjJH9UT2wQOSLbMhcGCGilE+OCzMiHtyk1gIK+lw9mEOX1yyUyH5k89QAl+qUImvCeS
EsHMx/JPlJF+rY9ooE+3yQiZjXLfankPBzXGRU3MdBHf+5g61n+R35Te0V0/8nlkaetoQFtdTHaN
B5A5bVxWBooCnfEzmWBffFMhrb5t/JPwkizGUVs97RlyvqJhcIOhTS9FDRm4X4E8jF8N5opNQZH1
Nyd5BDGM3T/iVV00sb0KK9ntridn1fY3YuXFMhrxkq1iNaHvvMN78UtyE6wL5A90tgvv//QvlfEW
gN8UhgVvxxo7F96BUd/WnK24PNd5zmYKh7nF4zDKENU8/O9Wue73S1Sr4eNnhzb5AjE9fNXatvGy
pp8qzBNkabZw/SSGWOrFNMsvlLhqfCAm1aehj7vYsV1wAeuQBHKwWquoPjCw8atuMkIrf+H5Q0en
vESkB0i+PTleNg4nBwSey+ZKTNRh7lPGmghGYyLkLRg7iuBwisbgBRifieGINeguUiMZrd2Bx8KW
8NEmyeciRPxj7QQO8jybgLiuaclN51Pq94PQXYuhvBS20FDIXSzEiu/ctj/wd9KFXc5jMl1uqCTz
Nfjws5evGMjJw4EHd+rnSV5U/R474chE5Dp/WKK2Xdr9OUFuDuTJTRDu9RD4S+uylJ1THlrNS7vt
bxaS+p8Yp6NOu/pIi6XBTCZsUnd+kiZr82OVnruQuznHNMabC8JsYSAB9DMzoP41b7S9dEi4Vg5N
cPnavncV1DzsvaS93VwueY6dPMKYItjo5hwwP6XX7X1w+4RRPAoiRrqChD6Lu6FDDJLaG8Lej0dP
qRxiFQYsMoLUwgc5OnzO0jlGZwD7cHzwACQthm3pWBBRxyz2sXHCj3iAs0BNEnlo32DpGeXMfn4I
IGtmwvDEXpBEDOEU4z+so1AS0cv3fl+/W/y/yWT2/Ru9jc85aM25339nm0ZQAOAdi8QgA1BIuH7r
uF8ODWjbhm2ahJgilMJehv6IslsoQmzrtIp4acAtvb4xkkm6Gm79hEDff393sek3aQ3PB8E4emeX
kZyYwooGpL5yIKvD7qWzeSn7nQAvsCiX8o6/yUi4mJlUiRaSykVjnyPelAYz5ZYxAnMQQHfsb80M
PwVa1FdveHKFwI1bGHhWM9T0tDQf4aDZGfYyJ57cyS1rRe22Z8BryewFqbaVFwEaxOZ1bMMSR+1x
GYcaMv3nqmtziJqD/DCpoR4czgu/fwfYyVFuQwn6zYzPtsaUZvoyXNeJGik1Mh2n+1lawTQAtmR3
9dXvd8yIG3UbBNqMyTFWKJc8zsrQnGrj7+F9BahxzxvraU93/y5yH0IaAatXYKnyuTEDJAlerw8j
5CCOT+V+0AeDCoJL+BmiXaBynmCLswTP2Ht9W9Ph8j6OKykFdYlUZKPNCba27XlRleKCPI9UBH0T
EqX5xPM+pBu0fGa8HdOk7wxHisr/z0eiXF7FECbisKyLWucmZt7/teqjea8WU6/qmkYpKq4o1mPc
7oRD8fkXd3b0rkG+yAWnXnn63Ux6mKsyC/VEMGpkndEl4EueewgWuRK0J00AH3YEs6gBHQVbrWnZ
6Q4bcBhA4OyJ41OEBAxh6LGmdBEYCN68fDr9sa/1LTUxxnHY9pLhOF9p+tEGwXLASXEbw4nZN98l
02yi/VN5dleN5Mq8u5UKfdbwyZsglmjdWcC6ZTH6Wqy2rQ/TaJYkLtgG3NRfXckAHEaT8E2NIV+t
1owzOIEe6qSc1hE/qBKOmDns4gqvWYqChSjMFYWnn8hDqky86L7AUjkcFKrm3SkjYR50PiwpUK3Y
oy0URYsKP4znIajJXOe5LVb8pFDlaaLdKCIZMNFvVW1RX63r3nMLZ3FBuWMFHCnp03tUw9yauaK0
wjeY3sJOsDlEuXSVpWVhIH8hDOLIrR3PJ6zClkf9XuljHfziXQwvOIDYEr310HpdquwEYR2ZqZlm
HdoT/kIr0Txa3oquiz9MEr1ZAhWgYFkZGaG93Lu/uTtRZ5IygMWsLPhmKQ6qOQsVeaJWhMDfO8hj
jV5/52ddOhaLEbSumdI8QzBsy11bpfcpJW5PCiwgMBkdOkhNfepRGoRDwn37GFkHVeSTpAPIGo13
Q8uU5PBq/TUIi2S1oBiGa6QY+P+GJJwkqGS3iQ7M44MyAO50JdoqM4Hpqgq4Sfruh8zSYeWSbdZU
TIJmK9uCIyWS7mJAoagzMOr+kMprwcNbg+91Q85v2G63gH0wrrR524iJqhBSlzi1UzcYkKTdfJ84
wr3eVQPbcmshTj1ZnTNvryke2bH5GG86MteTQ/YszeTGJHNsiamaIeJwg+1IJPktTqowBiq/GERP
ZrCXOJRio6UNosGseMOlXvcgQ3vn3fWRPzZpSaXcmB75PSwk2elmw8QU//QEQxuABWNjn76Q7Vfr
qMgUmvrkKbMFJ8MDN6LiQX1/H8/cduk6LzFXLjy5jER61tBinHJvVzEsWhZF1BsoLuANb83att7P
gtYRf+uUoUV2V1QBYPsOXNs/86P3KGJl+01ABsJfWmInhWGyl9G/cTwvVbvUoyA95wLV0rRa/1nu
vSGkXEE6jVevjqg2BS/jigua/6Ps0ygBaStajVAINh8+NJk71917mA26GLAL/brk622QA9dx/Joz
jChlDB3Rb2DmyFM0kvhwXrZoBGWoVo+fUtGXebUxW2AeXlY/59aExsox8ZIuFb3zTejWbmzx/Nks
FLQCRpVyLv6m8+jw2cUMz9iKYnVCFQUigJDlPSp+ls229sEGTMr+2T6xzVenVpAFx7s1bdaeWnBg
F2zxaSL0WNHbcHj0vxmuD1oqdOunbHOi8sfN32O6kQaNXdrqdHGYyOXgtfaNbK54NRy+3t7AUPrK
XiUx6+PCeGOvaELiIm95Yh3WQpHQiOeMq31KGjThYOoDbgVWcCcx6s2xnFzfcW2MKWm2bUVQnvZt
gJfbV9vJOVDaolDgrjyrEKz9KNY9/xbr1JKy9uH9ljllwQQUZeIRBZGZyrXJjo61QXIPmBXdAupM
0JRoIOnnJ0jymfDo9qaC9P5Y61+Gd7OAPodNcyPhu05fv4F4QCnp/ASfTNo9+fLiHEoAre7cWEqF
+cKvzXepPZ1lj+vL1K402n9WfsrKsiE3Ykov/5CP5nDCMMlhtt6krC8tFgpGzQrmhs2RoGOsFOL5
7KwePSwagj8cA/6EV2THpR9K7AVU9O6soW3Wns4Q6mQb35z/dxuc1WaqNvDwrEB46py4SCVjiKHY
IVZmnG4qYEi0mkLiZU+i59g00MTXdKMjBJDrFD9EwQ6jwvinbf0LHRx2PvBMeBpOiT5S+ZkGY3Uv
O4gB7n1NTQBWzt2N8v3OKPYXpPe2hPd11DoIu0G5Sb+ivjIokMJD8PzA76XF08586ysQvvLQEQrb
YX6evnW9gDFe7jPHhZBv0nhgDE+zGWAa5jFj9I8AXfV6ay0UAgH5SqZpbs2+HriiGNPP13iHNAvY
jLDFCvBERxA5/ah0nVg2sF23rtt9GKwD45xsRIton4s7gE8ECSt5LNCEzAraD0bHI5SopnmUBCid
KanBIKoSJF0KuHFH2s1wJkifHmXwO3LZqm1yD3lNqwqZaDHkvIEsXh8eKe1rvpPlNs/GFjhX0i6j
3MNK3zWZR2KN17WfhIM3dUS/atObUmn8pRb8R7CDuIziC0l5W/JkE+zRkvyAQ68QVjjJYvEwR5Lx
hsyqzpnHgGKlE0U4dz+BGiv6t7IP3lfeKOqE4RLekdxSx9lqpSTK7l0HoM4CO1/nzKmuuzsuP73M
aZNgvvATKXASqXiIP7fZMe2lUue9l2VaqoUmrjO81jmmDJwk8X49q1OU8DbDmjcnZmbODpOOCIUS
DbsHPVjvcjem8KtY6kc6J+pl56ciW2aOkrl20JR5THFNVKVO7Krn594HW+dphc88alg90lR/lzF3
pZ5FjXnmRpChS9KtvE/qWuqPydCB3YA9zKBtHgvRLjpXuDrO/op1+WvmpxwDc3QUmdDO23sIvrlq
s+AE+nTNa+ODErgHssvVspAfC1JBoaqkJ+vjx8hh8xfswV3s9XWXEu6dhqpDIqOorzhEVQp1EjeF
Yr3WLQUv36KaB+JU/tFyXEfyDlfmNliEGAFvTPQoTy4Z/MKpeFEltgc9A+fqSD55zk48w5+95oSQ
2wCacR9d9XiBqfc9d1k9+J7yzyRl+NW8BUG6pmBq0mtLmds//asIqWSdvKwvtg1WfIQ6wr58ZQrP
JItz15siKaXKQ6a982hPqwlsZv723j0SJVDX4+UJEda5X77cN/8EO9Y0KL1MlQjqw4M2nSKdEJp1
fqWn/ph3puCFUXo1t5oRGmUZhXmZ0bjaED5gP8iX+bFg3fdVAaSCDBXVBQ3M0sYvQjUEbnoyKRmk
skjcHs+9qhuPFpCHoPaRD2Q3zOxgG+n0Ba1L0wa5MkBctqqcZccPCYmOJ3c1fL90F4kVU0kDfbrj
ZFmbUVLK4S+3EsNBFmsYsLWgzabfLMa2dBL8a7/SAqRwwuQhrzIvauD8v+pr2+JOmQ2Qw9Mur9f0
EvCp7lD7XzR/jXzLQvbgjFRDP+y52sZfoiLbvbjCJoGkqGNA3k+QQg7V5hG1Tq8AzcbATUjLBDd2
YciywiBvhoEcDAA7c9Xy1mTEuV38yBYNhJrT1Z4RMJqnebo/UzOBq8EQTy+zuuQkyxGV5K8h4QJ8
DUl9P6j3FOYtJjMyyn6RK/pWXp/BLz1nd/WLmlfk2uwcCVIPB+pIPKW+ZU9WFo8styAjuAAVrpT9
IiQqBfe9gPTYCq4GdmAlC7kgC45oq0Tc6nki4jHdcCSmmcVjGGxlgwK9hs0wy7JEDXMLEO8W2ssU
DzregFVq5a5XLJIEkfxd2ysiLFw0T0qrPOfOPmHLlmgsQc62qYmvs6/1nykZnjzx6ebyxmSpkOdg
mAkZ1ih1G9UoUFrUzjaKUs+Lbso0Ga1s2xcqQExuIlweE6LPe4IUAABwiNtamT/JoLCKqTJ3bXB7
iXQg4g/CLYn6sOCcn4TwsW0FlicJoWeVYI/aQaknX59DPVwkti3yHl0V4ckOZ6knPnVtZI8mwdaF
pq/PY9xA4InXMWRHNVndr3hAiWtek4CY1jAF/ZydEDSmYFmMS9/ctlrX4ZaK4k03ku/JjFacPLIn
SbNrgiTL47Bweifis1tFOmc86spsw0uNjXwx/QGGlDfPHjplioPnm4nO97wIToz7GpJK9KimJnmu
edAZJqa90UCFLfYiM7p8XRpsK3nRtdrtpm3rVg1jYqKMw9nkVdAPue0MOLyrru1AkwkXLlew2JTO
vHcki5s1n+TkkhUyLQDLvWPBHhUlQ5jpRbTCVwtxftCYnop48nNRkH2ygPDRQzH3wIx7Wjm5xg4u
5MoE558/KspyGAGqEei596hnGnVbb2bK/pwDaaeYQoOLHVz+j+XKo54yOGctQNFA1E3mHpHAzxP9
0LaIv843eP++Yj4DqAW7GJc8wV6StxROhpGFMolCPmwZ19zMlEK7WQ0ZI9AtYY8+qmscqLU5Ebok
24rrRCmJibKqDRaG9tIIx4sCmrhJyIoWxD+PGuo/g1NX6716uP7ZO7c+v2/zgszCQPA130ZYtP4e
LfKe9pAG2maIg3snjKu/9dQg5kdvTBwvWqZbiyNcuhPX2/8L5I3hARt4oz9DMHojLasrAfN8V+u7
Hfpj1GM+ZyGpVvlMqiaIief1dAGCw8bWTdCvbLxONkGW6K6WbwyudIEUjVaSIrz25tkX91+S36q1
boUu+0LFYxPEKpGldFxzlDKuO62/5pmk0Pa7COAeaosVmmv7XPehEAEH0woBEpHFG2EdUOKnnZIQ
8dyoZDSMuWdQuWMuCkv9PAVy7+tMCMZpxxnuOikCXh0KsVdQfi3o/BeyN3/CQk042qYhjP0WO8A3
Anq5Fkrec+aBdkFYEOWlvLSSt3khWgZjelOiZKUo04iy/5rt8FUlL3lRT9ZsNXDcld9a50dWMqwd
Z0Q4kyvH1vfoP+l8nHI4N2TS4Tknghksfoadvv/JAbLOZ8pcy28JjNqGBcgBw6mgJqDq00GAtZAa
6+fAzmBaqalIR+uG095zGEhYfF06fALXcp7k9PIKGO8UmlqZ3Wg2y+r+a56gAqqezoTB73tDfPHC
gwldjYRUV2Ut7RPMg8e/w48EzNwQcDKOMV+FTeYT7Y8WvPyM9G4tXIkc2DxLCx5uCFVa7fRWmsG1
H+UKceLwH54Pt35SEqL6N4LqsZmawDTT922u+oNiFAOCmQZJM3tDH9oCbwoul60fGGULycOt0bVy
q3elFLwd0APhpMw5bp/sf1CSU7H+08DMyKkbL7y/+fcC69cFvB195lM84ioHbihLC4sLkYBcVf3G
DY7uhZJXUNCBY6ITHv4lFeICSg9BExAJGk2BHrf0fOzmBKkAXbR3VsOmtnbu2TpoJPSwHwMgM2w7
8UUPJCwEGCH7oY34Wi8f21n4kAF5oOewjuYORaQorF2wTaGQyvJr+O0NSvlj1eJAXG81LjBobqqz
M8wKr8/8D5nkftFEw9Vdrcyc2WvjlmzjAzK5xK9ei8Tmx7br3whBoDB6mGYIz/g0uHMyfnRbpwCY
Z1uuiZPykVgTtLABEShbR+qOAHFMzMdU/cnS2hKa7TGIQM42Ye/jzNd6mo+nfQGgBAMBpWM96ARg
9ByFBMVSppiaDB1KtNXe7do7frpt9XODclrI5U2TbjQXYD4pTcFHLT3KzUOQT31Jyexp0XamP2AN
UVtjSoy/xeCgBG93ukNROBgxTNDrbYLu77pRgyPfqXVh0bZ7kYAsEwUtkLLxPW29ojr4lElU5GNz
0KmnbZee7Sqv/SNt1AHSIFRq0D5hlKrI9CVIGG4DVm1h1rxz0Gzm6gpz75XisKdaa6nz/aTJxi4L
DKCwGmmloU4yIz3pKy516B87WGhFOQ8QbDmCk7dCaUnqoqiLubgXRX50/dLiVWMq/OYja2/nVTIm
sVl8N+BEzfE+Dc1l04YiKhX3sfrnXxJ8QVLxHKbx6ueV/uRvOkI3C4pueOILSeDn4I7udoWaZ7jX
m7r0bwG0Ezdf5N75HWUSF/yS1EHh/kEm1xG13P1S4szmjYW/oKAMr8NS7XTd8VCriPigZDk7VsLH
9n9oVX88hiSMUkZ48oYudz4hJzGuO7N27Q55/WnowOwA2NgM2plOK7bqrm5IXk+H3JfIp24W0mbh
uBFyNn0U5xLARbjBIoKD2d9CKi73KqcqRHgN005Pr6ALSIhn/G/36pKjQngtDHkDHuqf1F2fgOZ6
RkoANra5u9gPr8psrqV2qnoTkeUnZqXYsFYpcQ2p3G/G0uDA1EJZvOyg1HZvqAnJq6gaZJ4OVZyD
R9XX5fGUVAFW0Hd6Wa4Ve6XfmWVJg2xH/yN8SjuuyTvJpoYH2u4kZJRgdPqjIvj1zn+/8Nd1dzbk
8/rv5l+kg2FAiYE3ZIoYZDlcNabh0ywwLwCh18o4mwg9yflKRUCz13ywaO9CPJ9Z91X2FgdMFIJd
hjlVD+NCdrskbWHL1OjQ4/RmISqGUyzXYPgjqPZiYVrJlZnBM8+DXbeE3AtLejlH/dVMdlXOROOc
UcbeADAez4n511WbldZSw6df64JOlxvIHQZ0POWOsX2b2Ae1p+8oN7gsMZlCnbSJKO2XhDpI/JlC
m4gJQiCpxDbj6K0lbNmQK3D+oxPr9zPF7F3S1OnZn2PapkO9yg9pNtIb6rhm7Ic568Zfj1fw2Dbl
DcsmLqP/5O4yhnI43Zam7da2063Yx7oASWInWq24quxJ3K9QJPBy9poLz+S9DcTCPIBAXTmJJfV1
2DWNqSM3/lh/tIYUjbYbbZDlPNI9OlxgVOWn9HlQwsh0aK7+vooEGhOWobaqJnINmBcBEDle7kE8
BrGALExfgBjZuis2p51RulaGplxrOC5BGAzPwsyRZFEuWfXEdGZfirIySfhucroAKNCjb2bC19eS
mCfo6BCJ8wyPYcok8cYUqEebrhK0YFQ98Bs0Us14DjQJ+6fizd2P6TvdYMCHfrVvbxxvieHky1yY
//9gl4VbOZ+8F9W+LTKc9F3IfraqP8uURpLroUY8tjQpcsULW98q7w0plzD4Bxv1oOn9PMI+6tkp
iU096y10dVWi1bI71iALk0qtbanMM6Uf0dgSvcxBV6mLiZfc7XhEZGdYU7BhN9/ZDzlbCKMPRrab
VoiJWhE/ZAHyewzTjVk0La8x2W2BkVCqzRwz0yYhsXdrr3INGbmujJNhyil1SdQBfNRMziIE3QUh
/u3GpAf5lLEGIQTVzaHV7nlEBwka4m/AwxuZUbxMLULdWTneIkPsRul+vt1TrKIaCrtDdZiNHr9X
nKNPZwxAuVLTEL6Cc8EB53lXaumGQ9n+FHK9pHtaKBAKpMq96SjAhzPr1eSgvLIhkOXL2n/DzZfM
S9cNMd5Uj3N9mHUXabifyrb1a5Y5br13wnteA52vLd/hBcytitFnsTtoj/zp18mDP1y7QVAun5Ba
6oEaWD9tsPByQlFkSAUSkjQEaf7EwzPW852Aw3ufYRxEk1kexsUxdXkqL3k4I4IqAQvGeP2WbS9O
Ey4O0tKmiAKq3pPvnKVJCdwfN6Y1WY4uJvc7Uj09MIcM3oxKY9aNHoLmb41KMToyqtCV9Cic7L4a
p0v2fQ+UnDShDkVAhDdYoOntbN7mCuN5EhDj8NgyvMIHVq3QFHqDS0SfNPVxzflpkMvjh8ePBfvT
zrtvsKjwBoGByX2j+NohqRscKsD15dj5OADh1gGAaaVJifM0F8rBYuTwatnchXzsZcgMji71yDBs
7oUlJojyHjdsV2xTf9WcmiRvD7R2auTnHm0LwJmaFm++8SdHXNZf5lUSKOzT3oT1jDe1oxBravDn
gwObpLVwhVJazkTdaFCgLCW93Gq5DiMYGEu9zSc+VoSP/BCEaLZ528DhDH9MC7jlh1dFplQt9OCn
8+R1RuLUDO5dSv63SevrxcZyNi25TLHIrSxRPL+QxtbdWFQwhQ62dZmgm9xNMCwxolhntNA0BreG
EOqFQXrp2fodNuvyMtDOnGQ9isvCX+NN0V6b6FmqVCGp+Q3A+M81Ufeg7+q5lvGH0qSe3rEpFzfn
2s+s4KXSV2Fv8nSuPwvITVJ0kGM/nbRNl2nEW6aySzWd67dLTzIlXLLmFOm7LCxfUn+9gY4KSp6L
IN5kauUcbTNVeCMSFHPozJpvl4bfpatK3RFurtWkYb/F9QW92l/wWrfEHCuWjLwxPX23xOklW6NP
Kf8IiG46Vg7Pq0QromquYBDYzrXPuGDthlu7fV7QnPyj+jGXW75OfgV3LESlmRvQvP0sVAxTAhPR
yH4wntvJeezfmpGuzsGzL/39o0TZ9dCaUbDnnixtxRSLUw0jdvJo0JxCqA8cyDr87OOOapzsw2r3
tmLvC/vZUnvoGS1QoZ1+aIr65EMHryi5XU49nU2A4Kxebew55h9PtCDTP5IRbc2B/bGsNT0UTBUk
/KaB8IfDXaBGntwTDDnMNKR+IcFRY0wcHtT5og+y5PQYOJAjYLTw2qfy2uTn6jglzvYDDNhYsjz8
RdTTDT+VUozRhcWuk2Z/mtFHDA1Cw1H93NBYa6BvK4uJHV4NhxFhRZAIP91afOIcWGtCbG4c/1N3
LjbZ8n3+bC6VL5suaTQupyvip3WTpCc4f5xF/c22l+ewG2h6Kvb4OxlWEpquxxFkFkXMfvayGy1M
fu1X6Kzcyimbj56J4UpfaVFsP4h0y1F5Yufiq/IuZfHh5K1nMs5F1sF93zo2QkgEipWEYApEGSfn
fbLv37bLOgdkORJXdEU1YX0IMwOLlBwYSYBMKUQyGgx0y122D8Rrtn1E9uDE+bCc0d+k8Ux8XZt9
m8u9XnQeiXFS/oFSxB2B2CR9pYXQ+Wi65CPk8Lsm5X3VKAXEfU65H1LLAUkcSgfGrLy8Jy6kZlUK
stYrlH1OlcmnShrEuAg6leQzDCsrs4VgpeqIFB72hbpni3hbCn4PrYOsNF/Ve2gYjwRbpJbD4qZ1
nQVny9nu7eULrjfmDxB3iQisj+ifCNJXeWlOxS+bTyNoUIemo2lHVtbuC6FXrDBgxkLQwqoEoO10
j2hU1g5YdV104qatX3WHGnyVXFP6NFMsb6f7ZvDYvmytLpISEPwtZMAQteia1Ygutha/h4r3aKKq
IP5v4SkeuBJSH5DWkpX0DIjandM1sySAzfpuYVCN7dTYSYzTsjfx33Nwpoy844tXuYvqW64addih
zuRlzNuOyxdsFFpPAcSrJMNfPijooZ3KIE3SbDhKvm0BE6RZD3Oj08i/HyEAqBEd21WT6yJoKtmN
xT5oskCwnG8pGWPqYGLVpREqTEVM4Kq1+fYRUI2vcnfoqgCy7n10/1vLevQGhvKFklIMF/hC0Rkp
NuTL9m+IAVcgZWuMWqggAUksJdEYetdtM0rW+xuOmimj1jP9SeU9bHmjdbIIfWTEZHa+KFczJVv4
YPjGnJFQgCobtXIn+rJPY6CG4/vrA4fKc4qNrNfHLwcs8ydWc4bICEc/3ffR1wMrsK4E615rBRoc
gu0JPceGE1iHJfQrDAr3RAcarMRin/yxU4d1ZyuyPWKqgiCM8wuIiOL5dGppm1g1lWF6AKZYmo0O
UvqzcGTisXqJ2SoQqzhgvooAaTmUb81pK8GYKg+pElIRDwoKa4XLExPMLyuuSvPyqk7w3cePtnfe
OiDtZSY1FqUwSkFSd5ZgeC3a5AtNuydtjxlGPOX1qEKnsjNW/qNnpd3hRrms0tU4GUeTdHlfdiRK
9xwovW26E1dVA2XjHwNnyl8wWpicNj/jkVU4eGokZp9XZIGCr/FvXM2yZi3IoQMb2DNLIB4/Ouj/
b+WRH6dZ5zTCfsDmEJAjWJVtfUpr+cogNI0Ofb9EPS9aLHQVTcyIi4b0/Ix+mXOl1FRZYF7Wx7HK
19uZgZN0fLPlDGWLTPwEjFFC20TcMioBfVePMzF5foHG+QP+vYN8zznkzDn3zCoiK0LIB4OVtaAz
GkDPwmNz1iwPd5vpt2iCeOSzkE04pKPdH9MXflkAZhX8JvnYw23CfiL2IoEouvs+zzfIeU9HhMHm
WG2vqCvDrj5+vw8j51dYH7N4RQ3OavSiNnYhAOwkVtdaGlEETAsgI7T6CO54tOmHMfD6KYLf55gH
E/HcKIE0M9i1XtcAntDXECZapW8P8YkxaGG+3TzBbMSLs6MPpn7ZZ659MVaSyCBCXTKCGDOiwSXh
SXgoklkq3eJcK1rU2UurAz9BvJMjJymjwary7pKw8S8Of4/RBbkyAQ97k6o1h+qbnfQ4n+wzyv55
xCVQY0w1TCxorRh5BamecdM/GqweI7TE3YyLAKA+ZzNzgFnggoAKoDe//EO2XjYUcpwaKECUVE8I
Nwfgy8Ucsc37rCP9TY6o52bW69U6GTljacm2zi54Bv9gGTqhJVRos73Igkblx3swkZU5MKRWxtun
4ayPo5yrGryQOEKNxHfAUqRbAv11UnXFb0glEVg+eJXjZ+QMcEU/yJc6eNfVrtEHKzjUPfI2e9MF
5KoPm3AcwfCAtyepKYeUAwDkO4KxpM9TlqZja0TUpSGy/1PsTHSDUF1SGsh6a10Yc1QrSLP3rsXf
W0507aIPJs+X/1pQHjZNUUITUOfUcI5XWkN+vkHKBhuvMFJB0c8moUVMiAFl1og7MRKnwDw90mPe
EAqwFi4lEEUk0NiE0Q/1Lxoiz6DXMxHzgJNbVcrqCZ4tsp34CYhsShLEH+Qr34goveOkI0ky8AIE
Ffozup23SBGcktbXtmoT6cSPlHfPKsd4Xh5oKItXdf5spKetTushlpD69JvPWxNoXpweGGGVgSTo
zIdNNMzURgBIKixmiyHBywo8bGX4JhYy5WhilV0KvIj8tJ+L+nG2baCnHHboM/whHo6hXNv11JNH
n7oBwEd7/zAsGwtcNhLZe+sgRA4VgAww2s0EyN74NAnpsO85UpySnw8K21BtiVZcp4llS1ShNxUa
AxZD3Z2khbu9cgegWhddsOHHAW7c8HTikCRjghe/C1HZQ5w3daxHOq1a93KwG5F9WssY4MXHi9KP
MwL8f/gDO/t/BWwVdbnnEVEVBNQipkUqy4FFnipU1b0qPU2MbJt2Xy9q0CtUNmEqtGFPXlGjkClD
XKeEmhcd1IMvdQi/Br8IonXzYaf1mLfSfwGrfcGK4yPuYwWRvK3e21czkHlecgcRfd22fM7+lCBM
ZAVot5CG84xE6goYzHvIA6QahaEeRANVZWmsxtvMmbCjoYlr1Ncz/FHIdcLKxQqPZYLvKoybxyQg
4SF1di/2wTK415wFI/7/37/DGz+EA02AK8w08N9SbM8P+XiUSeyGxbuD1Nu0lEl6lPm7K8PLzgfi
Bzib8PI2WEO8PxsHa++4Gkqjy0tGWfi2i3p4yvoX7Qr0uLYKNWWbQoS+UfOaek6+e5kYOph7/7+Q
5wSrtW3kBf8z0b8Mls5FvryTYegyuQPeR+RW3GZRSHa2ympS54lIVmU4Wvt6X4aRHrcJOxeGLnOd
NpjUhFZM1iMjYXLZd9oJEeloHU7SYA5vDjN2Sckuhy4+N+2FSFD2n6DbH3etZQzvue2B6w2A3kSg
EWNVeEqpe7msijg1PjzFO4/DggP2Wzu39eydAgZ+GA22mStDBIak6pZbBvOB0UOJr1JMjJUV9x5y
LmdYb5I7Ok675QFb8ZYYr5Q+CYdkrW1no3N0kCFTjJ+tyuLwt3yH2++2byV75W9v4vZqdKOsl2Hs
isPrTm8EkpP0YOMeJupBkSJjtaY/6tuttoKDJwgJ5BFTV68WHyqE4b40nUD5twQN1OYlWfJis7g/
HDz+iaX9HpA35Ls40aQgGJivxHUouR/Lwb17JYjT5d+31uyJ/BSepYv+H0sm9jxySDXeqv/92cJf
iaVMyrUk8m4P2nUip4MVNXefmkbfF2jaypFMDpe/tLCfn5OQ7FOIlfnEqQKGHOy/PyLWRZwTzYYS
VJoJW5XXaNA3k/kqmgNdHWmvWj8hQmm9BNqbp9cIvla9oUwtyB1ztj4WQLeV19cb38XX4vi4lSwt
eR2BFhf1hwF6ktEZZC/pqZrsyJlyvpE073v9kAWDUwQg107ThBXOYxnljMwCTpoew16I8E6V/DA9
0y479Ray1sldTzpe+MuCx8iTyQsrZAAwcBCdg+U9JN8ghBykks9yAxN4hC1xQvVBG/cztedyYv7k
iev3fpdGrszLJysHdMXqfRHajX39p2CEFdRm81DNHrNSZe7RA9FsLee5QGDdRnxzjpJWbzAYuP3i
Wf114mVDQXw39fcfdm36zmieIgvonO5g+2ehAsdfJygRu35g+b5H8sTtf3kihE4IU22CgW6s50CV
gELSNAAPX49I2rWxaGCnsBBPdrZDNDRcyp/y/OuUsAVBzkPwI71taeQh7y7rg3t+bhjYUkycG8WH
aSzmuwCOi1Nw2KSuA28U3Ef3V16Zv8qDBwBx89bMUzjbZ4YCyVH/KjziVlzUU8Pbdddlx2wNmJ57
PfQEtSD+b0HMwYLquknadDRONC17PSXbSczEsluUSOrQIV7xKienYW7Nbugm9uuPP3vcR0hL4mDC
47oTZNWI3Ox2MezmpZSRP6x0NNN3fcHWT/V4tsCwBsoHbu1XuQvLunZnP/oucQPwgFPwzxNpDjtR
I2gFhJTdwBd7EmU4wvd6GCQlMs6foOkvH/+Q+4Yv7XSm3kVgP+8o8tSDHQGaz+6W4jOXBgkpzEjI
0qOuzFJakJwmeNzIvYBWVh1fF6bFPbvd8DzBhQhNgsoyrPiyO2WhTEDqkMBv/MPA5Xyav+6sOjvG
RcsYV0BkhdgkNgF8xXTDU94GagIcO20CzKR9SiGrXuvaPsBysUmhwe8aTb6rQ0frScEiHBTaim1A
x22Spug1xqpLJQPd3nPBIsqCjDyh89Xeu87VC0vvwtDw+LOfL30JzTYBZqq7tHlJ5NoTu42ct6yk
tLHbUz5UMXG6WX3NWOC/MAf87i8z+NJqQi/fFYFhtwsy7SnL+mo7OF5C/h3IN84Pa7Mcy5NlzvXH
oJl8+x62FBu5aa+Fl75sQ60DuxO5BimWTeT0MSy4oZAt/jmTITglMMgzbajb2AqJORG457XPNn3c
D9KWqlWg7bokl4Dmaa6NjXgyhv0VRfhW+4t+C4JiUmOqQLUYeMmC60WqoW+aoX42ulbuBI4A2nVP
mpL+HsNX+vyc5PXTXYvWDaDmGNiX2q5QRncqJ4e3FicRxC5TyXp7Dj4Yk6VVzbaMo9Pxsc55kkAu
SmVa/SVA1rhmGYH4i54tpPde7zMUxWQoRF7kyhhhlY3+RefbyM3MXcJTFVVGjxPayAyuVsEkebq1
Mv3Ts8G1aHASVbkXg18MO48GF7fo2jxzfll0U/cxeybCR/SIDfTLfshN2gXuQG8ndDuncAvhZekJ
gkpGVdwa+CwdNmHLfBEwhhAa4sbxo20p8tSi9kOugnhvaQRckAW32JpHm1Kgw35k4ZFw6eSU6O+I
tAGAo9aN8a9PIlOPfcg3vPr8DQ6OmUjuFA0PPxB/iOC2Sin09tNBh3Rzr9R/TAwrK7RmIxFOtz1J
hGObAvLSn8YO1I2vl/wKVFDvWoNNDTQ0eOJjQcOBJYItCta0nApLuvfLz3aOH5yEK0A/JOG2BLOG
MV/rzGI17VANG53qmdZ5aZABngN3jKkuIhcO1x10CtHU/kyaqnmWWl3y5ZJvx5CsmhVZ2+uoNUYd
FCVgJ38d9sr8EPf5FAseqP4rCVBQPApeEiwmySnNsZgLf1qQNpFrEr48o/4fz40Zs7w+G//SESIM
JlvZ8b/8fYi6vCzeMzA+0JumhdZrLgglL/DlcDTyIRnafB9rPLSgApq8rQv8Vz/OhArHkymM1uCf
CBX5uAzT/794B4rCth3Zvfu6JBzYFSr/h0lKcmAYPnTspxCHYF3BKCIBQR91AdDH964nHXPr3dLp
GveL0LzHBOJ6+yYrq5KT3dN5QzyuuMR/GwAa0f12Lbumvzx66cxEP1o087ksj+ukkVnyttLAmW2r
o0r3oqOoVbO33DgBr80j3pFz1Kmo8Y+LNuCpAQPhA9nL3Lt71efcRUvIWWW267nXrcoxkFMWwDR+
H5jcaDNW6PZ9WwoGLNNg24xzVxFGhR/GmcwkiUD6SP9sdCSF6Y8yqNtTaxHPOt0LQ8YI/iAdH0e2
WHUIvZRkbl9YQp+5Y6jv34AA/M6GXhygcG3ZN7YoELmHg85Wg3xlywa+5DrCE9gFp0pXa3nCR2F7
F9UNnaxDhB9i+Tn2djZw/ZmsDc+fVg/rOT1TeezHw0gri/N4ytzmXbpDEYH1py9fTZ8Jw9VoT8yH
9WMXAjQk5EYor1U9QKPcFkWwU5yscktKOO9vbWssRwjstUFyerXyYh8G4Hqb/DWhjK1weAe+6T02
vD3mkLw/5EJOeNs3fAGGHHWifu2ZHJ5+zkkVKMhABlQ+E7aIZFaSCd0EaMj0ZKtckGgpLHVlSEJH
mebIc0D6YWE5Y+g4BAayqfdk54kTfNtq/tZQOV3YNNwdV6lZqlz0xfYmmXQ1Tw+CLo9ENJ2tzrgB
CnXKu6DUcL/ErIgBCn3T7bwzPH2522UF3LsEqT88+NYQNjgSkkl0fTQoDR3nOHXK4A8aRkIZsRY9
ohAXnctNkUkk2lHVvD1Y8yjo+bK2deAbRAPX1X1BBH7WYt2mFge7+rUDfOUNgQ3ERuUekux2iH8Z
d5FpipiEw4NYYPz7/QBsiA/3ZKFmQqdERi5qDrrazkCYHfr7oSyiblTDMFLoDBLKHGpHIKqT0NMx
KSHPVvd5MUlBwgxyYcLcDFIREcNYFcwe4O/YXZWCEMi+iF9Ip4Blf0bvkxX3XNeXxpPbPSESD2AA
FvT3Vy6dc/qUsaT2AA8z/uyvVzPWKPP099Azbf/BP3Zj0mhVEJnHDsKBciNJ7jUZ80Oac4kMYvrz
ANw5/cWR26EN9XujyBNPC44r6bW+4tdxKjRX2I9xVsp5jTmUdo5KAF87y2AGWtxOtHRLzmmlILWz
iPeoNolaMTq60CicU9jN5VUbTDIQQ7fSJglskBEKwqiGZ34DRDq+zc1tI1mfsymVnwIKChNs1Xzk
N1tADgCeejvORmvCbhGv4kVdLxuKLc8LrUYvAx/SinRQFeC91TRqe7PwYhhY7xJgpICpjzbcInmf
DGhUvXilAdaYYgkR5P9L6BHteDUhsaz9YLYY0AEgzTUbbMTqVtaogNbNwURoC86RhD6CmY2sAXu5
AX1xsOX9sYp2aTJNMXYbumdS0ffe7zaPHAT0fm6komvjDuOIShs0cJ1mVb683bkf8TVAt0HNg5OK
/Uo+3Q5f764bkhz56Xxq8vxeRzaDW/QgmkSK04ybagQA8r3WqP2tXo0qbf1nfaUOa4i21gnHludY
ciyl0x1/8qi5s7WXEx5JyrfGiHV+MIboIfNc0DO1LI3XGyBAL+4oSLh3W6h8NmbSREgeOHiHHVaE
qCk54BiJGzs6aY0oqL2mE4+Ku2KrcBxRCMnv6s1MDvGE9FjuDYELar48sZdx5ft5fCaRo1cOUPiK
sqtdhOD88O//838ZJfIdoSY3YFdWh6Bg19S2dIHMmhB1ibnZzhz7JhKO1hZJSxJlNSwYAw0QKAj7
ksEDRdESr0QAUorHqz6yMxH9HZTcNV/HcD//R/iizCa0YjOIJncseAlk93KamAaIeVD50yeCoLyC
R1aqo+FkiWm5o+hIUfm+Jh6vhmaUDGiWc2G6eMvE43CGKdEKM/BTLeEap+7do8yCiaQpvqjpk46N
GZfsBYnCI5j3g/vD4LDvq8XEJpclxIdyy9ICIw5LyErax0V5fmAEGM7wtXjBdDRqGcgqpHgwciNG
hyZZmCkX7U7K3qnY21r5c1/FWFmK4C6yePAPAzdoS3VfmwWPwKUh4VJmwO5VihcN9VaMgo3kn+i4
bvKobbsrDLuvQGWaEmYFDqM08IjrqoZi/bzXah6tF0BFAlrHFxCkWf+grfUjUA5PnGAPIozpMF7i
aAw/jvQI2tw4Ku1/As6vl2Sxsr4cy+5J+31iSdeZUNXfECdoQZaYBB9YeKouOlm8leANclLYtVIa
GiMbP1IR7bA+XGAo5/YV6WKlmBN0DjVrLfg1W7B34ox3FeV7EbK60yurU3nOJ5T4LZViKeosWLbp
mpm0fhAnq3M4skuhViPdu/tRE7Q6kjADmqWQGt+5cHC5PcKmlXCFXYgk/IfimKuRfJhb9HTIOvUZ
oA+z5acdcZMBb0gwVrkl5e3g8MGc46Rl/XBhk+lSOnzmTfZOtGu0ZAASUcsz1vFLVlUwf04b5Yuw
XVFoXfo7XL2yO320Agf54P6aMII98oe4hzqUvkJuZgfRB0x5+ipugkZQz4G42v/YnSOA9B7IOYD3
GQbGGt2+KlHDsLGNSQqHiF5LYu3tMnWb5LcINuw4t8iaRbgl8efkKIPMmyh4ZHhpCR4xC5HHrZB5
3vQGqD7Mj4SiTC5Tkubsq0X7iiqxqoVXCezXk0Q+zsDCbW6CmLwV0PDyaClBpHkh8eTl/ta/06qI
zhwoF5ozzKHVVPDowS0KUuiuxbfs/xI0egz9vC5MfBp3YmTCUFUV80ozQervMc28Sq3Op7a8groe
zKjIizMKru5B18WSXoLi6Wj+AMO+Y64tWtfENHx7jut8LzfXHjOCcFPdDUapE5Ol28N1vpmgScVz
qoxFK0nO4GfBFoGKLgz18O4OUKY/A6TxylPXutw141RJ+T36wyA69cPokC0Dtegy6o6DDIH4lwvw
Jb/1j3NXVzIEWQ81tWdR3/FerwX5IjjvyjkTNS2C/N1cTvWZ7tI/g/ENXYTSIMdxYHTGCrL7dWYs
P8nOjaagJrLniE6Hfdus6037f4bN+5gJzahAvRIklF9/bJxv/mmiNVNz/Xt1fn1xgmGxJ5Sh8Xt1
4WSXGpVpxISJVoCJD5pHvt5e869LyvRHzPOY2waRcphFqtjL8i2pgkNrKjD02kN1fPnfGvY8eIXi
lo3mJ7iU7wIi4LC57AzeCQjwGNLea0mMN4TMN6kG9U2/N3+l4fAcyYvpXR/IHJB6s53iPRTHB6/l
zcpRxNWJEgKU3gVAGR+HLqqQ27eXi5TI88BgE69RldMuHIyFRwhiMctAGH97kyXTP2jbDg/iPtxw
mNODvf6MSrN3cK1UB5NMRqNXls3Zaro91LFVANrSbZW478MMq4qMYLllmGniGZ24drJ8HUopGXXx
3ksVZ/tlkNm7/UVFDCAeQfK1PXwsV5IX45lfTqzSs2NDb5E4yZdjFSBIZUTUmzfO+UKXhdIXJ9pJ
W2e2QAXR4qVtApENjZrdMHIGJ/WyM10m4exPPcKULeBuQvS2S6ruoolgfYMKARV7NaDAycucsWLI
nKeUIdM9QDHIZc9A/RyeHhAMFKNpXpMdETAWetwOA2aIfRpDZZDhqYfl4roRgyjGHCsc3fRM99WX
f5jt9mBnNYM5t1fopSqF22T+Y6jmwldbGGKz37bL6uSeo6PkfMHkqcWMv9ZM9NbtMPhOswWllU/D
wNSMqQm1mR4k6nvJCWkq2NgyBJys80oZqzQJFM2k8MnHvD7YHNPe+UIVjr7GwI34G/T/1WK/vggI
4pKFCBDcPv/NaTUuvpRjSLbMfId84oKsU57Al0dFmm/wTWSGeaQfkc30xUUTCncgL+x8EjqW/W2j
csIMkeUDrtkuD7WNUm7lBsuhIU8Eae4I/L2ycF5TTFEMX8v8ke2WEsB4ZZMJPrfoiewz2AAAWrFL
Ke6TY/15kGmxDwhisi+vC/vytkqRrQC5OthD3t7bYgbo1U20C2XW3sbiFUjOWgFYWkWdjYFrONhh
80zeIxt4Vd8FlwS6b8zmmnT4Kvb4cXCrg2oaET+Xikr/t7jOvcS1FNur/Tndw+0BsFuKt0Y/9Q9s
aSM84O8GuqPkFmBck06UO9mX3oU+Vlt4RIFkZxRSHIH/tWkBLPcpg6CIxGKyg0LIQeeCs/Ju00aI
YwXI2gAFnpgzpVJJdqZD3a3xqxBST77+2XeI2u6pBgRAHBswPjzRpQTzWLDdymgcD+kO33HGDcNc
fzkk17cY0E+EhibptUdXMaIyt9rmtLhGTI6qk4zDcoqHQ8QBX9S18139IdPgRR7ISubVG3AiTi6S
MLbXTixfWdni5Ub776cFSOx4Uy6WtBmjis9puvVm0JUAPehSOkFVQ0w7iMm/SYGNpRs38apptA7y
vPi8NeNjkRPg7rcdIWUnvq4uVLvwcUcHfuRe+Sj4iczj/Y6T7EV90G6MI0dB7bxmvqPxZL9HO2CM
FVMrjulApj6Rup2G8+GcPFEmGfBCidimbMjJ3gsxglEzcKZhX5jEOJxqlPKhkNbO/EtPpcp8pFkS
Qf3PEBBBOfL5zFX5bkuRIEOrp1KwFnoUG+sKH2vJZuxLKes5vbuVIDb86bP9Nm0m9K878iRgdCSZ
yWX1wpvx4KYPjbNItx7qgYhqLKiFHp+g7Knw9NrBh/dVEurSHi2gOmZj5D8j1MpN9vwReQl8W4XK
70J0aBdftnJ3D+G5DoGblDIxbGl2oYxIpp5ze6q0aCa0hKtLR4Q7xuYqtCrg0UWVNbrHtsjvo9xC
STV8II019jq+q5cZ2KKgH9f280OVRLquT+ntOCzDI679kBzt8+1mclK7MDxdVb9PJ5K6n/97zC+y
Bh7ODXugfhV82doePIKBJJ65mw8oTSUbNLvUNJir/myyOAHKHwRco/dsAZznQtev4dBop0SvTWJA
y5YXQjCQTNWd7DNpt+Q0iLDFci4FPxSkVhcE+4uT9o1DbX+m5RKMlbO3aS+oZMGNoJfwOIetZ0r8
VBSS4i5ow7+EUIabmx48VLIdAdSbXvr6v9Ecmp9hFop3fPtn/HZNI16h5ZWjGyGvYrKkHjcRr57o
APyPwhOSpMpopGzuin801qMo2D9zNdQMVoVtNcknpOhqC2nzPKMSAPcsbomp0qPHf11D682XhJpY
ktGdaCYCrq4hPL2iXJWNaCjCDqqwGfqAEp7Pm9WIZ0Yv0wvAJJ0RWzKy0eI83alTsTVAdBfoP2On
6Tql0k3KZrBPqHiE8N312tE41AYfepsJ2doOmGzI28DsgCIgDE0iCYLPjE5JtSh28V84nhfRsGk0
OcdL52Q5ogfspsQqLXQw2voudjfcs7nVJCKCwglDwNS0vRSCmY8Ic4YWWgm+TynGNNgN+/+oDXqH
7GH/RkRlI+lRQX/7KYVP7V2usw2+EZ6r3cpRtkHfBU1Dg2Drh4mNCa6obfT0QLNlOHX/R3pxcV6P
dOdZkoIgi+wCT55OIWsncB/fJD7IgR+hNcVXcl9MfjI5DHJrxYCgDUaJomgRsdm5OJsxqz38uYT6
zUlB7cHtDL7gkK6Xny6BNpp7whzUCiXpA7iWCiZElGLgAkRxKFwQ9vJsGbFAgaHTu97ub+jJu31n
A2HGDb8nBd49l6V89Ecws1XKr4k/G+bqheQ0JhvsJNZX+/3Db2lyXeBc9TIqRhpEChszvep+W9Fo
8joG6v/R0xkW9Z+wsdQLveQj8wDL+JUauveUmzg4FufjUNqcD48zCZqxt/SYvkaBF0hVcRE0keFV
yJ7odqG4HOnIXnVWMSdnMfL2++4RxBuVx8ApUcyPPP/R1q4D6rJlxrDdzLKMB2Aetk4u8k6MTTnP
J89FuAByZThY9BmM8A2agjewm6OBJMZA0hr84cieweVZtxG1iHgg5nICcmHZv4HKti0EmQ+CNODS
N7NbryhEsRlxJXwigv4dwYZ/s/WzJ11fcK548lbnhzP07NV6PsTZi9WT9CuntiM3MsDUc3Zv37Oy
A0ZJTsLfZl4Uln7Uafwp1/c3oQCUGDh67m0uR/8/jBpt4MuLGJbKFYbXZyi2Eotj2H2Deq91RkuE
54PD6UWV0+DxNa1QTjyVCLkCi4mEMmKhexMZ1G4HpQs7fpiwlO4XWRV8FIAL62nUGYyZCWc5PriT
t/x0Md9y9Fkl+Xa9G4aNIp+z87WGKkY2S3nx2+dRKWxfIGk292UmJpunMV9u6Bp5k7YJifpn9pu3
3dfO+ET/zdNbrrwOieEo7LKl1jo7YMNfG8wQMyIgLFYTotzhPqZb0GVEDoXjIFadIWKY+cQpoPWt
cocFJOB8MXTT7jBKgz2IafD2my96dryvC7aNDbrh19fYWaVxahYtGQwGdpOdkV0N6rYVCeS936Yq
raGcmzv17km3DE1XR9I0aAbBEZJqRdB8VYkBKw7/fQ/ok6i0Iv/CiXI0vQdOx57SjS8/M/Dy2vsm
ZPCPfgH8bSW0P/mtoJmzDUyNtOPgp282Y8NNAKr96L7EgOa4b0vIxeMqg9SqhPr8QBV2WsFxfojf
BnH5TcpQA/JoHeMGUrdSgSkmWJa1YwR8h6vrRxvSlCTviQlsFcELAl3SrQjY0g7AoZ431KgfbhaH
yJTb2QQFt1/x01dJ052CEhgYISplHy1yy+TGQoA+vLI2Pd6uUC8LrDHp0f6mZdeCGCfmHT8HhF7g
Bn1EoiH1nSPYvVjbyAWXyxubAEn6Wb4OXuB4UzJb8yqRQ7a7O0O2PbP2Y3YpD6uCpx4MaIM6FF0d
w/MamEx/MHw/9qu0OtixrbIzwRMnzRxi4JEjO72O+fUvE6ih0hIhpmTYQfeOoRUNf/XqQ/Jh+Gx1
PlWvAwOehbqQgFV59k/AzB/zHSKc9RGKUUbNQRGwP2XJL89EI/5yyHbR9osZrlgd8hq4BzRBBsiO
zKkvnAxJRTxv+MYdYQmzlE0qpmZa+eyobqGbpyXevXUhL+rVDgIEzUel8QEUZfPvKF8EtBcBXnt1
RMn/YUpbzLFHEPaFLMgv4d/0XJDhAQw91bmeg1D5tJdGoYbKlIxcRSJ8RSXCqc7vfCwpvjmPqQcZ
q5NnNk3IvtH++xU2hNT6MPp3i8Up/ylgW72EoODlWZiLaBDCFW8evshV0lXBXRpHsLSlY5rokvbH
HHWMce15/bRZCGMwePWHXuxTWIP1yFYGcaChmMUv5ZLpPhjWb6R7lAbGZDUkSi7Fbe7B/Emo2PK6
bQEa+Jz2Np93pBuW2kbWz2IGBc0MLrOnVj3n6d/22vamFq2msd2f/jUCP+xxyFuiaxIEp25GgxFe
Bxzhf8w8zJDAK8iuwUkPfmyVr3gISb0mTBmVy3qWUEkjFzqurQXzXLt1LoNiOmA1uzu2HKJQZ0Z+
yO07GQsFyBav2Z4ChI0BKHk6+p/sX11xtTdFrYAcw6xisajCMwCOl5j6QExBw8YiwV5hW/sCli5F
mNlbH3v1EapwTw4pBpL4ab0QsL6mY2iN/UZXpK3H9IDYlSd2giusErbGz1Wzz4sj6+RNrM9BrmAc
wVQiD55FsEPojfqtsj5QtSPhwwH+QnddNOIsMqqOsA/u4hA7Hn9Xhb+heGRavdMzJWTYKHsjCizo
/QzxnfJPWHp7DmD/RLPLCjrBNuSwdxs7hhFMub5nC9M4GSPU4OvHMoy91cbkCeOCQhTf8/goSiR9
8WiqWxLBhxSgpjiL4MRklLNO9yrnz/ne3kbr9eSkB6HZvvHS3msNcfSvTP3Q2iMqbSgViX1FMst6
zlGz7cC74Ba6/RpHgKkztdcDC100c9vIQRt4+RNlnRRaXQorTA6FUe8YzpV9F1RjGH+oUq+uYVWP
NCUUAv9e+mDZZw6A/bzVR4Id94vykrFWabbbpdSZmBRik1JNvqdeBxAr9JC1KNDYkUSAhVhr8Y/w
CNPpbMF3QVRGLlMj7P/Xx36a9WbCgQWL6EA1Q/PS0wZZeyyFheie+HxmpvX2ZmuZeponad9Fw3FL
2NQWyUdbdg9T12BM40FC+fOZVMl7Gh9s4NjlTkPBtLg1tZdiywiIe4frXD9el8rqTHy4CRjqiFDy
HW5pvcn/Pk9Mi+zv0h56ymZLM4MT4gGiu1OhEmNs66BqFmmuL6KIBUSbAhPcDX0eYxCWlq/0oMmK
LeZfTmr9GRghWJIKO5DKhu86ZH/mM5vucOOlBHJ9ez9wxWhNqEILfydcBJmHc+lu3dloOu+qiA9P
+HIw7BdYf0LZRQcP9jYF+FgxkeXdNvZLoML4FH031KGanqMAzAOBd1thEFI0rOJyBpGXjrk5uNJy
tl73JPSEJ9zRSkhFv6S1BRvXR8goK4eTlaj2kV8OO/aQonFrH/ltBkW3kstK3nX/MfKwI+yRDS3Q
8CXb1rYMewgw8xsahL6gktvpKvoRnRv7N6S9148fiYDQw11ljmPnabvFG1xdD4s0Z2gL9yINxOQe
+p3/erEsVf+5wT9Ae/ulro6rCdbxi7KsLqcoW+SwoVg82DlUmAhA2y61yK7X/fgF6rSoXtarC5Ir
1VDEsbtYYsbMhoUvmx4eEHxanic82xGFagPSN0MCUHRA44u+Yvh8Vl6W+p89L9mEp06boyA0l5lM
HVaDlx1Z3rq7oTLH3HlXhR1nc722KgvI09R9lV0Br2I2TMDVTax2qKZQbWFaCKXfZpM9n/TEsvAt
4TRoAf6e/OsDWtNg9kQ3bDwaBEBeH/hd8QTmPE9Dpb7b/0espkb8j1H+c+tBuUAkDm7w3WPDRu/b
gkBqCepernwdcvOit2YBdvbjXNGrooWbpY4J00gbXMwxlgIi8hoZnfBBNcLdF7LGs0umPSdpEjms
E7K7Jo0/TLStBxYDACjvnB4jkSiGsShf0lTHAxcls6IyM/a0PFphgBgXa6R0WxabxKVJt0QnYEGa
tkAtSa6ePOEpwRA01zLu9i+lkQ+SHdBDfMba1BRxCX3zLA0O4FBfpFgeApLGIM72UwLbtVU31AZi
99Cyw5WAX6k9ngKRtFUKsQVbY0VzDIRt+d7M/+ZunD7a48tDnvcFLD/KHMVuwuXhOzyHLwN0CqSH
K+q/guXtBWiyIZKrQ0VsmcsgTqEzSGa5U4FLNugGsDwPOIN4P48hHRYYnnq8gn6T5r0IFhl5Na5u
UnZx2G8Z0GylWqcmDRUO+y6Yj/KVbqVH8gzrNNy+oswZwpK+jy/aiLl1wtceUjUClKalmLaILk7T
KXVKZgRZwBjplXr8L35YLIZrLZgtNwag2tCxcoSSftObB5a2kBsJHZg2UA4hRrQIp7pEvU1yS2Q5
iVKMwZP+ZoFo9oPpdxMTizX658K30yPdu2Tc3HcKGJwBeIFakNQJVddJ6Gpevv4UF0PSn9PEjt+L
kMFnn7gJFYOHvGpcLB9EcM4jmRJ8d7Doi17u0afJ2RtTx4KEQnN9DQdbQKH0LJnRF54wwUuQlVxn
IsqzROyQE5M6K7QBCv70d8S5FPZapDphv8611zNzkwLC8ZQz4qHW/1cDCPZhFu2Yhyy1t77wzuCx
dQySe3om8fPuOJMaAiHar2tiPq2S2flXk07Ir3S5tL7K0sYHXQXcOwQ5H0f71RjJqcqOey26f+v7
WWrkibr4bHkWl5JlpqCQFP1rlFXXs6pTGw5wbisiDU+aF6t8YZtx8zr3OhfvsAnj6DF+tHJWMAk0
5Rh4jFB+b36QbG6yDqUUG0uGq46fWeZdK/xhaB9ibm6AlO1+Dch1S/IS7N1stVbkLqzPEF8K1qDL
eYWM0eUWOqfHOcWLeVzYXtUjN+lRspNxRd/5DXQ9HakQu0FSiSlgAm5e6CWRMdhW/wDxnCsbOiO/
VeiEzilMlMFFC8Jc9QbY6l3d/rs8yZcQd9vKWNBik2dmNcfrHsOAAUfDKzamS6x1k7lbKZOfwFUl
4+W2UGleNMCmFcPocxNEfSH0qyKlOdOeSeVHNuUOgnLdFCUO3zlBhZTZv/qeq0Q6YzFNUg33bu3+
yPH8ugryXDGZ/qhm4QZJDFMuLCkl+dNgj24Q9O2sxohb2XR9og+HKKxCHN7aBTbZ9W3Qb1Ga1REk
7n/YAAxbFdKW33zE2llUh7ZZiX8P0d5i11LjCcE/moQo7xnX9SyuFPZZXweD0xTLIoVv9UFNcxu/
DWzLlkyaT3vX98dxD2uHbhT0Wju8jEeHnffh2ah5vr6A5tv14Enu3hlSDEp99NkNCMDism3fXdUN
B4bzA1qAG04CQHgpD8cf+u7LUHryDxyZntGwWIy4rC+xi+VXIzfkgqdxIYlXT+UwjFENHn6lHzxw
ETPK1ny0HXCpvNdM1b1mgmF7nEfwdMiqrxNStWG6+SgKB+O7K2kfufcHUs9LQT5mm0gPhH3wNRyt
bFvlGU6ZFhT9Ldy+utJJu5DYCTmc76VWdynZUXj+FbWpR3LhnqRr/LwVoHRqHxjf5hrlfX40TxM0
QIGQ7k1lBvn+tNrE3MIw5HpAky/mkB7oSP6VGs+Mvk90+7QQ7u1NQE08pShb7/ai4PzoTu8M9OHg
Kf1N2K9xzSw/VvL5oCRLfu2b7ti7LFyAmHwNXKIAqjL/aDZ6SmwbTefTOv8G9QwWodpft0qK6PQ/
t8HEajRrsiwaVdEnAGw4cIhI8IVwO0mmzcn+REKOU5FBmn7cP9II1oOKaJCDRqNvWJ2YUr7InWN1
inQc/JuJG6g6lkDIQnCxgCkBefSNMtjfWHKAPfIc+7YmgBaKaoYAAXy8qV2HU68EstiMQO788NiF
cajxnDmeyHE9kezgrSNyBHyzY14OKrviIiKCK7lKp3e6wWB3lS24Wl8qoCa89hDIZg6uhekz4tHI
41l7ilZA4b5z8n3F5bIcw8gRTouAC6qF+4+RmDZN8X/i47GWTqS3hr5bj9Mx92GwiuGSTVE2GZlu
BsATIyFx5Su0PAtCnKa39BR8dzaLcqfuVyTAH2NGWBBT8UYWT+sUl2DU4e5L03qdr8Fg/D8RqqaI
WN8pceqWLPj9ilTXziY+7/O/q7zpnziY/Ted2LzfRqeJYhGVdKlyXOy+wCWwCXVVcjACHJESQeHM
nHzJNXgzs1Or9mKiySugzj0NWTkSsfZKWqHB0T5txyAJPtQ3MaCGbXFMfsKwedFlltcs7kpN28bX
2tj+uwJjdqpbTFUB/z7e1SDmy8Ma+RokR3aRAuze1ALUXKW6i8j46KNGM/oL9bHj/HFjavhRgHbD
254jIFqh46j5k4NOBUS5xqQ2/lSEvWPtUmAmCDbD2Db9elzfJyZYSWSgYblm2v3KgWOKckQmD31X
oWLwUoMPWm2CwKZO+GnQWKA5L+r9HK6ORaPXf4a1PfaaWx96VMvLzLBQZEOZz/3OQimJYR2MO2S8
yWs0I1vlFLCyRJ21qYANyg0OE3lexWx50RhecSNZb2WjMwLmV7nQs+Y7b8eEqqeMkvkNrah/azM1
VwreFOMScuKOlqUrvKEkbirdQMcEjJvW+KEcMNKyzQQ1PlrHGHdry1OMdOfdodroRogEY7lYPcf2
AMScyMX4l7TD/N3NzQoBXVNqValKDQhTGu1SrTGdtCP7QkznF6wBLuj08a4AkgEwItVorpcx1CVN
qg8kaVI3Rj10jRusHguBPEIl0xpRZU2ailK7CExlz3ASWpTw1JYmRXpZgxvBEsjmCNHvaLDQYB9V
ZBxtQ7S1d7jGk1VmFEhhamiI1Y7zcnsY68xtb+EdQm1l/WV3AEzlB2HNQx3UZQAgh6HQxj4ZR/A5
hbATVO71r/0oApE6ekz2EfsBFr4zjaBZnJHzJLv8Q90Ab3ohiE7OGo800s97v02vyAAjloe8RDh0
GkElfUxrR1wa52aALOPadKgKnolGBKMxgAHAiccUZAf8iRBuwyj8idUvn8ifWR11uy/9qPN19HIj
Z8wYQ2LWpFQbnBKJf5O5UgTScIGSB4bqC3pdNWbI5v9PzrSUj5hJBzZjmWWu5a/KRmAK6gK0rO5u
QJrFDHZWgqgxPvHnzXoEz6ZerLuOhaD+8Qqm1dDySw3Nr1kYFkrOoPeQK5P5e3E9gNGPs08L5qXN
08JcnihBSHWR1U684bT8bCN9k1BpDeoVgd/XarWnjTd5t6oD3OTCkHsYdf0g/ZEGuOLboZqv9usf
D/vH++suHZ9gU9kw7PGo9ggmK/Vli/smlrYSSMz4uwoyC/ZegDyOO+GE70OzFk0Wox2GhGfFR3ot
Qd/VtVBCD8Xy+Z8PMhpRgWGLvuC1FW4AFu7jMK171Bd5vjwsH90QngKto47A9zE44WjyuH9gmlMt
pJmUuXzEtTX7E3QqTvDFOTulztNaTdXdb0vEPlZ+ws5TCiG5vgLBdyp8w/BSmxUllHuOZM+BIOX5
nEMCcqu+F88MzmZyEKJPONjnDrf7JRAHaEuc2zrCgDA9fFo1fGre11VuCZbPQf04hVggfYMMKV6z
1gjybmuZcwXHmfH0mDaclwBufr8o89iD5/kpLVbEbf74IJYCw2q8Ld1T24Lmg6jf+abg+BzxPXSJ
+432ooj7ttzeOY7IXawVxszZl31V3iBPNCxBTmJWNWhq2jAaSGFvWVX/3MNIU1FT8Q5VTL7J5CuX
y+t/6jTVN+bqS/IVlXBIb+d4QTx3c3h6fkLEbMnjR4JJRCUEQwBAG29ehfa7VSw6pyXx2p9cEG96
V63JgnVCFVVwxYBryTWyuqMdaoyaKa4XRSLLsn43s42yeXkFzmdivf2Hx1VAhMgLEgjLXflAKWep
tKsmHOKveBM3fl4nRijxUzQhgJGfzXMR7KCz6MS16PBtIKMPDwNeIlbWlT/rEAby8vwY2Xx7ejG0
lEWthjaseA/CP0kf/FtW/69/JYuRIPzDapRzhSeAZm9n6BRpxHKs0PDpQQz6sJG2l15IPbaTqJDy
IDsTVlExUu9hqejZ93HZa0P+SjXDN7VJXmD3LFaLwLsEFJ4eFP6U1/Y8is8p7tz7+ffOwswHcn2N
czQzZoRFhSzBrgMyC9eN597u85QShq0HvJYV14EZiy/2KWFfFrdgVjGKzMsSNJ4g9wZaHsuIlNeV
o4j7jkLZAYGXrc1sscjwKbQBSYF7Kv7RSw2kL20cD61nJBgOn1TEn9M6bFqABEQZr5sMXYXolKPi
7YOyhTyPG+PaVstavgAVmN1ElLwvmIbvYnokWhf1CWy4ttrLdrHbO+nP9bZDhX3xE2Or1HhlnHWQ
sPvTmw0/vCX0aaaPF+IvA/iK4C6Q3Om+euwZ1CtB7NL4IX1hMOv4Iy0dwCmdH76rj8MsyOvFzC3b
15GtXRGAbQefaHTwwBVrBHeQJQAdMtBEYdUs27ed/YA8mJ8k/unR94fEWghjlMJJn2AzwYLh383g
bK2YZgpDJasZ107HU1wweTfrL/5GFJGxvF1/D4QiRkOfR/F5dBsDug9KlFyPqHod8mZ/eA18yg2b
yrRDUm7WFkIygrzZzttY0qIJvemHl7z+DJpWA4ws2NmYZkdFpyJFSFg5vhJTgu8+7CxTXbtHOsi6
tOHPtP8Zy/n6Zu98Rk9C2apsuh5RvJqVAi8xOihmogewF/RzaVCsHLWZpVky8lul26S1eb1je7Bn
QOzUgPzIKVs4zaWqxvMUwX3GWhMaaep0mSKld2HzhhQvRJmvYtyPu7d9V6K62G/7AHMVy0OAKc/v
P3uiOJnaS6Sy1trOdrdrnmY242Wju8l6QpcipS7ho7/a5ZOGs8Csz+PGsk2CA203Dm4nNCFc5V9a
Sx0Vog+cvKga24GcTnVZb5c6WmyUjWmpT+W6nVTH6haunwrv/uNPJLGjOqzxAy293wQEXIcCJc6D
I+Bkoj5uRE7X+BS81TL/QtgEPhGcfRA54ZQaW8n2qvhObFhJdZRxgX1AUSySI4gSkRqlw1aWsy+j
uoswsaJqtg4ZdUNHlgRjFi8UQFNXtw656VUYQ1Ld9SdR4qJmQGZ6xAmnW+WboNn/SkkaBeUwSOpp
MG7sKQfI1O1XrHh9nQz6Xq647seDIzQEzvNCrGuUWBgwirAxgHooRHEHAdIS8kOwZmicSVXUkTcL
RxQRbxkCasSdcDKVMNO1qgIolxpX+7vGRwaODfS2JEUUFUO5h5YZJKMMp8341+q/zgQcXg8AU3BX
eemRNFRPOgz1k8uWkEfvVod88iFX133IbXkc6xqWQh3MiIXRGxiFNQ1xEMsmT9+jWQZueirGn8ZD
JQancu5qC4+QefDVfoTtk7T6S+76eMI1v3MyKCaIfv30Fi9/NQdxJGxjGMAL7YAz0L1soMUQhnCL
v29B0JC1lImmEb63RsiMBPY6wTdHbhcOU8D5um5vkNbqoqjN2Uwo8YWM9mRLBBQ58ORqrlmtvC+C
DJvwdwM3hkqSQlHe7SVXWBU1Iro6xuYsA1YOPp2/HI6I0IV+r3+vWN7tsprH8RZIKXS/LtLqj5xh
w6EF2qu7pASi2AO4mw2wlopEBrIf/A4AHWi50gWuBXdqHORwlN6U7PrzYX7z3T9e7RwWKFlYrMZN
BquUG4P1b7Nhd6iXdRUQecafm87V/UCD+6ONR/1sg8wcBSpkSgZDf+SyuoPo0ilVR/Y09c4mm259
NAjXCyzDlK/yWqr2X78EK9jf4TmCyDm4qunj56IUBYWBWV5GQUie8uN3C3+21dAirPx9hUFIwy1U
gF+6Jd8kH6C+n7/G6qqgHO8n4ZOgQILVhIVunX7TREgvqqIHTlA1G7wElN2U9WENCd10Oeg08kK3
TnguLUpQhNwyIZ8UDp+49/J6XuY8bPN5GmcvQ9eW1IMYGNtMIrdrVowqFHCtWaFoUOWsH1EZZyF7
g2vMajPJTsovt2LKFst7J+5Sta5KqR6QsLFPwPx0hJFVDwIQbpSphkrh1lYazjkK2ce9i8zcd7xf
XNMXSFzrlWAHrvqJo5SqbN06MDmatffbOVTCuZeKBue51QKf3ef02GWOY9uZKTixk3mX9hnPnEyG
qUGTO/yUEYBD1fBQYpf2On8Sr6uhKyVkmwXLA24AuLLpFFt0SYlbGJ+zZbyAfz03Co4pL8DSB87N
6LTvFzgyQ/txx2Tz69QVVC4mGwfJn7+iLyTZ76qAI9JeTpjW1DZjrmyEkoWiFcENzrvS4oL0z06Z
dE55dq4g8dhVsDnLtZ+eEVCDb2zOA/3U80oDsR8CBX9/buazDQAz9j7/LF5hrrapyBKGz5KZTTcZ
w+vdAUNfmmpHsVxBnTaCuy800mT6PmkKYIGtLUvYq1tF2usgRfXt1USNI2klcelb3zGFJ8G72CUw
VVQhU1cHv/OHSYyfCpRqa/cD7EThWbxXmNcEtKNnMRm1SdRdlQhbscD7+saslohg67o4ng+QAXS9
o/M/GaLjHm3qcfAAE3FUv3WQzdQ+miOrM2yW2BgAF4+0r5cpPXqj9M++LWlBPjms83FfrRokxk43
gfmQ+wk2HcKSjdlilgVZgL63zGeiibdfnEN4mXqnnNnR8qo5rDnRqyW2KVWlqUFKm7xyAP2R4p/k
/YnzE/zmptsa5WQ0wawt/XQIjdwx7RY5SCOz/JVPW4fzufVoJzognI2o8F+Rxm083fid8hHcwR04
kc96qJTFhQFZvRrQK9BNney6S3S1AIPguzOwy9ME8IfqmP6CpZD/Gj2dW2HsVUgK+T6BxbaNziBG
hwjoHaAMVw0BhjxgHeC7aEfncb8pzV0y++vwi2f06zB8mUtxoeQsmCFNYFJU3JtSHzGk7GOnw8rd
L9jm/SZ5TpSdnbRu7+UqCqZjZupkiB88R4InixmvoEYzUCb6B9i74lQIyzEfvTokogBdQJZn8l8Q
SWK33ail/N+2L2kuHIIAXGti3nGDtxUE4ecSZL7axMRHoAXtj1yeQo/6gsP9+ysJ2oRn2c6d3ztL
1XnM4sVh/83uOMieYgm4+ReP0E24Dk0yE4uhiykLJXalt+l5YY86wiHQUUxHXD0X5hdXBWuZ9KqA
4XZrkP3bS78OH7Eq3x5QFg2Ugna2IMNXoO+uQtqxIiQG5XG6pCgZSAKBthX+3B7GtH+nPPXxWb54
Q2YogmdlvZJcZxG19ee2vJgCw6SZmTPCBurFlbqLw7TYCBQxaFtqK0jVOxWIx9n8u1dHIX228HG9
2aHG8PC9B6d8M6NM2NE2GaQw/vbf1NWdjvKuNBDhOMDNHiTkM4Q11o/60knXK4jJdVgjC7eRpO5p
TA35WJYHxyMPYbKEikO1L2mfn23s4NyG4XiowhQX8M5f5iSNxBPOZ1xgi+fCwn7qZB6xzvYaV6Da
OF6fIqDXlQgNrUiCTcVcBM6Z/PyZOMTVUl/+4+rBAqgs+eY1zhTpMBsKBJJ8UgZoTpUeBjuGf0B6
xdDBWQr/P78QsnAK5bzBWtRJD1jT/TF+n/soBeWREDJqtYxXbU/AT/HNlFSGKG50Tuf6QTtc4h3/
26FDeMYD0ynNNv92FLguN+Pbwl8sQDDWcWTVmM3E2mUSCCeUZGN/CeGl92UzVgCvRik4GtrVVtvN
PIZtp58uhlYNA3UdJ0nwxWW9C8lSYLwyMDPPXjXpoWKzRFUhLYlU3/Ls4bMOjraOegpPmpj+H32T
YGpNifX5JZ1PnGFyuhnBKAsWVBuO6HU8ChOYcQdenjei5qajhmaHe+1Nw+fMtp3EZiXMSZt5wq86
Kdf+p3pQHD49XJ1RAV1hl0rBQpKbxuDr2IIrBwqd6pN5u2aBPdtzgHx/KqErEllwDpB/ks0BPIsV
FFppagiXDoq/VU7skElR+tSiCNkj7JBf5oggzUBkra4zlOhDtyd5YwzEbmz6QmR5MnRbSEuZumIC
WuTtZycU+sgpPyEEsCrTw6dNFZoxZh7+Ckn8fA1T0yfXFS4SueuZ79fn+2ksFRPf9drAt20D9oRn
GVh1E2yl1Bc1r3xQR28GqxlN32Dg8qEOFp3eWC+Pu0HGDbMDSryknXIOQLjqgYIKqc1+0bFyCTVu
Xg0cEhH+GEQYPMwft6mlziEoq+9Sb5SZI2JkfS/0ulbT5xKJY+YC5ZeXFsekbULpNIzZ5lCC+CV/
cStw0rephuMG+n62mrRmz4Bt/SgZgSjijkzNp5JpCNqUSmWDqHFSPDQgn37CCWpN6/fM4TPw77bP
9MZdrVjkH1bhpH1VoQ8QNQlODabIZGi5rXpfZ/nKXGAs9HMlNAjHGnIyFNd2tuh/NIdREoprYJyL
guqhNNUroqiQR8tKmJow3DF2rtSNQQchqvuduSOMFZTMexAn77NGFR9w9+gcRJZNXudAUcB364qJ
nLyy1lhaLiodVr2JqMHgYiitv+DgjeI65D+lezhfuQ2nTvOMDhFAWMwEgoK2OB7jK58Wyjrpi9Y4
Vj+dJ2ywXVSVhGNsMsksr8XQF2E89QvZ9XNQvW6oop/D0iLVbbAf3eDh7j1dHJJuR403P/+wlJSl
uY56a6Ga52I8a7VfKg/KWKo0HPK1w+Ocf1NUR880VWPul6IAVkw7CO3kPDYoe2QrzovvQM3Hm9Xh
BDaYQ25q7KB5MUzfmU5O7fi7Hb/KTyKkWJ6/pnwlrFL+uxH5Vs/i1zLeKCLgl7UGuX9qx1UwwFk4
feNTTBsgBEMpsD5TSocWNltWJtfxUZLzJlhE08Uuz/RXUdyiqQqjFj1jcQHSANzKFkOyswltzmhH
uOnLM9LQutFfDNxAZ/P1A94waKgO4Pdj1tiKO+56/dvyHGd83l3psxmMwXeuFnvnRm8+WjKyK/sA
nlsNKavE4lrOgWZcggvjvSIwLaX+9vwuStDgtXAt4TnC4L+5mkgtxJSBDD4vqlvWIC4r8M9n/Fic
ZBAb5UhAqYFYAJWWPa30GiH3iInCGa1G1FgLVo/2CVpZcGrOp+bpxv9+3fQcbfKDurV+IrwJD9X3
jPzIW97uUaymBZU35oyB6BldsJ0+8NO6oohEkYVx9TGgqs1qNLOyNbZOoT/lxICYcUY37d8jf3PG
o9TUMVv+VfNSVjTrRnHe008HHfdCQhoswyyuyOei7uDwWcTeshs2qhWEmWZV2R+2G1IHk0cHjj4o
8satnaVpkuokFSalW4G++KnRWotxSXgnTSijGAOdpy3kX/rmlGLKzbbp5jRlNOJezYNx76Jo1W2/
PzXDdnMVl2T4ZieInni3ixWcysGnAvJxl/2uMUumAaE3Hakx/oTNjPvOuUqOBxfeingR5GEglX83
1/Z1bW7PRpPpGMMsH70L7PjgP4QMtlFKX8nzDX79lndwRUQfwdPnRpCYGIB2kLupyPBT4gSpPJwq
81p1ZYx1yE6gwnnaIwexZw06YNWn4DKMJP1Hr7CbQyJHuCs0NkTOJv1DrT5faAgj2oXKnV+l/c1a
EHr5iFTqqG+uw/1qyUhczq5dqZWUpyxtXSY2KA1Stp1klmVtGYCy27yA/LLwpqdSjHjysUEuYaBM
GahZxlVdpcNJ04FscmtTnGwtuyVpHIu8myCHk/6xOi5pMR0LUxDAqpWVd1Yj5zWFQ5bkVet/DygT
1xPwXYIi5A/nTkB9zNnM57gDEPdbEJIZF9rqcDHcGHjIM4ccQb79KpOtxD4QqaAhzwezzypfNpgH
M5mGBC9+jk8gp8nIq07a3RzBfzMN0EM4ds92GD+vzz0N2HiO7lI1uQJhZ87XukvrljC882C6Tn6n
FEAd22N/OT5KNP3to86BuJdDb3zpZGg9MX7qHBhJvarhl9rzD8MtakeUxOdpdN+8SmhM9gfRyM55
5XbDrAD5SbMi1j6sntLMUgyR/kIl+jHmHtHnJ2Ni5fXiHCLb6lJB9Yk4yzmSU2mmFAxYWuBXGA1Q
ZFfHKKX8KUQxwzmszKc5LUdnWYU2rFFKNpmoxoK2AZX8fNwJLlWUIWahlMYWYBpOL4CJsp7cgpTD
pga39YdR6bN9zpq6fRBjjnzeoPtUd9uimYP2ApLF+fdJfahufB5tj947vSZ3H56Yloits5Zd6g6l
kXZSi1o1rrHIZZFmM0QhFXmdRwZl2GJjfj8cwYLf/GPchJj873qflYL+ZM1eF9D7YX3L7mCw+rxm
WGDcWFL4N0Y5sgPH/GuclMZ1pSHUXITuEwwiesT229Y/s6ugE+Xb/3Kpsy0FpzCbjFT5lJqPQ7H8
wMnLT5HUrSpdVlprFoXdPxC52k4u8mUmthhkw+GehuQmrgl1CYoZXhEvPnC3vwduMDr/YTJAHVbX
Swi+104oQtm3VVesnc0n++k+GrI0uP3/UA+SLhmiUBoEky+xpGq26v6DoFStlWwNV5fIXJylPFYm
CtheCe8nDbkxK4CPT+H1T5YdxwGGhdFH0ojZdUkiQmtXY0Zb18HRYc4I+yyBbnllLwmgutHEzLlq
q5RAdvIm2MDh6dQoClLwFo6hv2dvmWBlNXZ3RVvcOM8R5hKzJglBocG+PFGr8P1IuGNENmd1XM89
NHG/HyDFtdWo3tmWQzEE4+DJ5Ty9FeZRzRu6aXmPcOQ91xRBjfmvOZzCOrSKIjeBXPoUySQ65NRF
saczjSTcaWahvy92BjzVmybOiuUhGKvwF3SI35hM/EENmNF801gV4vhrdp/X8FxPltyA4b/3ZMBg
WiIeoV1WBJd6vdUGLin/f1eAPWvZIsFDhK0+cvxgWIo0M9v9/VejjRtz/jVEeFJfe0AIOfyT/kDj
Hjv2BXeJ5o4EtnAJrNfN8YuFcVmyrt7DJFGWB2NeZO3fkopI4L8iWJOife6+VKIcs9XuqR6C6+ph
FRqu8g0DEcTLXRZJ43PBW/7dczf3TR2VxbkElT6n9uSERjdMBVqs5bzrNrFLaBjb+rkTvPQSqS71
EyVTiW37JbUv4rPjGta23kcBlrCA9x45u2q91YVfVKEpKo0LflrTOzYVlbmrmof3ZbgOPMgR0Kg/
mWII1IPnoX9b9oN6iaoPKL88IQAHeVYkggNdV3wORwmtAeAjK9Ny7GCyZZ+PEHDDU/Q5kte4FXJt
iyO+0/hVCXg4aGRIOTRSsO+1eGmXs/PNeY30S1qt2x+4DucW5B85mRqXh+kJ72OoIm4kvXvTlkbu
o7tMd+Zn2itkhcrMnlAB+KLi0K/K66xYa24BCbimHgjHKXzPqUsBIJYbiafT6Ue5hvMM6gURPYxp
fS7Ms9ihgvSvXDr4HmdpF4tvIAp8gLkyhghzH9B/l3Mym07PA94PGfBDli3za4VD8Z9IyWaMR8z7
1Ium5q+D+MzjXzIAYJCABWlsb0afIMc9kx2b6LAewQsBAgxAEYTwyP8BwyGQkzWtjpQ4rYt2krGq
FyRyJhvlLTAVjdDU2wOZRIWxgBz+5ql7RlE/JOnMCC/ZEebYAbxGFh1xN/teLzlL7SYejkKT3xep
sHJq4dZMinvAuLd+1TDQzPZiE5q7k1ZGsF/w/dxFTxQkJ1GG8uvRAhO5eVCQ5IJRl9k9hIiTb0zP
97qzc/yCM5TQKowcOV37oC8EDQPh7x014BV8RjtBbgFPVjl69wLf3v3zyogdOoEcuscAePC6ax2X
9x+plfUxZDpSei65luzWvijd6wy3Zwzy8O443ak2BjHE2NnMVhqErsQDrm6McbbFAzAIL5l/UW5C
yF6/v+Ntg+77XQPtC9WWypAZcRbmCihluRDfElmz7+2yHFfJoghyeIxjNsOYbFXYfU7fMCxxRXdn
I/JpZXsdgGw4rK30QFoBStfUzuISoynrDb9b/rX585bGBdXmyeJU/Q0NlqrXF6Fr2zoLnFZtd0ue
49r6RHaWIDNreJnN8NdabqoIiw6WFYBKtSZnbAdJI2xhRN7mToas1vOXzUBdd0VrH6s2l6Hf/dhE
xpgnehVCHvFAgdNRO7FKD8EANu1R+waMXQSkloCXxPLO4pNE1Fg0BMBCCtxiuY0UEvvmCLLMwg+8
/CteHjaic2AbtAwLY/rKmFQbLTE65Ko2GAU6xSPdANVaYt53z3O4XtEd1WmrUExsz4l9tRnYQjFJ
q0xNUUYcG5G+9X8FwgGPh1jCqXkvezAdUF7k+I9PLdFJ/aeTQgheGuVPuzPM8h8+Gnl7vD+ttlIS
22raViiurOSPGLxzTUYmGNRZXGadfAyqjARQ8zWTxt7XAG3RCUgJjLHsjcSTfo4mLPAAHtmP8Fmx
H56xnSajlv6BH6IOBZM4H5FuJdfA1mG6waVdt23CQzMZsifm1v2krV8sq3UDLOzzxozgzSt5UjeA
Rywtsm+hCDCrHr5ccjGNMggsql/ajRHg/FXM4YSQHdlHAJ+lSmzycd9lkFGCLbFe+e/sm2Ch+k16
Bl/UysQUrvWH4IMXUNw19uiP3y1NrfuypeCbwtQ7pD0tYYszuQ6iEoxdds/ZI09vWbOfegLXIGql
/h8khnFXUnQfIiJSsg5TEa0vVNLJxlFua/ZkNwse6PKV/uMYlOVU66EC3FaZS9brNUcyWjOze1al
8peduodRViqTPjRBms1I1q4pke8/hyR0UYjw7C8OPiIT1aIwbCeWy0KfUHO6WlSmGsoFkIZUA8hx
P9C8Z/LZQ00/nWG3wlk/IiNa9cD2hwg3Hx3jhnB1OLIjdWL0QfXpduOHqs5nj/LSpl/UCSIifW8G
Ok2th55L1nM+GQ6v5CAL1a5Sa48ZB4Q6HFrsjyH6a1Kyhn0MevrAcsRRkBPbfquvkFtUiGUGfZFw
25Xu2a5Wt7iQ4BSvkkTUlvqHJzPH+kQKH0wfpbS/OzAfapHZ8zQKodzpNLajJzkBXiB4e3k9Olhp
n8OGYJQtobg/HHxVD/pAxxl0W6GgKzLBJ9d4FtlbMv0LzRpX5MmuDBNnrannHB2sPhuPdJZ8cyje
A0/IHecCcPN8PUJ+JDoiXyTi0qcjBkknMOB+TsfpCpO1YPYRS+qaO/A0b8ILLt23cZEMlYYtoTyg
V8KkFi9uCOFs2BTbrGNgjDtwWc+3bbgDQyuXRp1ke7U37t68ZYle/J6h3naL8xqjx9DaDcOXkYA9
7aO4QNIttn69EFhADyky7SKC4Cp9s/dVqL4bhjquIkZD00A7c8zAVugwZT+8NwlQGrB4+6GT/0/L
/AhxQxwci3KsXm+upJ1yhMfTqaySAziJdXwfV4bzHc7IUKIb/O+r9RBiRoJSoDwbnRkEC0WwPgZV
M8oW4qsb5NOsk0yLn2oB3BpJB5s2U29rJYyDSsJ8uQ+gTpsp4RSC4TM3Xe1y7HyKWAzRVM5icXVn
xvlucwEhZb6n1DzyAdFIcZFJ9/4bxexveIiVGe2LtokSepm+tVSGdX+puYxeieTLmGJAjAk6PrQF
6/McdGk6geVJSCE2AtIGGgZKcOCgsp+DU/lP9wTux1UFI7zcdCfXcknv0ioZ8d4d3yulvNPjWdGO
tHdNYLcpDkugZKc3DY98qVeKyFHxmC7HTIObXw/lXdR8vlVxjqPUa46is9XhnMzf6iuXKggtPWVw
Y7IgvJ2M8vt2iiZpq01BfbFRz1oZyv1oDVJVnV84+BcpPAD1s9fB7fTl1nmMepPR394VeqCufPVs
byKu9p3qJqNDdwvNfGBlMU+Q9ZRQ3fXpfrIyT8rqCeBQQgysAKCCoLIIEe1LlAzsqmKGCuP8cjem
vpWDxkoeTmU7iok8qYJQBIr2xH1E0FVf+1gxztQCyl9kwgejKMDAwU9Y084gIZqMw5uQcqo5JduA
H7HF831vndBF0dk0GGRSWI9SduIrIJSC7JmzZruzLGFwfXGPrn2hPkRIR8qDuhEWWMN//eNYEYrB
d5xP7ptnkvJQNMnQdsE0SActXryxjs97SZzwi9wOOTxqNh3h2STKmTIfruML9Hw+k0aykSXvgHmp
rjGhZr7CCOwdFzB5DDWahoU1QJdlowq6Ln9onC3mkgpJ7MXd+SdNYxUEqDMe1NA1duy92jh7Fste
+KZPcizHTm389ksfctN7K45JWhFs7QrtE/LJ3N7kL3HOWxYgZC9QO6vbJ3mGwbMzraJsknsAUciT
r0NYQ5TreSYEY6nW1EhZpLa6kLq/Kw9qrE/rnofPi3VBMUTDOt4Xzo4CdErmdWrai/1Siw4HS4tM
SVrhGsUyqgp/+s4Cdc8TLnsWf52fQMoRdfuQBs2gZDnY58/qnvkj1t7xj0FbMWPYFYfv+VTbkjm2
sSEpApcGciLh5SjcIncg40BDox/2A1Kf/vgBWdkkutH0x0hy+NJzBEgv3NnK3A3NGuaHANSL5Vh6
q7biP28sGXYXalTfzICmiq5ctVO4FVMYo79rHTkYrE9yE7e2VC/xo+1yeWjrCftXOzc7QIVKagbb
jNlciU6BD1DUEi97F3t98Z6wE3AFOruJGsEYnzfzcZ5jQWLCWHrZgAJCwSrQNEl/vWTKe5/gtTzg
CG1Mr+NUFex7XDfiKhxhVsQziCpUDOtvOwmHuhZYk1qOIhE2q9j/cgl4EVFT7w2Yq7VTjVj1TAug
+x5zTFsQ9QerjIWfkiPylivVk/VTSPuJhTdy+c3viXX1VDk8zm5W/qlpAChN7tY26AiimjBa7hhT
j8CYGLcY0wcCAsFsGrYd0U2Hp5voaihvkQf1O7wa+G+NuVyQTBszwnaz72pbRGYoHqN7xBTi9+2s
0fyveoLPmenbVDatkH+jexoCjBkx/FAah2SNpWwE2jU1Njk94ABaj0wGOcgP3yutx6Wc0oiPGtjA
lFag3mj+FCcoLKhEPzmmYH0n29aXwyZ55YYIVSLQH1qvd4V4eYAoaQtTy4mQiF/u49vRolr9/6SE
xT2e7wdp7D1Rhq5FbeKjXkGMBcLFD24zg4nrP2W5bA3k2DRtohEV/do3VpuvdLJttzCB60G2wz8k
hhe6ncO/ekDLA9OQbzmYTfMyspb8HIWtr87pKBwX58C3wgKpizGIle1TtcgU8kBChDS65Z6QBbmP
ayKIVV5mrDdninQInyra4t5Oqg111X8+WfpuY46AbdN5e0MDEengLlIrZv+3hw7hr5uTkVnmmkQk
opuOJ2HYmlYcrdMb6Q0Wlep3ZsnNZqeAwxHAV3Wp0KKGcU8oQADahkmG7r/und33DbtN+WE6tiZe
XE5vNGjb7XeSm8nEYz5YlUKWhKmJkcoftCjY9iLN423LmrtL6TwSkh+cM+RsFTuDIBvgAQgjitZ4
X/qMWb6S4n2Z3rECL1g3B7Knhjg+MYD/4OHJsmZRn9KjrNVpnYkZC5CuwNcgYXsIART2RXITJLXM
1GNBIPFveHK1yVnYUBsw6vIDIp+utUhDS33hFHw+DnQ0up24BtI+cPVXxICAG81FW0u6qrSaXmoq
5yI1G0dDbl2euH89SixiniX6bpNHYg1vlnaiXHxyj+99s77NrKD9psP6FD6FlAkKZATfJLN6sIxP
tuDjz+w7cRBL0zyVR5TZoGy+9V0iA1uQ8EMG48mdKomYxE1J7o9qo9jGFOoz3SUHhjoptna9OaIg
H/vU4u62RTPaO/QF8PruD5lyImUqTohdPuC22OEDqpmK9bIW95DjR160TIXWn1pejKjdmWetaOGR
HMjqw6h/PfP/U0dqGFG4pPW0v4wMmsc6QkrSDLFGTZf2kpnazPKrnJOHBuH2B31ub6Paoqy4Ls2h
Zy3KitiFaBjRdvz3sNkXSX/IlR2DvCXhzBhQnFoSRMTWU8ogeCeBB+FjOu4Fs89MeQTtcBCUOWfa
FLPFRZGgWbSIMhfvFg/pO5GSvQmPUkYwKW9zRVOOs7lLz9KlrDRraGV6SSplO+2ZlmbQOmt8Cuda
CfzXJfkl8WMB1AOsas5brRBPxvIU2gvr3TqzoO9bCq+6o9SZ2nE+BSSPf0e8KLJP+cediDUdFvQ/
Y5Ez/UmikCuLeOVZ1x7V+gQ37yHKVt7XSXZincg0CMcE0KLOgvDgPsnyTj9V/Rf9AXLdFBGHbFD2
cJ93DpD9jILv/BGMBhUGQlUjd0O7XUr4Mf5FCNTiMa9WBVYLxs33zAYK6XgkBd3PlZenOSM1bv8O
1n8teRN0Lee14FafrxPbi+H+HUnvVmqz8qiyJVtj4/VI9O85DiNH5VHiLAg/Kold1SQzekz9sg9k
PSQ0kGq8wlSvJqcFNBK0drPEoziFj7PLkiNMre+Edq6eXcjFkIPBO1YtAKrQSSZp2hAwJGVRN3rL
PzJsphXhnZ+mqq4wHIEQqGzanEtr2gXjJ1u1pbfd4fZCu9pSUhbQA211Ezn1q+/C7Zaw6IjUpLQi
6NXgsnhmzobn6MF1Ty7LbCKZJh83X0gkumwiJ25EuPegSuMFhfXycKCk3Fn/PErjq2WJbYoPgQdY
9SloOetr1ZZdJxcIdWDpNHKIrIXdpVEQHT2hrtyqbWAm7jNIgwbW8zrQgyEcURoNTeNxgca2/B0q
l5KNPux8GPYDEdqDyiAmc4T4VWQD0tLyi0sUbm7rOcFY7J0T6G0PQuFHGicPy5dIvRcrUj8MMEEc
+Ue3ZD8MCDHP4d2nZ1ANWI+OQ9YEZcjWttAx04lryFZBbkuQYkZEuyzeb+D5lQkJ1+IZACsfVvcO
OykbxTsf7mYu348vsjZC4U/R0nmmdr/HQgd4PiCj/KzfzQSRFtcT47Il8rZNBcpWKccc6qwAPhPt
JieGiQbic3L27nzwF8UZTGxY2+MI6SJiDZ1N0Pw6sRUf00bYx0zwxo3hGzspP/auND/VTxN9oZjf
Rz4w022PiwVlz6v8iueFiZeaPMrFBwEzhQlq78m119SYnGuOKSYeAlKuPQuHaigmSD3kv2blpl3w
bJ1bRea9GRXe+MfoRSFZQthaWgBEUliAZel97KWoDmO5xOMZxdyelRP3deyLKAJMvYf+8uWstBvN
ZNCPBdaz+pLqr9uud/+nXIXvDiQAAqZFd7CL8yI7RVouF7xh02F7PQ1RjsaQnxV42fHN3Z4W1BBZ
03B3TgW/0aIA0aMRwg7a/iDDgKLZsyzRE77O0RAR2t1pGvV0CZdtYRtKkB+0JNq5eoFxueHIYM5j
UfOb8f7aTP2ikqS0pUhFynfLMpHrlaBUORcg1P7Y411w+rfCZQMJ1m+anMqT75PXaYvv9Xajd0uH
qKuZUEhCcnIzsfL/X9Zld4900MIGbfynO9yCG0O2yASMcZy/GT/b6sb69IAUo+jFLb6rDEsqyTTL
1MXAOd6e6ClxlU9QSePxjzyC7ST3yHEsn8H+Kv9oC/s4kLf1UnB3pJCE5qpC0KHHxONG8keSk0hl
4dhM/YKlsVQEE0leaFwq3PoST9tqfvbYO8YMKEGXyiACUin7QMZh7pOwWHBC1G6J+Oipx6kIRE4a
iX3cTjAi3xf0FLcZP2OZfFNwW+OT4dhiKnZhlDBGhUy+urak2utb0b1QYo2CSPnghrhl4v1sGYy/
wAVKNa8rpqTqmqDs/2I1JX86aRyhwKdiAtFriWML+FxjpNp08MLPxaQx2rX0Utuhy5+uLQEi3l51
PM813lgPhLWgduFwN0dtFBXdvk50C8f5NKkjOc46yn9TBWCHFv9s81/RYah1qyvpZ5O8JUhLiZRR
64uD3aYkxcbhquA9zykBTgHAJgnxoefng0xTxha5FB4nt88wBxVlXC6ZQpWmIlX41+WZhnbKAIJw
gq7W/dhLLOYTxD32Z81l37Uie0llTZmzRZ3/Ro92TTtB9IStJ+Rqi/pCRLFXDeqhkR5kHtmsrnJU
q5RwX4BjYRi2qvD6PJRsWlZHe11g0wOyYpNW3da2ysbUKvlVhmqKOfz7+SAjwIprZiuQUHJBwl8D
apGBU4Q1WcaeuM7zKUDoiIfi42K0TVVWB1jDfSQWfyY3HDzpRw7we78+2vJo5l2EZ+0i/Qb81pRL
oHghlUMS/+DoO3I8HrHL0iXlKGhkUxTweAF1mQiBwbVqu+QZlZ5ztLqUv2LJmz5a+pnUZ++wYuEV
vL0XNno7zvgB7esvwxiwy68WRQO+9B8n6iYxW2m/ZkxvO6/gETqGJMj5CWghom81qOBqWZ0y/9X6
HCF/l0ZPKX1c9hdvu/IBzsWs/CAywlOBUXfvarOdRLG5H7T0XQ49WUKvauQMAezMCUz4vIH4tCrL
75hm+C18WvHRXIPAdDW5/yICTdbhoTAOFRuKgFnGlwTlOwUGk3UoiS3XO69bOXE7fdgRBc4hPS1m
n8W2eohGcWhwITBClqmaD+luxRYE59H4NwJTne4Y+9YPqROV1O6uLgx2rhTzirudCSLx3ntEkiz0
98MUjnktlq0J1CUAZhLcsjx3WcUyTkHVWqcLkfu2QWAr2HoJ+lPk13hpq+r1j8fn4NaLnzHlkMGb
63KHwf+AmkmVRU1O23KHFX3kuqFhvexrSq9Bp5vIM3ZpeF8NyIuc2cBu5tinl3uRVmC3A+H3CL3A
WxLN/RV/dqeP7cq8Br7f04wpAZUQbqVovF53GAPZVOBRlCyF5JC/6rTColi9CbI6FOjuMbj9Gk4i
FmbmInZITARDFutfcXHuloM+2uoJFTAiYQ31sV7BPGuu6qus1pjvLdL+A+XrIzOYaM7Q541xWUax
UD6ljPNMcCqE5qkkCBsWtx6LErLZBdxlHlcgCGRjg37dJAKz1PmKEoDZ14BzKueJictbSm/p9H+/
PCDhdolcefZS0Zx0j2VXdB5632RoutKzWtrc29rkI1jN9b5vD3gN2HqZdE86OYRNSQDb3Vm8JJOv
X3jZa8Hvr0+Zkh5KWlyqt31o9i7ioc7Xi4R6LZS215XR/QKZ8varHGasRCk6+d/9I4Kf4cpe9P0X
NevXDHX+3TpfAfhaEAwMt7uwS+uZfzanTTK+CAN3DowcPRS6KAJV2Le1EBqmLa56tCgoHi2As07a
IRHmXqpLAvz7ULc8ZuEvqCtzgJN+ymgBmpMHbzrrUwXqGHufKBZyE2vF1qMS2NgdruXXbFIV31lx
Zu93sTOuX4otfEMCqt/GPfKbEGJW/Psgwonkqg11hVLok9RqYUQfCCHlFFb9W/t6LL+hmz0Dnhbu
HWR0BjWqprHlM+0CFHXRBLzBxU53DMU7u5mhQ5d1mBHivTPqrc0R5H8gmYwb4Gza+ChHfmwiHvcQ
N9hkeH6XNUsAu5UOeVxu7wzWRe++F+UkpqUpZbOWe84x64gXywoGy/b27/IL0DhEVKhb0O0pL+kH
/w7vqTyG/kG8lPuwep944dippTkJR28PkvsF69o224IeifdrctkX1XjlQuqzpjmOUXlsX2pOfNKa
+rR/b4RlqXz8BFD4a4mfJLw2ASIxoW0ykt4pajWYFuUkPh2wlvlGtAGXMQs4miEfH1I19j7KPlsF
PBIVlTCLfGmBlV4Lf+VxjWwi44Y/b5xM1DxieKQ1zK9ay0i0lXfiFwfGP1HVcf9yI/n9adSxgoXZ
3NCHFgfuLuWZTWFrtm/TfmkRW5tXr8a1ms7r0dQX6IL7hwlLbJ2aVHneTtkcEgW2cmkuNMy/q0kO
Zkdduf2krndURCKohn36+V9HkkQhwG+9rVtxgO7ApHKornnleQHrxsxXYyYgVIvzNeEW9I0YYiPP
c9x2DXatCpX7+obe/TSds65IBLEM+9w0VC0R6Ts9JV5d2tKL/2ds1gjIJOVFM1XPg0OQbVYorHKk
jngUzDm+I+q2d9rktLzARNd0q49qMYdpHLeXZu5eXrT9tY0yrZ9FoI3YwgVGEx9EZwPwcjsY53WA
zb3lrzS2dj5IOmdP/nyl5dGWIfznMreVSMVUZuVpFUHtHM3aSwc7FVBg8vW8w+Yq8DZO5uxf1ypH
R3LKdFcFPhMOUNVrp5rIACU34ykUItyfyDaB4NG0c59v9Ov6bWs8zXrxQIAAM5a9uqcf9838iS2m
wDAqnc9iJ6WbhbeJmfOdIF82ivIGoc859qdGS7tbPByN3SeyOI5N/pw2dm5LPAo2QUz7/8c+Tpci
BRM8Kt3Noj88zeVRBlSzpOizymXJYhHutwWBHMRdvuRC2QXKI/BgbjV8ueS+eB3cOGqyku9/Weka
RIBMLTKb2SsjBoylQbAdbZLjXy+RNqGxkcLdhMQhlf3GmHC6X5gVjT6zgyDnJfIl5+QudaQN7sGN
anCyJ5CdoGBjTcx3NRnpFdqcU68ooB7haYW9/jfMBnyu7r53o/13fipI9Mp85/m2kL2wX7H/d8kb
vqM4UyPM0X4yoFfk1DzzGBY99CsVhli2mr3ODZyyiZbqKhf18VyWAwrIDhLChDSpP0CPqgdSWf1D
or9nRoR45S2VIkSw1OG+NqGEV2XLQ0ZZvBNOKr/C0RZzqIYCdSiYxaRD0WLtml+vd+nEkntcnkJS
BlCGZH8uhQq0H+ti+L6p2SVfGPounA5qwBeOQtZQu9VwxyXCsxmc/E4azRc7sf4mcQmZXISEtTXM
U4KlEdqqujV58im/O/yhZL0zHJeUtjML6NtbsFb88kk4wXeBj47Cy2Ip/zEf2n1sVJESfrI8cK3n
fzX9J4vLrvWhAScwlunxucgBycSf7WFjSqmA4wjs0QCB5HHmWybNygFUqHM81PfWVXTsTGDydcT2
NW4+BwmEOa2TGtj7TXyscaesa768+mxvKgYiau+RpRE7IsSNVeXcD3C+utRIxtw/vf+YlE2OUbgM
PbXTA/WJHykogNwypmNyTiEbZmvqjI48NupSkpP1aYqtJzYkQ9G5wfT+7URcfvyuM0PP6ayQYkSz
yqUn3/uRr/Fqz0DJC/pwPt60HyKiKkblNnvU6oIFlRe0iAqxKUmol/turWmPV8zBrPYGN0QiN1am
fSYe82g+xxS7HRS/LI094/1Wz/DeRbfYuPHayCsr4jH15w9E4Got1mF7Bk6oxgfKjQfV9rZzy6+r
nttZGQIgQo/G1mE3WUGm1YuTXh4wyVR1F7aUAo3vbJlV6VntJFIN0wl9sJF1pogpQYlgpkylUhZf
wAjNogM0EsIlm3Mvv3P27ALSDyZz3JPi1dBjsfHLw1JePfiaSeiLY0UGBbJkOtnIYokzUj7/jmBX
eZxaEsjhkIqW/Pb5tt2nGaw0854L+exVuXT/WdpYXkuEa/tUls6iWn6rdJgU3hIgJaaGRYDJrWtl
5hSmk7KYohOjzBdpS2ZL5jlIDfZ1fnbvIb64bT2Nm/O3+23i5e+D6s1BC4zHfVfnthgPtJ+CZT9y
sd0aDaFboTEoBAobKwMVsPbYZ2fpKb0yR1xyvCpA7qnQchn9bnVlvGK0WzX8s4sF1hWrYKaznk1G
rjehP4zQUxdDW+iLCrJYrBnzAaXfZUuYyA/b538vI8RlswKTxTy9bgecPLZz79K32LebJPIJwBa/
+/gyfXj0LCKB9hmerye4Ywy0hRGf3JbRfURobQTm3yDf0Aj5XwQHu1JaJjGA8AWbNSUQo4MDG9CE
1QwZYpIByL+h8wlpLbkYAGzYt9Ju0PLLt6ijCHwSpXQDSnjGG4T6mjqd6AgvrXTetSM4TkAMvxK9
rYaywlRRYRz7yblFct4VBs9IIpY2H3yLEkjLvwuPj1dRb/55uJVpoDkmbsf4nzo9FU9nDcwLRoJd
0+7HxlxAy08F8iUt3G+3HmqqP0imgOiYgq8DMDSKM1WZJIY/wzgZNpGDVABW5U2ATvWfK5DCrblW
fe+DzPnliyYGoehM0U8cp5gvkjI6wqLX/3dXDvGcHJ9PuMjan4SbeiLOT0qgVPrv9NKvVlBD1wHY
5Ek3Bnfgy7QJifLz8PWn/DFfkxI50+hxvr3hdB/e14aZKkmNiVlSoJ/ACcvfH1bQgmsZdkXgGW3e
4Qo65sr22lMzkhFZInSMe1QgAvMc6ULc2R9hD17JBg7bdX6kRDV6qwKhP+FPy15ytlBweAi6hVFe
E+NrLjOctZx+T8zc+J5yW0Mej28o/v6njT0FGFaLrdY1xJNRn1CMpHh0pZdBzOa2JVSsT/cMTJqm
ek1wVLok99gkwFgVThF2xG+jnvXVwY3sIq71Hu25iZvzK2U1Gd/TAjC9Yo9rT3G76jJPUC3Wfjve
2qvkry2Jasx11oWYgHDuuowG4U14jukzliJ3bJwd4e9hGEB1BDZ4lwfoAEHKpUhTHA3qhKBJTITd
7ENKiMGQCA1FXU8ah4zyFK0NB21LlEedYO18kSAJ6eMAsOumhfqmoQ3OT93WR/2t3O6KhfNycEYA
tMjfm4gcuXCa5ewDS+X3am0Zfam37qYLpQH+5I44CAW5xy4bmkRdQrus2gsJ5oV1l86X6MKZwUIh
rcL1TnDcXKmFbiJXODNSfU41KvQWg8B3QOX2EWqzv9wKOm/0qg3GsfjNFRAMF2npoBfG9pdPciDf
NN+U1hH26mVx1/ct26ugGFJgBct/9WwJ7gH7gpd4bw7htnnzeL01Zhi+Hjq5ejlPJnZKYFRA6yfh
1Pxt8J1JB98cCp1+n6ytALsw7P7yNQG5FyI8TuIJpbJYPaB8UgZQG6yH/WmNEMvpXHv0SCO3YsfF
+JiFomrQQPxZxdjUfemwKjp4jZ1eRE11Mqb9ObN8zC3IfcFj6rG7uyz7/N277OAh2aU0kblt5WBU
VydtSADMmrl3MBHLbRw16BW775Rn7oxBe9wz95b8QJlCmJgKg49xqdigVMnb7XmVOqtLT5jB3nTO
iNOaA2sgjL/50DytwAOmcffaoFeWgCuoIH1XOjZt3xsncVAgsQNTUFkScRWDP7QNsv5xMvFrP/o2
ZMvdSDlTZEuJXx1v+385KI/MjBKLN2L43vc1V3MWOoB/2W7Z0TiGhNc+wCODCUlSNlU5m1f3P0Pu
XQrThnRujQlDu3hPnUBqa8XuR9Ead6e01Fe9qwMja7g/5Sp98idKHj5f7Au1qVnTNC+nmLqVm9wQ
RUSYM3vZMgpnz0BE5BFBTEzlp8+dm2od1JRq0HHIhFHkyjgVPwY0q/RCuhz/+3iBk9fD3PVcY84l
j07A94Q49j7Xba7VapoK2vNVPv8940lb0/tCr1RbTe3mWTcjLFOhDjF/81xdm0cVDrVUmwwvfIZR
UyM4M6BH0fU1QSaD12oiPQxoomVSDUq6zJTqTQzKZ0WnLS/pFbMnJdRPD5xT7GSayDhWGTh/UHVD
JFtw1MHnn8ElZENOzXWCF+bQn0V5hhKAmcL5DBcPFy91+iF3kW+3OcNZc+rxdmR0SitdwUmd7Hs6
Be3kekl2DvKLOBvlX6lWe/polBp+G2zvnOMRVO1pn5HAhwaQc3BUBQyHseD47GG8P3CqNcVKwCF8
5xSnEOkAGas85beYFwkMAnmz1A3iPmXkCI5ryMN+nzMP5zjwF9Uhw3pvLZaIVuzAmIQRWEVU4QX+
Dq07cs9aI5SSibUVHYnBQ9Pa+oFbj0h0dLUVBnbR++TNigDHjyav6GfX0syYwek0Sfi78IxT3j6q
Ljp7+w4pWkIW9ZYQxCw22OYB6lGgnHbk9XeUH5GbG/zyI0bp2F6HUHgkD+Ii8I62KNlGYG4l1fNP
1UmAWGxONQqfYmmJEOALn6mZrzSj+roZrDfbhqkF+68amJXXIer/RCIxS4zBic1oZX6fMinA+U1D
1533BKf+fxnNoEaEXXRpYxYunlWnKXZXPXK1AL3RfAnnBGUPEtpsPgX7sF/f6pcroq/vZUbPdRip
SKZJAB9oPU4B1ayUPXVGJMx7Wj38aMNbwhL9S1NvViIh8RYU+aPYwbXkhKZOFoBI/9RTNCs3vF5L
EDFttmb36EmQ+ORWhadkxEOiSQV6pn2aWDe2XVC6LSEhfiRD8K4e5KEFERxzr/mkW49ripCooEsh
JIQgOfRCnkjwD7xU5HyDPd7IlUg6HZcMOAoJy5DBP+CgIqv017ejep6noMZQAjidy9X4AwbsNDuE
YRhHK2zY2YpBJqio4vjgPwz4f41vlBaWE1AeRnHiOpKtxIqpCcwCsIh8GjE3LvNVvEyqenBBRyuO
pZdwDEEK6mYbghJzoG4apV/U0kS8FSmOgxKBskMGxBXYSJe+NZ9sPREPsF5K901njVFPqjn2MHFl
sZ/n6xSSnBFtjepwrmxdf5HEQu57UaTZ8joe2771T38WGaXuFwQu0aZpE5kY+rrkUJ1X/s8lthvT
AJvAVpOrgq9WE1fmLNSCUzMgbcpqSdwYCgPaByyUD+E27VQChDqD6rKS/ndBkbgv2SmAtGCo7Mpa
kbZ70L/AymvsDDXJl3pqgNuHlENMY1iPer8+cHerwSvf3QoxZYiGRjD07yDmRzJ9yphV7HlrE5aV
juLzoBdEefJqBRyxQ+wYErJAqGTlFR/KWC/VLlsozfNs58TFrRwiDEKr3oC77lCKjwwpMW3CTzuy
LUX7fQqps7iXWXb9XEnudzmH1oqnGZIgwwmL9tV41PQwZQdhrAcZVD0g1oO0E/MyAVWPhK132a3H
Q5t0KXD2AtKnDEx7o8rntNB3nUDtPRe5RjCOB9WYx5E9V1qLtoYNmJ3b9THULPqJye98Og2BMDVH
+XZ+Bgd+kmMysRLgrJwsOYhUEFYUldCQDBpF6gUOyFzm138Iuuljz43hgVzYc/QYWS1iqKZksby0
rsSJpAlml9PoPrlAzzxMhv9V1paVjqZFvmjqq8YLKVYVO7kq0ey1DWZbDtNinfcW0WUZDsVm8Oub
jzZ5z1koFxB2NSn5/cov0cviqiYc+RpuDBvo4KEfNiWmEs86cqLwwn57Pi58vN91+4k5ur56io3V
9b6t1PetA8VylWYxgBCLmWNarBJ//Hlur6+wHYeV63g3CK18Q52NoL8bxK4Tp1FwfcKtJfT27Dpy
EIFxNmwfKKu0TTnqFAcgmBVBoGUrZ2TS4EYgNF4chrN1GZfEzueYvIaZo6AUozOddOeZMe8EDwqL
ZXfThNt8Noon3FzNNsx4nayKQqb499RpTfwmVdHt9fc6DPEj5wBLH8rtFPhnCh/SlT2B5Ww0yqaa
65FbprxVjd/v2goMWsIAGS0bZPtIGPSjfadE8zrCf28MsIcWhvGoC+lUYdxw2SSH8Qj9nWdcGPyU
BT9SrUEzjRg3YTSFHgEFT57HpkCgmmDoj7aP8bQfUQ1RK2moJy1KXccfzXsXAhqu2+0A61Dq7kP+
SUV8URm6zfHa8Umsssf94X2uH2nzonimft9VbeXWqlFY/25WIat4mRIgeC/bN1lvplTi0nsqfI7y
iTuBX1ZhJHyJbsjIiUqA0o/p7DCNPVO9ztW1G3bYd5LpBOmdLWzNebz5a0ROyyBux5xie+rUztFd
MuvtEerynvYMgRoFsBwUvJfBLoEiVJT2BGBMu6APONGo15Q51Tt70IAWS9TzHc/O9oTvZG6hM/xV
3Hhi8kWOPcCJZO0YYPrxaiQHNayqciMnlPBdLYy+cTxQeDNm1f+pCm6F9V9Np/HR+RJ+c28CBtyD
BMZ5KsEsHb3Eiy4h9npTXeNXrp7bV3bnV2E9xnMj5b26/Z0ipzYqYtliBQF1RXIDkE8T/jtR/vYM
WBi4ZwP/rbmPb4bRusX1yWZQEhhJ00UZlXPj7E+6M43yeH8wKY2F8TfGRP2D8f2Vo1s4WELOE8gf
T4Qud7J2QYrnXHlD7qHWpmvUT++adAy7/1/KrG8nUPb581GXhK9pZZzuDP7ZphePi/okuAPb3+S6
uG5zXSqu/t6I7qK3cEdaQAipHdjhmMfLurz8zkIBYGNl0HRkzcwuhK755Z17PmzOIX9lQyWYBLfR
jOumOXUKDWNpe88Wjb3AjSlnTaWlHKrb1tT/SABPLcPIK6TpWYEpkfGHDNgB2DsicTytHtuHNZa0
a2gmTKxtDvmI2g38BjMvuhu/NqAQNbqJYpm/or/auBPIVlQWA9w7r/Ittz3NknQvmdY60AAcSO/6
aOYIu8/otcWK6iuIPUo/gG2cCXGNPM+oTh8vZDD6imDeY1pprmVaGCvBIpwOFXGK52h3WlHYpu9t
2vfNc3OkgQoCEgU2Nzdk8wxFbKSYYF+mAirE0jePQE9J8Scxgp0MR647zv/V/SQQwCdx60WRXH0x
QopdL8jMzOnUSc/BWzSJyXg1CKaIFxmNdpuZVdd3AfASpzOMs1uctVeOwPlDlLI8qhx5UBDM4cvb
9ixHJNPvmWluec3j0LL336TTHSdnZ8DFs2XFngybCG4ApytbSjV5S7mWgO4TJcYsbdlITGw8YzVR
x5AAOHx/ohqOVDvwaox4ylBR9hlRzNCc6SHGvDCuKQuii9uCURV4S+FsDPuVyISrfNcKrxlviJbx
Sx8w935+4rvXvfCkMeH9UP9VtZ0B2X57G4zHncVijTKWUhv1j3Ai2As6OgID7qBWqRHkCANjA7Jn
T4kpGiIzqQsEgeQbj1USN16QC61b4/LCPhypJVAS/WmRoPYm39NB9UPLostHB++3lkf9j52B8d58
GZmWu5UNRsfoLLGS4VtucWi3bQK3x2my9zP1GSdJpfEKsAEQANpFsmdkof3Mb4tgKUfcxJJmTDos
yH9Rhv4Gpg0tSWGb5cszlEJJBYugqdDul7/t8EBPg9JepOKJMDG61axkph/cvchWSER1drFX6iFa
N6f8ISvIgYhJQqdSfS1bf63DJF4ORyq/Ztd6HmsbJzQV6M8RLy1kQ4FO7lB+qkSvPimkyqm1pATL
wOekuIAu4M+QioTerRzVjCBTwwYOCD7o5mwGcKBmSp3Il4VoQeGSIP6slmWzabulRbwePks7cyH3
Th05tvka/aqeEMAzdMk2RFudj3DMD35/w0SvkUXooHCAGoHXV9+r14xad4R6tQbprnIZpgGF7Pux
v/3+S7asoErTPTZ6AKw4UpGkk7vwjQgZPu+f8JWpOMf7bSPEzKvXNddR4gqYDXmSFgD7eUEmPSH5
Nw1XTsMWvTIRLc5Q3pJq3J+IK1KZojg+L5Lm5NwebL/SIQ6z3WF3y1jvYLMhfRzHA5fPloA7LcgX
DT9zWH3Q99RkYSwoYB3AzwqdY7bQvVBc9ea8X2DVYsdydRj16W4HnAH7EdCy+KL6PV5urYoQYAs4
qonb1Vx6fTlYf0e1wrlNqxGIPggekcYb4qLZ9y83joF4M7u8a34CoZDawkxwSpzl8+vMOT7Rb6h/
IUPlh/qRDul3FE9d4VF6hdz2V7pV8BGykpFAOpCfAZ9fh7PH6HLKhr8HKFz22RzCZos1ARqMZF00
gmReQw6knbCtyfZ7HqlpY6eB4Rbs6/+CWri3uKpu66qwoELssHnqjv6iljs+xfTtBMjKnWN4YNdo
Ep+zuQGP+YPgHEn3GHFJNWjxfd1n+fAPHX2tXwunBMKcuaqCQ6KYWYVr29r6HjMBp78ySdkVmbRe
tag+YeeciYlTb7/bg+66g4bgvQCg0ZIDgMtPMxGBuoeeyDS+Hw4CmfXhcPBjzoH/6cUDf2iZjLW9
AkgbfUq9nESXjhJPQAVzJ1WoSPaV7SN6gwzCsDX39ZZbg4RHSTKNpBrM6iiFX80fH39O3aplQJM/
d04v28VmveOkGvcB3MSKhY96eTix/LekQ+pwLNEPIlwAKjkmAN8f1ccua/QZu56pDMo9mD9Zo2+o
3WCT7Ns2fo2LyY6KPe9Z5W8xS8gaf1ZNdsKMs6FlzQpeJ1gL/P6yDM90NtD8yxnfZSzs5bLuV6+l
fzV4QQfBVjZxjVcjEGNrFYhbW/dHuX8HwSflcZubR+bwlwfsoJiY4GtFlE4cyr4i6vfZLAGrzvuM
78BJ4BLERevsP/jU90P+cVgY+Rj0WAHPTkF4g6r98DNa9z/NDyjg//yDy4ippTcSvp7yTLnQfdkN
mrjV+Wn01T97rXsqDAo07yoeLxJIy9gnqV9nvgnfVAP0xfOT0Jf7z7fF9qYj7gw9q2i98/LbJeKV
FGP86wF7IWJDbCrqGsL1FeZ6R8kvqwAsxrwaZWtoXe/uptOR3O+leOBUQ7jd5+vcOLaFhkvhE+FZ
U7uc6U+0/Q09Fa0/9qmojcU53UiQ1U8HWkKDXTV4Ri9s+2WiyRtjFpTXUhVppfs4hxv9ayeUJcHx
nIJlK+zDe0Co55s73nNYZXmt9GcfVjQvS08sQMOTVmw5qpFgiuX80DMJn8PvLAPP6MDO0HNV8FmA
HpsEET7GBPRIOeUKDwTfpHaKrSSoLA/gkf0pZwyC8u8Ao4TySOfPsn3n4uynWp3UkYtiWPJWy+lB
Yqab+JXU881RrUNN655aKkNjpPOXhPTj1ZRBXdOYFV/ozfnCD8YYhefPGagyX/ZKLvN7TL/eQlkE
zeAbk02dzpOe9KUVh8MqxuCpfKO1R8xekSrChr/bbAS3ZuwIRd7XHLESXwSyobZDoib2Rp7w5ve1
gXp8SkGYxrbCYi3VPQvItZqWsNDgtU4hKacFZtg3aAAqs1LW9E5Vx2HK+DJkWQeW1LW1LWAY+Jtc
neDqY1hhgb9y8ibRh8SDzvE6ZnHNhX1H9hikPR28h360LklwXTJiQ7vfQ9SVgubbA4qJkb27gPss
3cgEm72AgcVCUYHr5TM597FUGhlO0xIanv7G1AO2KgaK3uWCVKlMpajtyVJFouv9jP5LMjl2+yai
ffTxNXt6foYkkLFfAM3NFeVMxV+rvoigKS4Fb08mHq12aPMC/7FhfqyxyvNkvWDh2gdrHLlbZ2DC
TBH6StvQTNFnMyF1QAd3Y8jFz7bcxsuzY9BwmSb41DhdmbHmNqC5yNoA0elsdwJFjGme6lUwae2D
wd9a4k8kTe6VGncJ/K61+g7Eij8XXyS1/6u4zCISy6DChbDnCE3de27TbDVwhKUes4zQo4C2p01n
KC0a6KzKcHNk4q3tgJl0NKu+Z25xfc4JcYSUyx5hT3ZE5PgX2DLGpmfOIPwgE3rToKL1cU/iuDLL
uGoyvVHJapZJcpdkpfd3B2eu5we+KU85e8EAEDhgUu3p8N4rI6+EdWhpp2xG4+h+xVph+RbO0msE
d0lcFmblbSmzSHic3yuvRxfzGJL1ZziOUR4HDLLGtZmU0YZAScAfL5LoBhrzAjf4BiUYFcyWfHcb
jX9WBL47CN26qIZaNfT+Pi62Y7wVZS7i97M4rJVCR/2v//SDVw+OZlFvCvkc/igSgvgb+QmS4o3i
DSSReFjalu39ngsX9e994Afxs0BWzRjhqpuqW2fEI6UN2yd5dfGuxepJtmw3qWLhXB6J/6ZqiTdg
dpRTcDuBDMIlgOtv5UQwOuKn21VXCJvKtenhKn40lHFyvx0cQcfgpOU1OjB0dyEqo63ApFkwgXBt
Va87mvUJCrParQveUAM+s8iVSwWeibJ+2DEB+i34qgg0s7afWpNh0YKPdQbGZzMCIJJsGzMyJ6d7
Ua31aKmdKNsg570RgwQ3LqIUuCX3Nm5zl+O4RgkQYsVxt26ThBF5Xt29js6aLNvV+kkqZLy9PK1f
7QZotZ/BVrdihBveo37xYm8nuUIusYmidyt9mk946UTS8w+FhiJSv7JVetpK0lLBCWTks4ZqQhEM
b4TJdDT/Bx3dLdCHVOxUQkLp3AzfkCjuOm/nGvIs6RZwzgtnhc5bK5Q79Dg6nT2efufYuCrPuivf
LcyX/CNhY6MwVJWsPN//VqF/xgvQDEI2ZRiA1oxS+whv1ibwBJBaow6v90UjFlJ74gUa3L5GT/OU
uQwB81mNaYEyupAXq6goRnP5ck3KPnctzzc+cEGYyik3igrwbATAmcAt/ncHcbQnLLTa+33mklvN
ubxREQhFO1ryPJwuGaW50/9flV/HEu4ScH49s+u+5ePAqo5pzLgpnNo7NyGaQJsT6QW0ZMI/IFp+
LUocb3zTTKK16ySQaxSdHdo+KZ4XOumOOyA5MsGI7gj4eIA91Ljrf/UXgSlgTcB9zB1vDQLeOnUn
XWW2yOXo72OVfZg+OgTcKinkl5YXxmN3G//l68gvJka9raSPmZ0nUw8k5gXUfJh4+V6OUtDZt5kC
NOk1C6J9YIKVIY8cDOjOo7/MB2PYyJggfNIm4lJz+aX2oyy0YQVAOy7PyYf05PbOfvCoKWecpo+X
CTzshqOJCLrvRjqB0ktf0fWyvKxp2Y/e5dEnYLVPEBeYlIC8D1YmWNxtAoxHnXF3zEif2JgE4DJz
xnrofiO8z1cMcoFi37kcHxx4nb0am02PPjVwlkRyn0k25bZ43gDkC8kjbDmrTJyQIdSi6qOlnBsX
4dNZ/u2uyT/UdWY/X3btyEzrCoTUY2hnHg7OmzPtuvK5T09MWzwaFJwksZGkwpdLOAc50ZsdKFUe
06jUCRNfP35T5tdqsfUDdA60bG335k0AZ6b/BYLGTarzLZPvHHkuORfhjU2weThp5agbC2S1B3oN
gRCg2t4H0aw2bDOXv0EGHv+LV9qlQZ5ICyBVxcfQXeauAPbP8opDpIhGh8QVsEsAd3Lsu8AhQPKU
XcunSHqAWQtec12HW5PsB9ohT/Sjp9ToAXxIipBC7gJvU6B4JWfuXTaBHtsXJmc6Vd0ZCFCuipo4
KwBUHQ8Zoh2MXlfRvh0jLGw0YyP9d75HLCpFMXFZ5qNqUVlGBNBEVBjcYJbbxfKf6D5bIrkYIdZZ
vFIuXwNSxLOi6B1DHI4jUz+pRtazmjUazR3s2FNPUGaKFpOfU9TArxKDvi+XGTZ22w7rtCi7BGG+
1yfwa03BXRyzfdmtXH7+nYJPh++quvPwSqdzrE0Xzad/2IfI2nVHnFuyXLr/2uzvPjfOdWCNgYXf
o3VyPOGTh6pph4oWQTt2QLYBOOPmJCx44FpMMyxNuBvRRKBpPHtWmoy0Vwc/5oJKjRkdxRUMk6WH
7xukF5NrHk8zX69hBW+C2XLU2s+pBJ0fYaUzUvNwr9+wJiAF7Ami+HqDp+H4rgwPai+1IKf+QKHI
ib/Xq4vtd5DhyGS4hpnssarfO8ZKz+Cb/fBTGQvE0I9yKOAdxKrrvfaoVoJ176pS54MuP7/ZLR/R
xVVdjJh9AXJTMa+0DQIKFzE6e6Dgt0DZFVqLjEbmuInVrAgx6oQUzUV4Gm0Bz/Q/nR5DHBgZ9i+d
mi6MuxkVNiA2cG59fHvLaiLf2JSIyddGifCJXlfukbhYDoYvM3gE1XEQbOY/aM7EuUD0WGx8N6aZ
V6ARV+jk4/9LdU6nCSLkw7Wtlcml5K3JwvDXVPdtTRKUi9vO2Vb6KEGFdtZD9hZz+ne5tZiSpdh/
rE9CqYq9xoJLOSRg+5vo250NlLm6WxDPQGcISmZcmlPBv38rrGemINMqhr4jhRco+CZ0KCgizFhw
RMZRB3fJeF1i4njgdhNDiioWRjv1u7sPlph5MA2f9JLdQplI5974kH33XFHI7ht/I5734zBO+e6/
5c5456jXfpnAC8tvRvVoxGRj0CXCR0w2MG6hgFFJ/sxboNAo22aAGgduf4d46YhnW4K0uGODCg9U
x7GIZtTvs7+75haLgQuM5484Zu0u9/zZWe8OodmA1TRWPHycwPtO70wUwbp5cPuYtYaF+C7Wt78B
9VEa4rH+2r5Lo1gflsELQ9F48g2gcNsGg4U009S8f9cKm7O8j7wFjxxlbGn19RiLQQD3v/iPXrA1
vipd//CwN4JiuF8mJ5InBGcGUzmg31w0Ei9/QzY6mtPTo1stRzAzgy3tNGhLuRBvlDXKp4hYa9WQ
8Lw8cX8CFoCfv3ZZhxIiTb0s1dP5BccZVl1h7ub6kcQ3KkVSKwa7CQNSAD8h8e5x1JDyg/NQcKF3
GTQlqLyrIOt6tJmkBEtop4BtYPZ1RwxGqvIxULUWfq2jAMzzqyQkZpirxr6C0TCsHy+N1S0PM23X
m5BnZwXAbnos5l2KgscjtITsUheYeKgZaPmryJnOLCp5P+vUL10WTu4VUBHxAdzS8VJJUoJh6DnN
Ja7wuDEEIuYj/Ruw/9ln8srey3i3a7yuMxgksyqKg5SN72mmrf04+WDH3emwUkJ8AuCqHJ24Q6Gv
9TH7aCKbfapB8qbKfj/xj06vSBWmJB5etq20gHi2Xrwy0OcFs6bEYVphXDJJcrdwng52T2VXiBVM
uulQ1ETJ5Jta9831DtUgMVTm6SUAfhpJmDfMbofdauOJjmv7iQ5tfob3RPIa2iV0LMumSIO9dBNJ
AzI6HHu0I6g1Fvd20QfZEiUDwnnzV244k66M47HE9LXSTv3T+jQrDhHYfiWrOWqiXYbVTkCiV2il
sFIdJt5LCI8vunw652ku2NXBkgwJ9c9qTIBEk5wkTbHZeJmZQXPxFdzASJYHu17hjAe/M4LP/GLh
589UvzH3V9p3+I+waHGiNV8R9M4rKTYECeowC56Zg/WXX+FbjF0vRDwAdOacLDvG/VVd0jew6+5s
Oiyp5DSRBsMecu4aFyeZa2ppJbtxx7dF6Kthlo5sW+X2EC4DvXp4YWDWCjE0E//VSvPI6m0UB3C8
ZxfEmetO36OA9U4gaI+qkF4BEkc8/hywD78w5Qd6osY/cLxrGS/1TZbNp65bBJWffbN8TjzCzCxI
Bq3TIlTG2HL72WTFqLGdtitAQu40XC48SQB9fpAcw7eOcnmGz+1zawZTK56RkEvBI2UDuedjfGPL
ly69NKDD+KF0jENl4uOYT1v74oYJW6/6HZZrJrh21D/aCOWVpe4k4LEsyWY8HzkiIxi9LrvMz5nf
iKn0qheRLXEoDkndeQHk5f/pGB/istKA3f8eAl2bKQipFd5G9mYLMz+ZgORpqYJx5sKy7Ey9yzjc
Ei/hUZhKJTx90GCfpxma278lb2YE3oHx/q2P896vXjo1AT87ZhKYCeKVwmtdIUswbkQWFjmuIINv
KU5lijMxpANgwN4o64FsapnVtQrGDTUYr2KxxsXwTppoQ8mIlS4OhK/q0mFjVi8D9gOwh4rvowHL
qiIH9NE5fJqOTEViJGF5tY6gql0yz6BykgdUH7jifR286BUQt0wgYFR5DegPZsf05pKPJ/tEEJ8l
653zEceWUbM3rgzH6B0o/qAx2wZhtDgFwU+yro005FAq0pOhWF+migj3s3y6K6PPtdquHAB4OQ5Y
F/Onk6RUXoDtfdPl7T5OTS+VNtkqfcw1G7AXoPL0+WVnPslvJEZ1ss8iUsQvtfvCFLcGvJQSwTKs
8OsahOwfaecBY8gl9uNvc2XkhUhkLwkYOtxNR34FWBkL7XkYDwOZnB1hPek3OZXuJP7CEn2vc1ng
Hnu+mfDz9XImokPy4QfFo9iGesmycPHQ+KknPbWqVVsdghmIz/MWOMzUR+5sUuuneZ4fZPKE4vsy
j/e4wwGCTwMntHF9Tko/wvqiIkA+fKm9To+cQvaW7Hq3xPbbDCwODnFIm54i3BI+rCeRy3YLNi3g
5VjGYmX4EnwkTQ5ItQMdCgYxFp4CtbWobx1aKNUhXQCbgSR9JVxAFH/JRdCk/RSGEllckWdMvffV
xGxlT/aJUylvofbBbw/K/uuvdLyIjTl0ntdGh/of2ME0sWlHWFr3tmnszI7j58yiDIJU7/bmbUIx
2kXWKz3dkvA82lbj15jKhLsgMmg7Th+04oCAqI263W2fuxBNHKP52EaBFQYV7xQnTPB0sNIM1qSb
LsBf5L+TYNTBRGp/PT8bmqsBZotQXJgfYqdpU02SBBa+jDCs3VFsmmSH4blzx61P11yyZGT9IA3b
AXoo5IgWKQ+OXd8byZuQ2GyAM0O5QtFcdUO2medZeF2+XeKrMusQL0kSk202J14eh2MZOEeF8ycA
UYXGV1uJ2VU8QqcZhFEwMQdODQ0N2fJqJHkkVdbhlBewnxZ1eGx19KW95RelgIZej6BlUhEoXzeV
ybqX1spx/2M24EU6/MvJwozrjD+t4BJo/qnm6vI3sKpqfQOyfkVyqeMyh4LWWfL1f2h1gkDKhrBU
/62fohfm8FNUchRIgV793PMeA3ar70eDoiq37bKwnbwxIoKD5c4Qo+1FaxH3DERTrDN2jySdhPDD
eyfstJ4VoG13EOVnD3yBXQ4UYEojq1j3GW2mH//9V+MllmAcG58Knvoy5DEwBRW4q93pcjME5NZO
+hPXI3H6oIi7kUmd569SkV2ga7d8TgzJ/KsvD93KGB6fVwu0k8HqfP6VQI1WzXbWpZ1Wd2es550Q
PZi+pLHt3+wt0kGdHAeV1lUuTvhsdntfwRpSdlU/grK/5w5y/Z+DuId0ifKoAM6rqyjHsHurDfgI
aumewFWeVkkPtHPg+AV1FD5yHG3e8pm5EmgA+JptUKQB+fj8oVBiyPNxnZdpFHT1Z2eQs5G6w6pB
a2TlVvPLBMbI05IBi1rejCKban/gbE1jBviI+4acH4AJclHiuDdlAPNwff5l/cQEU2Vj+lEoa45U
QiGz+l/mKjl2VNA4b66oL6MT1MUq+0Be7S6UAGZBZGgeP6SGpY7qBfJTA/L9B9ZsAkAiXi+OrGT7
Ycf5PzktPnIxcVgOXqsWUYW1uCqDAcK2rFV8TIU9kBpuvmcf3PCEipes868dRDFjnUNhJ5clkbyN
IKxxQvZTssrVi76DjDL2ZHQ+LaaOKDcOEb5jy9PsPsouiQ/cTcj7z3uw+Hf7UvMb/aPfO5C/XcAD
mUs0T412T34blmhKatrknG/PVHe/iYiuxaXM8YM/httqSPpzQYqPE/Am63tCYDdGVrbDLzpoziIr
cwQgcZVsxCRWKkIxnRc4uqSWtqTgkrE5yhkMx6+3QW0x0ryl5Yip4azY0B3nW00xQrk3fMzqiS+N
zuu/I9rrMeo6MmQ52mW5qaPKh+Aae2WEduO815Ng2wxbuYaV2zJsCafVHlHh5a7UUghc8UfHYHgV
VoMCw4SCYhDFSZSF4cxcoYx06pppJJrhBjyOW4vv2OBsn7r/TMdEjLkmOsORMoHHBFaiAU9KD7au
kD0fj+OIJ3GzqZKK94q4RtYWU0wfrhvC4mTy/lj/VhEEfqxAiiiUmfV1Rh4hwJxWTVMD8b00IDdp
DH3buqR/r/TSiU4Q2BSjQJS1W79HnHIFA/EPD7ViXR927NWS+yO+ROSuZuR0sULgY0EzA6Z8D8Og
3BsBwEJ//U5YFdk9i2uR8OAf6GB+UxLZuAslOJtDfaeeJbxujOQfnMNhjp5VX8VkQCHiMLmwtovr
M5dklzXRiwu+2wE7+GCizXhzebVeSsAxI8SK3WfsS6pADY45n+mNxtGMM6Q2vHps939uZUfY6Gnn
csPA1dIrOA2ITBqqwMjIdJAcAGYvbDnkY3IJ3qYbrjZRVT2XSq0LSaK28Dl6oimF5jpF7fBvBJnw
hdA9x6s2IWR2BzBCXBzrifcrFjqdtN0AKPkoYa/ldPaq7ieNGAKOxdgsGn4Ti/8EJN7wWEJ/wTFF
UnV5gHwFT4naZWuA/OwEzVrQaVpTmXBmuo1jhG6ZWOP6uDdDQYkyN3LDIJpzvF9dDj9f3Cw8TWWl
GcUjebnUmEPPj0mpkGYEXLr/LQZ0SPKiFbBoVrHs+OdbHXrc0NXCxiWfH++roL9LTgsVDLfV2/Zj
SZ4NJB9Kz72bezh8Czm1YsGbg4qGIoe5Gew8tiG8gKuck/zf1QRtJCFoquHBgLVY2iUMpqyxIfvU
rg3qSAsCQaG7vIsbffGOodosWd67ePxDy0B5kLBHMj4Uy58BWN2uakZYuLygtYneCbRx3lkPFWPy
cl2ojqYTV9InU5yU6wz1WGeJEewa2qkmwh4mUEkYVwu90Wipnks611vIr+oP13mO7kXI2pDszm65
BMtXtzuEmpnd+uRPD1imK5Z/rk7UWrmlhDxRQ10ZvADE8oYQAZMTjIQX2/jHk0T1wITYNeqxIflu
g5ruB6kbqrU2+8EFYV/DRW5/agDNMqL2xMLcJd8K5J89p06AZ5o2uF25GIkLU/uwHXFjwkeDVVNH
yFIt4qsCwDH/bjjd2/6Jtg4FZ+dAwCaig9TL0N5PNNCQddItBB9uw7OcFM9WV1XLVrK8K2P7oYVt
pIIAJsqFcDoF94kVmEYb9UrsGt42w1UhKwIzEw43ZqoHbqnpZhbU+AgzcsCFy04DSi65k74K+oqS
jsSVpY9FXt4kSOcDoGCrLr5JHniMVgbFK7a3HqfF78Hm9jWaOQulruMyhVRiLHyhQjuW1zoXw8FG
AVxlmERvNMnVsdoeXJJW9ckpvlMCV3xueipUflIMyObTJFkKQgvm9DCiL7L4PdlCa75Ij3PkQR1p
5bDV8k9G5DdOxOff18L3w+JVAwSpvyDpol0XHmcF/cMrcwhL3nh1MPAbeCHziVMPzCMBylLi+075
GUQ9ubXqU+F8bMcr/1JZBzked9pxGFpfejwcC5vOL8JXn4Cmc/CeFEj2cJ4IBPbN+U95vlTcHR9L
kYk4Pdyu1WRviCbBM/+r/4cTm46CQthte/OnGWiv+Ac2fOuFuFn3cVgmDoF4xTO0NBIur6ghh3vO
N4nXWjikoxFV6hu+MMbC2K12W8fjRHmSVMM8sEjJEGwIri2G0AsA0cbkSHdRP/68SmxsnTT1wvDX
4KZysJicM4gM5YGVZOP/BabU2N9fSA0Pz7iVDQ+YDt4GWMVZED4a+DHTz7xEi28tAPUh6bFUrK+L
YklwJPA+vQ0I6OPkGxH62gqcAziPmQvHwtpnTo06m1c7FsXM/ZCwQvDH41+qapMsVdcRMktwSrR3
6eg/KyHqc8hLiCiPLRmc+FYhgJvY+ST8AJcViInpcnp/uWJbida8pgYMFv4j0B1NhZME6kvSJVlb
usDTjrAapaM2kjo9tIn9pzTPCtmRsSXEQv/PisueRtvz1paVI/51jcuiVWH3px2HPWuef7rpTROc
9CLKqzpOaIl7+zXgjG2KDvLINY2NrImPYieUg/cHUDzxUL8oz1RpnSB1krfAGyJrhAb0TBbN+HqV
DLGVSuXRd1ul7YWBv4FPkQU1u5EQcG21We3qMC8zp3w5FSDmtVDeQv8N89xHA9lHN3urKtuLuoBB
Uq+36fEXi2DnhnGv9UnZBgz+6mZCN0qjqJXxSWOAijbjAY3ylK8NlqPSGDQE7G68V44aP6jKJkO8
BqoVenakWM4IrMp45sjXIZCxFsxIXcp4lCBRk751cQeK5V/41jdxFSzjDlFINuxGaJbrtUlgtJja
Nz+m+axOckiR6aSfkoS389DxLWarW22v5i/aYsd0/kDNAsLSbkOkByBDfF+0CrgdlHZZK6sleQgu
8nom6O2yZPy7I4eZlWvhFHsE4UFMhjz6KJxDgFd8ut9I/6LHQdPVQqEYHJogClhLkPnBukGa/Lcr
Y1EKqj2QvK8wwzrKauiKRGbaVQgg3zzbVA+GZTqqexeim+q1Sgmkzsp7UeizPsWZhaN5TqxAkn+C
hBKCf6OSxrFEKf1Gfeedgk5zqJZ+kn+nJBrIb6cZ1CDb0hRwvW1TlCdyWnz08aB2blc5KBGjCAKa
7fvLEUUo/9l5OO9KdslUbHWgZpq/ryDfVdtzHj9XN75IXmtnUcHTVvMjEdkXTcAQRyR3CnO3SnpE
HiEXjjoLu6m++1cegEXrn9SIB3j21CseFsrD3IJjdi6Cyjpgx8tzAELJJapZgBi2hAUV7tDTgN0z
ssubG8oQ0cYMvYlG/Al+RVOfKuy4TV7b1YKcdhHmvkxBIMONuXBdmePc0AfiqRVj9Q3jB1/Cx0iv
1KsSL0ocAJKmvLJen/croSy6RngIFr8kgCSZK9UYRMFYkmUgUqKLjYAR5Dv/PcSuZujIA5SPKTsk
nmT8NQJJ851/geNBBUmaX/rVdOSp4KXQWjZELOK4MAxZiTTJqomlD8xEIdpwa3DXqa2xM4+kcGEU
W/+SPIsNkeAVILBUBU2zYB/weG3eWzjge08fztzxrgEy6OazVzbGM/u+KJZo2VhNDJ9kV0jMn94N
t5osMToXJQmXvJVsejzzwPU1e7d2H3pD7AvOR+h+Ru2f3ZYLM3h8ZQ+z+goAwsueSeJeS83KjelT
np0cth9g5hVtYhqd9d6CUxCmgbIFa+Fw+uUP3YwrTNKuIFnPFlnf1soss4+ilMvViV+d4nagIZRm
Ka10SSAqBpoMZZK5tYVMYTmjVTyZh9mrJKXcCyqaLqB7sdT4wMy1gGSEdZRba0Q49XasuxA/l7c4
6fUZBd+DU5kKgf2PgKeRUhVQdf2/itkdRX8ORJtfjHIdPZKCJ/81FoM1pCjCt7npqEEqwbfhdiMF
zUFtk5Y9Lx2NwegPSoyDLUBLfB7ic57fCott2TlMqjWptEcrJOODAN8EBW5Dn955ptbwmFimIYcx
EbUPioALwVrhpjTiP1zFoiLN352ofCwtJEU8r9k/YBkcwubEZAIN33Riox1wi3I0/CB9RoHLGzzz
N5dhMiWz5m+ONY5JcyQVEV35+fTsdPG1jOslgX3cO3xX3NZgGyD3IUZleOYsF1/g/l2PoyGXGYk8
yHr7DTKwNmAE3jJDFBBdcTyakPMdVN1nPtUVBDkjujt1cXvbmWJzL3j1NNaEOfK+h6So+VMokW38
t9+9EJy58o/ZoPfIexx+GZmiFhwlCS+AefP5Jc1MAn2YP285Kj3obP7Un0CXLWdBKhR9RIohkuzG
bU/swfxYAuD4AM6mpiyYxs05vcA6ggJzQ4ZUWaepH9hipmcbgYT/s/fuKlzTCeStrJrSXdKdXHgt
U0QqPUbK3nyyC9g3ggxYJ1ygIWYHqGHiK7N1hMY8T95XB1Nb0PETc0jPGWYJsn419XtbotvZF8gS
kHrMXG5mpz/Utpey6We8/KQ12f24TRXyLQwSAxGKIKsr/I/1fFy/y68MBiJffxgWAQ6py1Bn7LBV
xRAuQC4xp4Ad8+Kg14Hw9pioQAQ/ABkBnKGyZPUP4xhBEieO8ajutJyasxLlndT4Z/r0uwRSzobx
PqtSfg+Ausx1Qo/40a86Qh2xhgmhewEVIq5jJJ5tnsOtXTbhFJ1jxmTKb3IS4vp1olgrF9ha1EOk
0TN5FF+x2gtJEdfBHMeVXt0hvsM0YpCd+T4asg5xUTovwa8QALQfMISHIlK+MXRJObIzIVbvk/Sm
gE5m/4Z2TEL72xqD/pzFYg+y9Rxn/S6AeQGTuoLpWm22Wqtya7kKf/S+hW5GkTaOEdNjNIJSwIKr
XSSzkUm+kBmNBJNoyKSitNOhyy/VVAXQjIhYPMJvNGJXG02iUzHfSZ0inOcYU1wrT0O7F/10rHOs
TtS7duSSytB6g9oXDvGZ7LwWmoKcSgBOsFlMYjvLKS2SH4D1/5w9bydfcdHlErji1Gbdy6gAIRpg
vNgq2nlBvoiojG75c78K0FrYJGgjyxrzG5QQ5SP+JJh7Zf8yoEf/+7lKBo86p/rboetcIY7eY+V9
1KpI3SI7Sjvu582LYJDJ+P4BmALv2Xq/u4JHVgU9sMo8YgpNH86uG8xwGBbri94tIyzfAdnmFYjk
UhBMlUcbf8bP5fRipbNZC4hpq3NrkGc6C1887lrQEkXJ7Xbsij/6L4d/2K7fEBVO7/c+98MmKkwa
5A2gXFjRfcmqUxZmw0/kphJNMqugsAEihuA+w6Q78yns+ZOCIQfsTkR3DWAd32HzGxs19nD1C9St
QD/IjgyFyf69FHhqycth7Q7KRqBQZGksoo5jhp0iNNb7f9FK5t8cvHw4UixbTx0t8DBvHky6oR7I
h0yLyhu5ZtoWo21NsQ7S664M5kijFNo2PxveAam60Wk2SBiPDqF5RhzBVHuwYSnNq0DuQaWz2Yhh
q63WnaKhZz2VGAcbdLkh6PDUqqxfskxRdqE6VsPVifWnPn2gJthWzGzKrTOI5PWvnttFgkgsvzAq
8+Jx2TwQ0k8UqOnqa5xtH7pyfxm5g8vF30z3KdpmFaIYzE788qkUkmKM2t6U5w9qgvJzSX8Eeqa0
mrWJwxK8RUJegBBq83sgB9ts5/vykZTgCP5ZNdmjXRzqK6JTyotJ+HIY5Cpccu0yKvTHFhT+Mvvl
fRnC6kNIazb3+QS8JlNUdQHndMbNqT4sX2clsgMfhvVi4hmg/veCTN6Yz6FV2NgA1zpjoFjFgD2q
zZN8ggXc8lanW4hv9oMy59YJ6SVpbP7RpJJITDhLJCqAgNtGBJvZeF1hpvZVf21vsjc1OYKbH+At
XwNjOH/eiEwFkCSB61izVcpLs65WR92XOwY8ukbsVaXaOdBzcVgizP+AGgIsSrbyFQzJ91xoqqC3
MPzFlea6xCKKCbb16V0UPapSVSKOOtv/RXGO0oaqUXj3FyhXGs7SZDt4V3jn2agTLDj9amcukKjb
eFEeeBfIMC1kR6r6EGAkJBxW6zNBdiEjso89C2Yjjy08XQ+zo59gsRMJh1/SwGL+mlZaaJIOt0ZA
cKkjHxmGjsXd3hsydCC/nSHPEOeBs0Xk6+ljetjBS+1ct9t449Bt0/6Af7RDtk4RbxexATpdQtij
rLWFs/gzSXOWbY8T8GF/ifLu2czoplRUSXanz8pyQF1bvQqe6uFPA51DepCFnpRFXVn3o/7OmAHo
4WNzxzrb37w1SyqAiVkQ7YOUzFItl46sy18249EFgTodxy/eTipBDsIUPesr2U42yGl+eIss5848
zgAFxOpofPWG8J2O6o67w3lhc2L86ah4YEB3wGSyIyS4fGaYMH8BFuwnUp40e9ziN5w9iQG1ZJEG
NvvdhGs6wOft0GXQIcsXwwMRIUe7JH7MCxiSepHVE2F4fhIj7iXo4lvEd3x/tJjxvUtE/9uQE8MQ
3YHAyZ4QQSW7rudzVlSHbq5kWR1yA4/EC6NQXK7klpR46/vWY48ZJkT43J04a8xNvaGWSWCmlF7J
GQKiVM7NnVsuvv3P8QWqTQ4v6LvfxVQta6egfuR00D8oH9jUqDNuQGMsbQ5HzWK2vd7HRdwk/A2n
x/z8ox7z23sbu9Ol3Dg/OjM+2ADJLuNwdIl9xhWjThfHeKitz1mlgipbLyNDoZwHnxk/0QbXN9MC
5BvpdV5LGYFw7zUiUJ07Jjf8REezqPKIcenEpCcr/1J8qmvVjbQ++KFJtSDidzuN0g1ekHOvbOfn
KzrIhTHSfiZIIqIPC5n/d4ZFMW6pJKmPlTq/vuKb+lQM/LfHUV6NXJ8V4KCkZPkjys7OHA4AOHcv
tUDWftkHS8zbsxWIWgYTkOTt1vaI05pXthyWSoNUHEycep3IZLXM4qSIT4/TvkzyFEX9S6TU0eqS
DY6bUxmeDp2wTwqumsB6uLTtmCoqOLuBevPMwQPApZ/SQJfGucpROc4A251rso/nLy78bmmfeAmS
CxX7gPLisbXN0dAkZ+7pq9cpByl6Kpe6hNL+Bmd+4XPpDgInAht1+q0p6JdxTZwuUszkAXMRtn/N
EHYLrjnG38lUL4xFEfBanngmUiZzsl3zcXP89swDhhksRJr1nvUidprTXvas55MKiPIeCtVtU5UD
MMWFXwWUTqz+J0XdcpSoQPtxixGOCjZEMTLSpF7r36R+Z7Ii47Z7afTdqhXDDhSv/mDIQXOyQmIM
tgc+5TshIDpRHLPRifNoeb6bD5hNuVjBG46xIPUMFpPG4JC9tHzlDKSXUxRygwaFqRGVA7VlHGcW
DcH9D20L9B7f5LCZX2AkrEcuq1+Mhyr3Bw63OyVfzq+uq9g4jhIbSeVPg3DJt5i1NlS2B3t9zo3b
L0U86WkVlKROzjbScyyj64ixE+C1c+80ZjMMq67Jeap7U/+7lgmnr7NrZDHIdJXOP6M2K0m6+Uny
vg/iUPFJ9cd2iBiNBuLrKpTfPXxSDrjOuvoX5RtukGZs+XgupK+8ZkPt+N6nV70W9txuhEp6sbgm
ryy5MyiKh5cS3HGkauzWbpQ1OX699Kwp88E0gr9N8mGJKEtd3jc8JRzov988rVUFGulktaszY+ld
j5tQaBXpXlhroLh0oR/42h0voGRJf9f/7dmEiPHYmTb6K4PvOH9qbPPKQ8vISi/P02LfhZwZ+vpy
nfrK9zYzjNXc1RmCCPBntVz6PJtzPr4yZ0uu+3VG+t2z790MhYVI2zE5Lf+/HkYMGU92QOd5xQV6
NB+CQ0g200zzrXS8eYFdce7ra7HvFQeDTtxOGZSq9jXLBxcQNdZx4tGEthXtyH1hQhk2xjzCHyyD
Shpr+W0LMj9aJuiyDofWXhvM+SUwr/U0oLaaPbNU1SYhiPED0Lb+3hKx3xiXmoepHcwurZVkiVnv
c5+MN8XE8utpt+xiCiqG9dmkBL6uk9ufkF9UGWR7QjMiIqQAEOSZ/fj9kXX4Wokil+SAkTdDE02f
MMtR0dNzmhw03gVQGHhcuHvLGRy1qj/i32PCexrx5xpcEcvby9B/5TS+6u8myL5s+rWTg37mKPby
HhULqtR5aulcDZNhpX6V0xlec7cQOQ42h4KM2f3Hcgd1N2D1wQat/UJ5Z6NP5AQrCe/OL5KQ0XWP
KYo/lDo+9TngpIbT8zH/RxW42pHOJ3f3Kzw0TTwjxfmLlDJFKrvqmpuV7ffFh4s4QoajR1n4GJ+b
tjCvYpk82mKw9dTLCQ80/ObjgGG/yzymgsFfGEGlZPkL71d5649waX32NOFzWjDpGqyHtffPK0kY
q2FnEAoek6teC7EIdHTzhzwCPco5Iqsa2DGzeFBMAPcjIeU0ABJLSUqI8Zua3e0oRuSyv5Aj1LMH
kNwtn6X8ObCNmYL+raSIpYFIM02dgtpXpaA+TdU7AqbP5OoHdNJUUu5QlL+NX/hUjDaiauMxwLkG
R06pY9efjCDqM1whvVfOvCOZovEVnOm5eb32K6UvuvkydJwbQlvIhlXaVKElWnqSQo7Q2OnBKtQR
5SOMxrGrTvyzqAuQUh4kqh8ljxWqul//IWYBSK2n4XsMA8dvZxZVY6qJBspQMyKp/k1DtdI/G+bU
5rUN852z8nUV8bCZXEr/bIk4W88p1PA341LudwYd7NzXgnuMSx89J32TAmXeMo6Ouy0XrP/83Gph
/VOHRSTS1ZUHXdembKIOnULUTr7ZNeF0EEwlSjfpCYPoM5PwD2S4AcDe5+zgyNoBf+Q8Pf+d6v3+
fIdCpF4PSB9U0Cw0ldyjdiIs+O6QVoZL1OhYDtkaxDx+jpZiiRulwXzJcGWUyjAIzIkzR67z9bl1
BqE1vhGQ6rQJDXe1Y1FoZseOHNuJ0z6zLD6+1mzXIO/EyicHs9gttB7v3P4gI7cbihdN7c1CyN8a
oqcS2EaHi3s1ufe9/spdwPwIJ6OP/SYD4IT8ygDs/QWjQmA/h/2HDk7LerQWHjsRvJ7RYDD32vRr
kj9hwri/0guHP60XogfF+A12zvtilD+t+wubMbeKk0OoHob5bH3ODJaA0nhLIIf4WFnPL174sBHt
9Yrs5pE2m1yZgxzMf6prOCxXvjYnRcWSW4+QwJnSffVQv7fki8CZ5Q5vst1UQPHMJgjwURsmxAtp
lnI5/JHO44Hyd7Cw9XvC8I3QkGNNt+V3SS9b6XntmBxLZxNI+nCoSOEO3r52TVeO5UDd7v2hdxzt
Zx7uWCgeWfO/7LOFO0qZic9jzaY644e6QpXTqxFg3DdagL0ehavW1KFWIr38jEVxZDhHm6Tq1KSN
4ILrpDJOZZ3CceoALHKlIP6t27+oI/sp1EZZTIMgHB+QLh4RH0nxX5IjtKD2D4+8uiW/upJcb5ZT
WZWX6hR57V+/Hfo4uPLYbsBxFGI4TtCBWe1MtS2l0j+9ZbdWFDq2YYOJJzLgkHzc4ZMaioK6qZFm
be+WwVH29Co2osAWFBBahtIYUZBgt5AA3y7PETWUTW8F81qOUBW0NhPB75qPlmPpjcChHLvI6rgj
OvZwGXpXR8TQVyC9DaSa8EdFFhZtcMpOZxY31CxiK35SzAN0/dVtmEN3cYCGpWC8F6t9KpA3Gn5D
I/PhuDR6zCybFigfG8shAX/Ty85WzQ4dhAqxVpCZ9QpXB1ThQXjKtmaJOtwrFdASVA9cFNWOaBtj
giAQcDz1lBVQkYk2q8eTkZ3b3OeLDtz7aCiXklVFxTwkh8X/h//f2xz8O1d6PG47Ga8628rQ5dsm
JxnOEruE4xUkwC6l23Exo9moaNcrkaMISWvZqQaTM5A3adqUgAU6v4bwdC5/fTbiHdoLjLA/A0n1
wmSgo9d3AoQ6U0E8csP16wg7OO5FxUfuilVRNxXmHfL+K/aclfTog2rXkH1CLK1MUgLb+ccDBXtJ
zkythqX/wbBwXcp0Ti4LsFH34RXdItyppK1mRZf6bRSZp0ExZ9u6xul6X7BA9ocBzlUbx144JuYQ
THUF+5yC82dyPY92MBij1CM2w6fv3s58mfv1WLb+AJCbp/65vRJi8NQpTlNXCXsgPnVFxq4Ykrme
47LlzyXD2Mo+X/uxoKYFbm5XGIIFlJCPJU6+nS9CPdMhrs5ob37fJ0sFXrkC4xjFPXcug9Ewx1GP
U2F2K4aRl7MkblmINlI/Ld02yZDuWMx5h5UEJmGQFJS1qeDsypu+citxFjSlY/EkI+f9PuPB9Tny
gAX/gEJoNhmGn3MtaE+gqPtTwX+Ke2naTyDJJ62amThKqMcVQ+/nooPpLyWkYe+9l/1zmNynQEE9
DyDkRInhwI/yVm9GA+7taYlkL70lz45znCeIBa1FIIXP5SRfY9YOf3R3WEGM9/7AU8aO4s7UGFwJ
PAL10pHoyxGri1cOijhd2PfXeOoWWh5R8sATbTjJxWysYeitspVtCeykWTTzetXGxHQZ2OXwF1nv
GLujlfkOUs4XpUu8E2KZH2gJQ8ztAhrgr5bj/8cW6V1fycrRI7YegquBuURI/MALZkMhUMCdIEWb
hfd1+wpeNxndNmc1bSL4xgVtgO1yFJiQHqVEBPyLXJ/8tV2E3vVJk8YLILdD7YLgH22nGD/ph/mj
oGldrkXt6PM8ccO1AHUqXfTDfN3CI+T0fqXW5EgTPFmPI0yowJVCQR2vUI0pzq84k26cGC+iD6FE
7gHyKQu3Zo/b+8Ngao23R3Wwamqs1+JNhxUxktb8s8ZED9WzC7hHVkZbIuzC8XrPDnNQVNDQty6x
Q9oos/pGgR7+/0a5j23lYKCnKndM2MGqSAL9pIyyBLwsJJXOE7Cgvc3UqJAS2K0enbtb4LUpOhs5
rpvjktYkpSb4oFFt7OX6qT57o2x+nHi+ArgZWjZzGNo2axABhHU31AULWqBCoF8IKDvZEQuRUDkD
3diUO38js8SHiKbnLPcqFvZTVRTuJF3tuGlm/0Sl5EPQ4Xfgpqral5KthHOqgdqawPR2gco7EZN2
FFZajKKlurC2KEsZnA5lHEQFfaQiRwn6cU4U4knehqWRe1wx/AL5d3U1eAkHSZSHrgqQ9+xLF96j
gdzmpzG/a85izBe00EuuHnNQjpMDamIXWyaYQgHqwPeRM70gf9ZsOIBeHQT+1aHHJ5diINsPr0Gx
y8hLWCgp0FFvF5Icumbdi4oOlIDwNWiv65D0OAgzHiW5s1DD3WtvKiuIkzVZOFIWvaG+bYOMgJ3P
s+Fm97nmUFn53u+1+HOBJi84CzPQQMxSkJwYhO+NULHXI75UKqO5M8IbhtFx0c7xVy7X+Yfw9iBn
YBdbTVa7iJXmPLUXEY06T/PHWN3QKWEijH5SnIlRUPi3hJgj6Sz+UATAr/Q6MEc3hFHRQoe5Ovwf
/3sSLXuCM6ggXMEFk3CWhc8rv/NfUp4Hh7WSi8Bx2/ZryEm+0u8FspbTt+d6V/sYXBCnCe1YFRJ4
ObZYgc0nbIL8ibwmvpE+p7Ayk0V61PFC+vOZ2DYDHj3BQ3LmjYXI2LOY1Ql0uTxE/KtWkzCbu86R
9gLpXBXLqy6qXjYoAojCr/DOSJ5P7htImI1LXzAXaWSUp1WS0Lu+Zx9MWa6LJKSjQvisMCYdav7O
uhz1pbH59e2NyKJNqMqweuT19c2E9tBqcBQaB6sucI4FlbdiNkFNFB4ANXrYhJnDQuPua+NitWN9
QXBtv8vxRBNldVoWu/tGZ2BXG4fEwhrre1F3ckZ0qWUPYdV8EzVXY8nmR0fifDGTzY61kpL+ZyWC
EStt7NkMwWonovB9dTlgKt1D5mECOK+f+pExF9CqQLlIRroTMZUWhjwy4c8jdOeCxu0AlzBnXEwD
JEs2p+ND8oMRZ//IovsSGzIaMbeldNs0/5ycdc+Z30pFLTfZxbXddivskCrqB9KBBqpg8BfvtXqp
wEEvp8vT84LsYb//IXLqBZa3uOuSss2nCNc2wGDRh3H+GclixmTzENkfmq90wmi6O+770pB+ryt1
d8P5UM160PAlXX/mTOB/t7/6i8M5nmAcTjlsYy3mm5wfF/6uuloJbOPj7BclcLEThdWflEdnzHhb
3YaGvWGcklOvQCrsHseWEEK39rjvSxFdV5ZED19V67NslbEv1lQGsJs9Iw/Cy3XQMYj3+miCCH71
Mz6Jd02EhbAej+Huqnbqw9dqi9knQrteLDPgjGHaaco2TMDB845OhMyx96oPLBzJVuj6nCuDVS15
nREZ8f/dy7WWDj6YMjDO5/nI233FZWuCr65MbBd+Xa2ULg2dyApeVfcbvPSZI2jWG4R2x2ybEj33
3hMmHHpUBeeES3wKJik56gpmg/bY7FskZM7SGpSDAQype4wkd6Q814Kjwwd4KY54aTgjoVPue9gf
ul2R5SwP4Y5mArPDELiZfb83RXkPmmmN94/+ewvgsCTvsMkY6GOLuInriyxoRudKhOKmuObSuOz3
m9gQAXlVX+d0zatQgtZ+vGl9vxuBOLSph+MaCjXOOOiTKuBwRQ4gfFzaYKUBtUTmNZx566069+hp
3dY4pEkgXWHnT2KbZ8dWEGjiXNbggZoO+uZdEnmnP1xUqbreUGkB3jqzIB7kke9EhAGXDxdycT/r
WSRSzq7Ck3SPJ6EYvJtpzgxNP/WCdbND2F3yMlRhTeOydCocNQtMJq9V1zpvN6Sn68FAUa20HBLU
DC9IVoDYZua2pWMpFbRigEFzvYJ1ABdAUoFn4OeGKXfuvz3JtIScdmXwV2VscTEUJT2n47yZhV1g
/Ti0XpmOaOYvofw/ie7VTVJC7d7EBWX9SZ8Q4gjYOyDZqw2lJpxy2ABOHfvf9W4af3xqN9ceoGVZ
6I4FPynXbrdW33bTnCuAtmB0mU43U1yWQ6a5yoaDVtigglYgI0RTp3ay40/8TWsi0Y4vIoBjmRPr
yQOe8LNRrbe6SyLVHCo2zpoKs7JppuhXAhqgjoVD7Y5Xv/lL+GHPGOGE+Y2hpPPrrwjajpk8g+WQ
iJvjBX+YPeGVEaxgLgcJVZnJlvVTOaWWHHAnBWqk1r8nXuizatpAev9Hz0mHy/pGEZragOW7K63Y
rM97UQOXflnoXgplVONZC+59QqiOtEPpetpoaqbyim/ap3Uas4xbJvee/SGHJiASMH886S/qUY+7
6zV8r/rhMZ++Xo2EGbYaVhgFfU3QGfPZYtSzmK688+EvENCXUudwwupmMaWaMGLdatIKyFixNHE+
5pbVTp+We3cDuQbVIFvsRwohuLCfEFWPD+6NX4B9DZYsm14DbN18kqQlRhIbePmHxnajXhVkJ7z7
6kyAuh6rQ/NuChLwBvaQkuMce/Znn3JDvxizTKvdLqi98s/UAQSUwJJatFpP0qBOVEpwmrl6dVm7
1OlRGIitQRGU/mkB7m/xnabaO9MW/E09/9mrDoeK0dI75NoIUpJxSnuuziScvC4tq0zVxcHdxXgp
MKEuxL7jETnSGoTXePT797KFIU7ID9yLdp22aZTqKr8aNnkmgS3VyKCDKNlYmfPi438ysCd5utRg
fm0daUoHVYfD8lnEF3c6Ypi6PqGzgTiZ6MNyyI3JDdUF71wLB9rHX7bDXCMzd4K/i/Jqd35f6R5E
XIwlU2VhTcSLnJn7Z4EEyxxgk8j5CjnD6m+M19QfXYOT58oM/UeWtYUprgBY634Anl2CMlLnRdGW
GGJyaXV0ePLUCd1kaEaR/J4lMDpIeWCBx8sfdlkSNSEvePzw3aL1939AkrpUXhoIZQqxwiJSKj2V
YPm2K0WFDbRX5KY/TqEBR2jbg/IwAuOyi5PJH5QtmMDzu2dBysR+pLHOw54I5DYVYryCVVq8Nqip
Fdnm3iDWrqe4otmbYdf5QVGtsbqqptbZhf0983FEMc8n4TQDn5u7fMmUXyQfyAm9OxnAn1AQsynT
1rblYrWIf19jrICALIMf075a1jiXIZAy9SLGSuBM+Pu1c6hDPh6ADO8IHJWkw9Eu8YwyYhm+sovX
ts2uMsAQIzZz9Yu8Ex0KztZ35n9K478XQwfHRaBrfQCcIUlogmX7i9QSXTpQd0K3SAYkKox5Gnfh
K/Y3ucU368mPt7DKdFolKHHAKVhDbQCxvfQUFRbZgiwPMZbt5XwRA5tnOkpDfJw6gP82s6AODQ9U
fgMFiHj5KUxv3Drzgbvy0L6kBjNremKmYUYUnQmGCU12P7v+D9VqLxE41ZAfIwpxSlcq0ziLirPf
nhNisEn6dB+fTSHeKcIHuheoxjrcSt2tW4fDESueot87MN2ZUDDrec5NqwNptEtILCbdxbE+OQDu
OXQ1mizCAz6lTixhBZLv0phcH5Me2I+BtydekWf4qr8OXXNgUh/0onNmeUcpEopYr8oFy6MFQiXf
QZ+XjQrqU60IygXO1W7mtzw9fQlnPPuu+mZUB4Shnsle6dTPu20yJkMc/pFka2PFsu7/Cu61r531
xuUtsHy0wW2/7tTfN1HEWct15oxVzJtwU92haZARy87RiTOKoBCizzDCkOYRH2Z26jhlegK6cFgJ
X6RtJJCE6pvVGAX/VIQW1b6dZ4K/UkEDOmxm5xVwRHy5XuNDoUMAUa9fWl/HLSkWQb2FgZJjQ/EN
KXDMTFRnvB8wHU+z66MRHoG0I1tZluOcy0DkfH3xb+0ZPmzhlrHq3lQJSmDUjTOyeK+BXjuihkNM
je5v+DgrXnTSu8coZL+VV/09C5ewzulP2+g/12a4V9jYpI7nRU9eemQkQQ9YuCgmd42yy1a5qr1J
KxpvKsNGTTjwY6fHw+x4GGu3i5ElMlSREa4QNYGHvvnxKrU7RD2GQoCMYz0zBwIbY0CP3KTFxGz7
v6OntQPnwKoZXvhPxIxcjCcJ//K+ZnxQ14Z0+TKqjv7M/d3Stc7Dqqi3u6sXVYgafJPcgPrNTAme
sx9w2ttbwv/+soVwuZpxVm/TbLDsuu7900Rp7NblfiKag1ysd5yCzhFKXxyIdib+cCHi7At4NWgn
3pcUu2OqRdBHYtmfXiT7n4Ws4zaOsME+P3uctYMFZD8YyVA10a0Inp5sjc5szGRCFEioB6dy3jTu
O2IkOg89IsuBzmX2fcPXs/IyC92zB51dNcJ+bjZsZki4gISCnmyfeCR0gU7nwY8GsGiEcpEy9yC+
Dt8fdCS7KTSqCblwaHFMF6ytDi/TYlPeaMLcrioR6WykdC+mvdXzLx8c7/FMyLrnzdONZuZ7UHPo
nMj7Yea0qSnEGiK6dhhcOtEOShEI08hgaDl44PWX1lASzCMOlKmMLfB1Lwbh2D5AQPL29QtWRqQR
q94IIMDhMH+NnGfGVWNkzekr1nWElK1QIAAQGE8WzXUEpvyITNNm6TrqwicDuJsnUxyBbzqTZ4x7
iXyCkeEuEDsq79tI7iR57cyzRwoooehM2shWqyOLRJVa5+nzLv4e3wT8HYzaSQVVLgXncfv/pnm7
b8ul4RHyvqN06xz7xcNDVbZE461nOTIVqn1VKhLb3EUghbUMYch80QafeezsuA0aK9p2pASZZHRx
yD7+gjEB7pnE18P/hqA1umVAkRbCOLO9JkuDYcoAHHe8xihRrh+YdYOZ5jPjvSenFwvY+2G6Nmmd
OYBTMeYF/OrRfDi33GknmfFzKoaWmIdAPXF6miAZBzXjQMbzLm4DndSxF/b6moNGWut4D6zSRBdv
/7r91cIAf+SdaCqizojLiy+AYLyd4FQQFoFUYFV1Hr1xQu637r58Od5eLNPBx0NcAsIuchCE/JhL
O1cLu33KG5wlJghs6Gw+okFDVFWdndop9Gm+yhmLP3webFjxqXnEDN7E1wshA0AcMmpAj+08zC8C
a4qj/BYm2iLtpvhd6QApkhuHBwawt5yRUZYgsTdETq6q4+U0SbIO0bcyKNUEo/Kg3SQ20+kfKN5J
ivgBEdhDyWIp3h87sWrtTTXTtKX9oZkjIv+bVDMur6zGNx6E0ffYGFa2MEeAIrtjwReBsUhWwUCc
YFYXaR2SLbW/YS0jUaN2KqfPWKvLwJWZnkWkZzdsUxJ6eQy/wv+4x+ROqQaZnyz/xemKrdb47w+2
aU1ZERZJH4xwCBXKDa/n4oalfvTMd+YZY1o/4QU6EiNGWr5wkdxwoGMZkjyYbgzQkhnFxwL4RNjI
/7w3wByqH9AgQjxTAxrAv4dKsNNqbZ1IllJGh7vKBpNyzLm+jpyEcuA9DgV3ioORpWwxsysMMvKq
fRKMTtZuRS44+95/6w+H9PI+7u9RHC+WoEZdsvwOYXn34kDeUXBI1bFV374U7RGNpKyUuG0z/s6Q
Ak6kCVBFN4z5VsSsORa9dEWiCIQ7oUXquaLNPjDoJYZ6f64cia5/orpY3MMAIFgbC+mJ9WjfF8FP
SQ0XhkSO0YfjF2DG68DaXT4Yc4TVnYWhORJuEFqjHXVu+6sdlmmgdZRoxr5zkvh9HXrpGwDC5QDO
qsyc6jChgKJDqs6T3Ei2nTHewCRgqLCtV6zyeUqskZ09Nvc9nc8/dM5Lku47QFnxA1ESLmvIon5B
baEIYRTDg5S88/cgCklfEOkwbeEqGJHb3s/Ejgu9GK5rrTQzLc74PozdmZdd/VAax5vdkiSJlKvy
n4+zBhRpc054ZpmR41t+z79Dq78ZvTpClUeIJNy66+mepfPa87tFsqWDN/WVMISCeq7RtxNJArgt
gxOCnF+zCtvjGuWj1QCNtV9vOoEM2YExUmzRQmYqK568zsEI2r1LuAYga55gl0oJn80RqQler091
0V1fJQ86mVt9Mz7WQ7ERr4Dw201H2nFw/lH4aTvsoJT/ahirVFDUVcYIPwRJqkz1p4A0ZUG4SNGm
rzuJXNz+F/kDfgFgJ+rLWM5M0I3R8icATBVt+lICoZW2eiJ2ta3oHdFiQXhQg77e//vyebS3ydLj
ILr8CNtKJ4AXEEImfO1kxtE/9ib4Lp/eRoZfAOAWd2GEAn0qr7Od2uOKHh5ygjgrGlrHs+o9oYwV
YdmatNa/oPNnO1Pm0gECrUlAa3GzPiiE1rdIei0IhSZ7/3xoIp2byHend0gu2+N5NYhmljOQebBy
gwKI6Qq0wxMkrSr3PhBCuiet2Vip2IS4767TfRfKRJbi4TPtW/k5qq56qu+38/OGKz+jGb78loSR
rSpv9PuMlMwsydVoMlgqNaNNjB28CdkXunN9sp/GFXg7TAVbTnsPjGrzu1+quPuLUlfTMeKWYh4i
+9ZxATgu9dI2Gw5eLifx9NBlT1L3XCzGFP/WVnB7BzBC2SrZSe3BvQRkOwGkkvahO1ABLVow5FkT
mJucwuVI71EC9uSKjHf1cWytMBwY6Vfijau7g7XL0tahn7jjCA1UCeaZUvNKmkVdyvQbDrLCyeFe
dajkf8YVHQP4QKJvqZgDN7fJnPkQ8ivy1ooNXrGcmefrnf9rLxAqFi/r5aYzvC+9tsgxtcbaaoVg
+Nv4tuZWt3RwYzTfokvpllQ+nRGr5ZyQpiLD96nJDb8dT2CcAsTzjVVcGDaDWDAO8UHlf8qxpWXz
Y13u+32+RpoBRHVAihvRhXERd0fm9IqYP1TmegeXT9QR601BCHHa4ouorIF/DDsa9XIHaCXPYytb
eC1dqon3egoaN4DWxBLuZuAxwCs3Nctvr4M6o/Q40tIkAtnWOm9wGo5TNolv3f2y7Ifclb5JuYZa
RAXhBsbWGJpKpvAETDNQer3hbeP15WMV2yeEFgScJrweejloFcFLVL9gFl0ZGWSUMwSQloW4ehVT
Xf95rKoxA6w4RuZzVmu9wuh0RuaRRwJcgdXeZgGzwtRslzjJakF+fp4QBxuogXvi4jUvGVZFymCQ
qKMWUOX5aFdjFS6I9mgRXzHehlp+V0H1U15AALcDoxA62BVxmCLsxo7alXraJ5bOD0CDPqwVNyTz
/qyLzJ9y/7dTpjEVkmvThpQBYfKlWPZaYYMTrKTjBGzhn8x32Gnr5ByglJOkLcT5XU+bo1jVYWT7
TuR1hzRFrXKTwSaNY2q96LYvH7xYIbopHhHUR79dwjEZ3eKp/O8qILZkY15BqUXfjeJMt8y3uFY0
YjCXeOD4Ij1//w6I9K+ycWOvRCxcBN7FCkPvzbd4dzmxmHGLE8E0LQYoWHjKNK6PNbJLK64IKe0A
gytY4AprkFrc6jyptbpWkrm3aiNdFzvDIzIDtbOhqq0jRl1kpPU+1EnReTPhQORh//8Ue0KbrLrn
LuZJHuQMjZO+ho1aSRGxwxCTfl4hgSVOWvKsjx1BifbKaHXvzfmtOGWx0SIZ5CCQHSBH8LMX7Uey
v77A0e/n5zc5i3T6ESBDFe8WiDqC+AdNVHj6oKLiENKXwnDdtQ8tPEuiMhaofjyHgFukXdINy5Vj
nFv0sAHu0WZmOb/cNmTByLs6cDCZ9ZYyAhuucVrQJiq1J+/08oGtYwYza/HF6KZBXPMYRpfZ4pqE
1O5dGd60oUDKXNGpxgoaY74+1wdSVNs3+OHINsGBStFOb1rkxDAknXKc3zm1FzJlOAqSKbQDhFIZ
0rjoYeb1TIdhIQko14MTDmM6yOZS6Bq70mWyDG/TXumViFRd35gILuJ+r7BLL1KAKQMc0uexfKTm
5n872W6K7fghdINsD2JGcJawpeWMmVehEs2gmBUPCkRZotGEtkVVlabF/oEJFOYAl6b7voFlInlN
gaRxwr6tQ6LZ0ir3lYDCd014sP0wAL7IMnMbjhCY7fNL1H+uGmFMAblMe9YMiHMriAN566WO4Q5O
AxRdospoWoMGitSSVHWyVCub0jLKfZS8VUvs6HZmt7kxiQk1KeWfZ8cYWWyALrz3MINSsJY6KI+E
10388JT6NqtuYcjuTS7s6f84jnjKNWSdGh1J5dhJxXqcHVwCStFUwzSLQ6hl7Dbj1MgtQBg8XjPV
pMsCOPOrcWpjHeoll33vHd5041JXYISqoGLHvKeKzOt+JDhMr5GB65/3ZIClR8oRKoMadoDii+Gx
4Y6mHpEE4Tv956CICqbiUVpWBdtxuY10DOsfYLrlRhAVZWANUP4uKSyxrlJsP3c6l+NMsbwQO+ib
2SysEw2fy7OUjPhr1cv1m1zcCDFfFCoJfytg1CS1ODNDKQgpupsTi4sfLPuGHp2BiuZkiBzDt8bH
TqywXSFITVvSGgn4HY1vhOZQUEnX9CecOGHOkYxzYIAkbs65tf1wWVRvxojnl+aU3tGLbAwXgaDJ
SIDVzmmP2isDy3Dl4Axi0HpcQa7cBWiVmPY0j+w+3tfuAcHerYox9o8ADSfBDmVPPPJcuNCcK2Uv
dnvoPmxeN+qODthhPTMySeHg61O90fJzFM9Gwh8VE+Xa5bkgIAGbViC2dJeISNd3r4GxqDu/nOpt
F18KztP0LCQZhQOQopo5t+OKLgxxvLRLGsThxaa09OmwLQ2K++TpOgQh8GkMK7vXtBOjLwZJkzI8
/bdeD7JE17URKk9K3AeurxGEzghSNcTHr9C/zi+MLG9ccM9FpkWvoDpcRN4VliYCGxyJB8tOW6fY
6ILsUMiCQ1PfBFWWJjSbJ//OqVhRVsASTJow4kf1CgvPty7a5wW/zdELWrw48zgV+QvIpmFzbamw
8eKIyTpATdsy/0Rxlt0VeMPj1WsDHyyxpUXXL9++IRb6YBgs8gvBI1dUa0Zms9FoUPaVrJJzWNft
6TqnqzONJblfX/oIPRYp+o1CRKPwGgPWM3dbgUuU/I6nh0Kbmx136XfhvJcKJX1YFbshx0mUa82H
WRs1lwovEzxjIL3HpVMPDEc1aQb3OKYXjWdcX59CB+YfZJ5GbQGIZ7lBziTqjB49SAubMFDuxfZT
ibaOtojP17rIuaeHAZIM1X3qCk6RB/iOvWsvWEfe/Rb7nGTDA7DYyO3M6+Cvtg11nx6a9uO1mCzi
EN0HVJuWEFJ1hSc18snFdiR+cfNClJwNs5KtEnoxhWhKXs4x//LpELhYQg/9adIaxr2wjSMcF8Td
N+Fcu/hGv2mz5pHrdvAEtofgG1cttpFnwHonkjS1tGSPfaLiUsx9nznwz0i9eek+Gxaw5Su2rs53
W3N3IZJ0Av4XZpvVSpxppzDa9h5bGriv3V0E/U2+YvtT0KYF11VqT6n0WAYHmtWrWFlGtOqnByH3
2B1P/+mAkIVTl/VB2jnvICnwIa9oLnPyfWRvk9n1NNGbY1br9031X8jPCk16UBtkPk4j/Ww3eRfX
K4dKsAL+FBe0Ii0XMGyGh3YlDnvAdOCiSd4VHNSL66DWZ8qBnNYcFTzU/HbC+NvQFL0rQ24uf2wX
l9IdvSZu87dILSszDltjaWrzElGMERd620507qD946/K5cWe/73DmhKTh1D1Q25WkXGD2gxIuzX0
+xYKIfTT3OvmeSmatugknqzIis4J5GGf+FY+DGFompKCUlp+8SrGBuOyf0CMdyxVbueyuRm/BVCy
9GEFF2ZmAhb8bh7FW/YxLefl2nBEo+LzEAAhBoskHo4SqcLnwPRSVTy3q3pbHFB150tbLdAEvdWs
ROkbqt8Zjkr5jfEZ5bd8lsfpQ/3MakhB4Io6U59QK/4bcyv9NMbhto+NH2zeZWiP8VhBpOQrfuUd
G5vS8gvT8vYFM4m5R3n51nA/bEAyLB7EVtR68le3+4RFUvGISLiUaxzdBbcOk0JzIZIDh8aykUCG
bZRogU52iO8AIDOS188+pt//6v1pC+iMFaIQO47lEDhns7oUimBk9Flab/50Oial1fj+PkQP98eV
0vzPrsjLkNe2nks/HE8cgsYioXH3FPqodj0iK98U0E//0AeCadqsWK1s
`protect end_protected
