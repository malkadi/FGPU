../../../../../VHDL_Files/V3/ALU.vhd