../../../../../VHDL_Files/V3/FGPU.vhd