../../../../../VHDL_Files/V3/axi_controllers.vhd