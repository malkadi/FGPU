../../../../../VHDL_Files/V3/cache.vhd