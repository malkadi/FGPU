../../../../../RTL/CU_scheduler.vhd