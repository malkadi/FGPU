../../../../../VHDL_Files/V3/CU_scheduler.vhd