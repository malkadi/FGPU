../../../../../VHDL_Files/V3/WG_dispatcher.vhd