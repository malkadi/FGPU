../../../../../VHDL_Files/V3/CU_instruction_dispatcher.vhd