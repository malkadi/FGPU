../../../../../RTL/lmem.vhd