../../../../../RTL/CV.vhd