../../../../../RTL/ALU.vhd