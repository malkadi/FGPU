../../../../../RTL/regFile.vhd