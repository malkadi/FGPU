../../../../../RTL/cache.vhd