`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
bx24XPMbQl0ZuYgzgnvmK2UJsn5v5rHRrHaBzymEsRVRAjuRN3xRCY+goyOwSGiaL5BZpex2sDSK
2sd0nljSnw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
CSRfZVLMWm0HJLEB7NOFzWrGIhgXL0zMCnVPoqKjG5Ur0+RK898D8TnT1vzg0/m9z9AJo34CsLar
7ajBwWmQaStI2T7HakgiApYlcuC6de1XuIEH3rZRMj/RWcjpTLbgkrbMj7lCzKzQdvZHARVRsJHt
n6KxqqDLGxMs1/m4zV8=

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
YDR4T6HZUUPDmkJ3uEF/8DG9RH1KIm/Soi0XWVOdqKCDBSgk2PKH3QgKdeu/Ygc+E4sEfsdQ97ZX
ZNKLn57bC8vQMoMyVXHXP/gB1IkATHDtiORbiLIN6gz0rbLre/0AWJ4pnD6+ix+zJ2ZtVx7uSjJD
UeDwmSaYOZQhEg4QN3w=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
b5TzJrebbTGq/pRucwAvmRYTRYSTXLJ31UHhj7qPdtWGaTRXaKbjtJHLK6r2fdEku+xRcQgb4iwR
VR2WDz2dfhkKseFS1Yxa2DFJTK597UszihjnkRHDocjQO3cUY+io6Cbq8kFDe4t/wEf721IVy63Z
z1z8RoAbpBZZGG1+seGG0kHDtkTe8wOMD9mRo2qsutfBPBsV5sK8/fmf9Y9E2sAlYwKjVvsGOjpr
dIS4pkfWNQ1UbQXn1WlPTe4wXcRDxSDWm2NMDLpVsB7PHxXe/ma6En4gcBeXFN40LqU3TWcyfbF4
Fgd267nviONJrvDRA6uaiECsHX40iXKsaxsGyQ==

`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
LoXyfjLEjXF6IqzWN8H3K7nR07wwyqyXVISYV16h6KsboFmbDcRTEPo0gH2rwN+AX6fpfnjiQCDi
qZVj+jq+3Jpyaex4T6xZDGqASKvTFZ53Vog5975jRBzfQilhyEnt1jyw4Z0UhtEM8LILdgabJqA8
cXdC2MS8KixvDgzWP6ABnTAwC9pDqbLUIqs+coqVvcy1nM4qt9WlS3/X4SHWNrmKgZ5d/HUtKouY
9yGUMGTi2nl4U+Zd7UaI2yJjVCW8JLst+BTCam4lPyVXo4ebpoEbDK6tTwa5DlOxI45b/ZooNuYE
Rpmlrdz/peCtaLTTS4+P11HF/WIAxGHuvcXpOg==

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
splRKPjEH+uTzvqD2tjFWmYXGYcB4TmcJH8LhGT8ueKKhMoa+orNkr7mpiSfxGo4nOfb4ddB5A74
rXupMEGR44uXFXmGFms0uV3Mo+LAVOswYWiSib2qqWdsJAVPQV+uS8kwf1pFIhgSfyhJYccE2+LN
qen4ppn5nmwPuAnPwhqNoxWgV6I1SCeKHMvOOim/bGhWBFyFuI4F9GeL1p+BC2DYSvijB6DHJgjd
lmuMd4WuXe78W//Vv2jhHriZx5nGgRFuRWE3VBR/38AWtMEOOrO4ijdAV2GyHZrphPmDHXfSwU6z
9JSFgLsD3Pd9zxwPDkqCeFOIFV991nTMDEBaMg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4032)
`protect data_block
McOR5osfN7FhwOeAmCNp5yxj8N3/g6Bq5Q5ouU3XTxl7+PasnExf0o4waiyX76zG70RaakRXMbol
AlUwSoxKhNyjkXCvIiWxYvaf7X84cSKo+JEKv/b5Rdm94q1QH/SQ7X9dRvORac1MTtDuCtBO+zBu
5zKvhrBmefLEYWiuiuOprr52zY8OMEGTbI/IwpCKXca57+WnR7nWC4FuVPbQ21m+6tXR4EzqRFsO
cqDqMu1Ab3ovVp3eqCWQitO6rEHDy04pCb1sKV8c0hiZzUHzt4I/g68EwPxa/XX8j+Fs3QgqC3Fs
8+ulEURPPs2r2ZSyn6904jQHnxL56kZS/iblOI4x6yQ1ciP6F+Va2qJG34pTrO2+umwjJpUU5hmW
LsQBb1R0fQrg0LtM0ngeP7JjVgoY5DPLYYIb7ClA9aX6RCdKNShQpPNTP+loGzH9uoXiIq8Qat7y
nKDTbjVHuhsNDudTYuvhv19rtdc3imoXRwdQnfSVBI7K2lBRBul2GnZFWgYhYFP9HB4IphnsU0fg
f4N92OMVfavI9rW5cK9MHLTjDRpFn5fnffpTwZ0oqRoJ6SwQ2Sbo9Mw66VDcBSFB0IkAbEVttWP8
Ew7KyPPIv7Rsrhi7gXuL+4fYA+o8oy8TtXUauSsAJk8gRzC1Z0YUosp26uv2Yw7p5hBx1yVJF2HV
DMKd+V4rqgBhNUMrJKVt5CmwAvUssDtyHWgYU2wZeQjToi3h4hSDd1A/wqrupXzihYHUQLr9Ugrk
KAGBmUVIibQLWSJO4JfypRlH5HxIsvmmAGjycOfh0wzd3B9EDH5gZAVvCp9fdf8pcJY2DmmF5Gvi
IV1wR2SZ91KO0kSiQBiNy4h6hw16w2CBIADVTAgHgU3UPgBsMTb0w5QOE6G1I/GntqXTySIcumi0
miNxaqrGdv9JeirHyOnIaBLjsehPCnq0h5LP6lnL7WzCa5XpuJWdLX6PuQjCluZIAj5lqVo6UXI+
sawtxM+pAB8CjfHjD/Jyjwt5bJveVQTXY6C/U4M8Qc18rmxFoNoeUb9cuAgog/tZ6TkAvjVJK4wp
M44SSLZfkpb3+VC789N8mklwDh2KsIW2gfm41E1uNApP+K048SvrQB2fyK4bYbOPbdrUNkFUKhT0
WGI+pNZbGGOvXkpGbzjs24NuKynVLG9aUnYs/3OZ3XPXxhXZhwkqig1JhZQ67SUksqLdwOmqAvNC
lbBWSOT7Z1plXe/H7RBjS2H1KjU01dhUfr6McHKLRBkUJWQLWge0UXkjT6xtCFUW35ri3ZRiLTQ5
FveWdaCZersd3LWdccyiDKQa256MBw4ZruZpPFbdKS1+crF9qH6mrXaL3T7VCeV5dQLy5LJtIA8l
dKRBxj7iKR5w05SRZ8VBmm9moHOG/Gz3Q3zER8414XEAIQpNrZEKICsk8BroS0HSNw4jt+e+7bwq
l9GQHHq1kVz/ZFp24x6yQORyP8Hd/Jo64BRAtFjQq9rF+DtFJjxhGsWnUkBrS4ER7Xnvj0Npkcc2
ClbCoRAqT1oMTTAEJzrRC8d03fgztYZWuF/t1L8aQeQOJGCzApSEp6PXOd9TtojP2u2uAL13l+rT
zZQsDx4Fwyphlm8euMIHjiN683sEcPln21+0pwyPMX1IfcM697hC56Q0GlEXHLmcgfF1U6kxZXuB
Qg67FIJ1tI04Sj3+IcldpvTCxWYd3yXNBghK43c6xsECkvGQ0adNYwkd7zRKSd7mgbzrsnF9zJF/
gQWAxd6lj+39h0fToKlzy5j7SMTP8ioL6EQTCO9u53X4e8EGXAciKQ+gB+U7et/nIrx4/SeEJAjE
ILPuyZQX250V7Ds3T8RpVEz9LRZI6iokIbR2s9G1837uM2j/+2Z1E8iZEA8vp7+5cFgIDm+SJ+DG
l9uuMmc2UkL7ogmO5EA7iTFBcI+CvHcbvZm4xMUGp6ZevdVzQ0WfvCSU6CHHxzvuJ/MjVLioO5wt
/7fQOeP1HSZTT9ZLLXlNThOUN6oL2Yhh94yiqWb0NV5LVh60oVEspG/Vweg9HELym6Gw7+cip3IA
mfCLiFrx6uifIVMZM2ot4H1FuH7zxEVXFDBq1LGlit5SNw8G79KpJPVJHMLWQz0+vL0BZIq2bJB7
96MU9akCIrltQhqZZNRltAjQBlYxmuUHHDqnIUoeFsmbDJvjb9RFD3hVjsNpjS8rqANz1JODRW3N
Zzqt4AbX3sS5B2UbYnJPA1IqIME5nBS+7ymbE4f27xhxGnNf085QmEYNxHPfmEWlhjJD9OA8aIwF
S6Yyg/V3Z3aiD/9ZK9t7JiT33x9tt1iDcmVCzAYPm2x7m8ejsYW3BYrg9lVjqTqX2WvkELPlLpk5
YC+bVpM7B8HFHAId4ZD/6IKkB4Pdwc/dPpskWy6xVTzRomvgLjNsI0i/sJsyXAvO3/bnOzpKklJb
BIt2/ZzEYg69726qokqMPRb8oc92lDwY/R82E9FQ4D2RS9uuCGcNQiuo+1ENPIEJDqjUgOVHUlAn
zh3AuBc0b5ADWAegcRyjKWBXGZCrMY/EMfy1HZdLk8UbDulcO5JHl0B84XxsU1QYKih0rVrA5uCL
aF1bGgsbcOYXIUahjDkrGKg1k7GlE7Tq7TV9Kx6tFBZDTgXOVzxSirAausVE20wIiroP2Ss9TgZ2
0t8Ov6zq+35t9fCOO59JyQ/vQLKL2lDwCWpq8ZFtALBAq7ghs81kqCWLmIAs9dW44QyC7ogopUHe
p5ttYELifTRauybnRDHvTEYuQoreo2ZE6vs5itp7px9TuIEFSTmF9hT/CpD+LnCkfgMBYzSukSwj
PUAy3OC9GzwOOEZvHprUUzbGDKI3H9K/3FZnbFPktrWMjlBc+8u23x+O/xLp8Tt7CL0kfIpshCzF
OiYnRosTPfDIvn7k1ePCEO81qp/6EuyMXfEKfEvlbyUPMEPvOyRR0yGrz5L3crhmE1pCCEZ/sxM5
bzS+kAJgVlGXRx1ymTtEWwVHlZ+KaMGIF+9er9WWB50YBOvG68Ud28jtw/HrArymVEAqxfFxcoeg
jqRjESDY5JNSpfcgMLm5c94xq31E0fSgBofcHZSutlzHcmI2U/7Tc85arkAOoMF2fSJFBqA+VRrl
lUvbLKA7LDHkKyKghcx18amJxhxxUsCN6PKpx+SM3e3DWT7aBSFIchoVr1fM2CpsJvCbp2nvnwUO
Ua4GV1mQVYdCHa+j7XI7hfAgHaxwIxtqbpSapANoF9rJR6S7Y3G/x3peeJWqgvdN5yWeNMIT+1iH
JoXbQvERUP4HE+hM7B+D4yVb4Vkl6Q5PljKo99dvgUT9Eu3vTCALY8MRn0B0ohEhMf1qteGoZ8o+
0wn6PpsieC96agWBj89asJVJ1X+rrhV9fATs4FqY0uAZRgnyW78VI4l/Nuse7Il42aKMnFmaIbQx
56mbV/LrFWKk67qHKSsFfHTZZRxIqzBhhcdgr8i5rY+W3TaZPprP/J5vqR2/3fBdzXuLhwoQSuPU
aDvp/FMEMyI+onya/xYmtfqDPDa7wCjHIiiQzwxWXZkALk0yg7WYtqiDcWoXMoy6xTqbJ0rL1sBT
P+Uxfc2XfqZUXeIhPX8aSBngz96pCLG0wMRcwdCS0BVHr77wNNfNzF19HMRL9NbpZT1AwHENYlWa
ZpiPNjc1lZ67lnmsRB2en8gnV7lY0mXIpSse0oTfwyNXY8y4ENxgmCAi6vVh43zvKz+GzqrGsSWL
nwrqwBvVhHb4LZ6tbOK9j8bHQbDeI7DcGlryhvZYhfW9Mju/T2xai3f82PL6BWkGjCeM4YXyB7Ih
5fbefL9h3j18d15W2AseoEmL8AY3gzJcL52wnUj7AO/mbgtC/FoiGuN1NtBixDS11lViMLsUMFTv
DHPWpwufFBYWflbuY1hyAGHU4CZ9qTVuKzk8PwqNWVHeI2YtzcDCYWkFILok+EoePZj5dnFk8vUk
1ZUsCSVvtpUsaKaZ9VT7wzp04XvKWQUQy6Lz7Ahy+YLa1Wwp4xhxpJLD1vsvB/CyVr34v5Y0lvtt
tpP1lTyywI+YG5dIChA10hAezCKZ6bvlm4Rld5Et0shvd5zED6xgxvXiLc+nSpS65UPf8YGdtlDP
EauT1p2sT3d9jz1b+N7gOgI96eoLLEy25q2NhoLf69VughJ2rqKesuEdI0rcR67YHmTrTiLAp07g
9apSsof1L87FgFYONBnsw6gzwnJxqTU9YqEFrp2YROnKfYkR8fT1ipwhT1ho0ND3pWKXkaIuigJs
JxW1RMgmhzJQFsYfx1aZNLpPc6CbrXZR64CkVrctRdz6TTyJgWsOFHBhk/D3PI5IlUCSnVfzJmKi
Bfqokc7rzBv9jBnmdZCfAaHbGHYU/6nL2jb84Bi10gTJ7ZOh/selN3i9FqgagYhafegpSd56F+Jf
6MUpfshgMyKx0nD+EmhVeuFLQ4xMIlPvL5DB9kXlr7Tb0ElY2UphHv58rgZnjus1IUzqeBjhwq2J
5qlQbEdRM/5ukq+q2WxtdpIv9vQac0x68m9Nq9h+1P93kFUrry8RfjqT2XSdoGh3cSL7ehQ+PEOD
ESIOE59ZVdLiUM2hTbZb7QEHQu/uuvHPwt5aXboJWgYleUGeWHMKCsCQQqICqHeqonMzf7CwVZAb
/G7zhiOVcoRQ3TReJu34hQ/ku4K+6bsCTjPqipNZYoNItBl2sO41Di2Wcus57D5ysVboljgcv6PU
ZgIXvxc804Htzxabke0oV12xVcAQUpebkXGBZYo0KBXIQBHNXIUcA3l3iUTvwNlnwQOt5NSV6Uhk
oaZWUlXSprRfRjhBW1Fi6WpMl53f/HyhjigJgx3T3koGZvFANLwshz6WyUaBNlBGsWqywWQDUpGj
iM30w8DWcu3oJ8ougFnKJ3QsEfctWOPO4gJ19eCStdiKDOpdusoxIEeUsAjEssHXRpvdn0HSfrRY
3IJd6N576qUW3qycOopn2ozfgXXu99mMEoGFbiD9BFKlqtXsN9Votw3qqLsnDWtJkcehlpaFrd6C
dRa6334xd/NClt7P1OQ9/sx3DDrxbKyES8ghtOfs8Fg5HN/KqQ8UAxG9kiK45l+iFaKvoYpyrENE
2l70wILQW79wBb7ypUAa5IhCx/wgtO5xYgbO34xC91Pba55BU3GCXlmE9PqKRHZCmdamOlPKxlt2
J2yqTvoBxSGw8KRRgZK1HwlJ1ym3kUS80FpVCQpAyJ5wLKCN79gnXNgNJKCnaeukdfQFGeAP5IG2
yD2gRPS7x2p3rVPNwp78TQmY4JjRdOFqBmbd9k4x21xZA2YdzhnT0EFCZQvupmIW311R9OWLNTcp
ROfM29FCRSTChwLvlADN2GRteZ25W1xpU6dQjtebnB0YvK9jSqv8mtTj
`protect end_protected
