../../../../../RTL/FGPU_definitions.vhd