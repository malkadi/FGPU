`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
pg2rOGd/KTcwDdRn8tBeCboOFrKztHkBJKehCtG5izAvyAC/6VXlCu46n5x8UdzZVRb9oGGVlYYE
EPLaBek/5Q==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
E3aUffY75oUaxWz5xbDFJvSgNJuxEb/vF60QmK+TVvXUT4kO905WjogNo/4uayw+RecdY/ITxnbm
CtBn9t8q14n4cGdAAdXMMc4+mG6cUPf9YQmOBKWmQbz/D8tQvTYba5pqTk+7rNV8R3tZbO3QIGv/
/GW2wfn4eyTXlNeJKuY=

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
qktdtfJMime75Ja10jhweJniLuEomGBQKIRjLt4/DHxBPd4f5v6IMUBc/AAL18Le+q0RBAZI2XYg
LBy71Pq6DU6GKIEvb1CXCPbf5Gc0vUcJsgT463ap+c8wSl5XhDplpCFHmg2AhwRj9uZLrBunpyOo
emofTHryL0pAPlGSCzo=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
DlreQrg6ErB/t+GCadQbLa/zqOHNaBgF+9roqR+06XbPb8dCiQL0ZSQRMJaGVi66waqEoPiqnGl6
EuEPEwu4o46cAQIw9XVZwnXzXl1hqYIMIEXVCCMDJP1gNZ36RbtWoNOfCJ+SsMlYUjyFhCfKRvEG
z+U/P26U2lsXBAOo0xSAptE/xxHpIEJ6r5Ggeyi/UljN5bOvkRvML0+aFDAxXqyKDB3MH512oQUt
HogVgoz8pIEnRD86bmxVcQ5KMsxicfY8HJ+BytWdvviOTqDPh01oEWKMAwUljKONAsRJjmczbNuU
+U160KK6tvUtKviO6HGRHyfZEjfNoCG8fsGLQg==

`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
fMaL/MA4P7FVFo8k5xbhVzAYHxt1F0VSt16y3t+grpO0DCKNxMad+MI6JoNXUNsnJMjjWvrnbp08
CXvzRQrrPuxA1P8Gn0GJQCTsc7aEeiqrU7RKAsUwphxuQ+dp1YBpo5kfyK2UJM9Rqem9InrflA8j
qCQn5gY6ibJJZK1kX3sQ3tqzfcC1gNskNbkkmPOxJ7Rh3ucQB3d7xXO6tECKoTPUNnDmKUotkcuT
28w7DbbZi9mKw8Rx7b1+i3ZLvOVbrjTEEpdBjIMRn+7NFO7OUeTeTa7zKL7/JZLs0JrQniolvYlt
zutGAXsg6zBHMCDdn5O/QSyGAkOuF9U7eOFFLQ==

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
pGCOkKBVsmzN/NTvFyge3xNTD6qIl8MVQ1M+wFxHHZ0wE9rXiIt9vwLlnfk4CT6zfmKxBzuyhMmE
jialmhLvhJjc/I9lSWrYlcBBAD+BK0cPWeV0UtGynTZQqk3P0Ja8Ah9PgcIypiXysNFbkuALV11h
fTeI1UyErbWB9F9qXj+7NgCJKZ5zwSDDqzH0TfIg5ykflzX3o34qK9uvuLdy3hh1kD/HB6mcUXcz
qc2hzC0ZBQKni3lkq8LIguAz5qVDTUyOhrEPKar/mgn4CGBEsjY9VT0QLHk3O0CPeKo4ydaEzf9p
XbLY52GkzGdXT3er2G5hU6HFgylStOK2fRoGnQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5872)
`protect data_block
0Ep/dM3ZqQUHqQzsv2G+GaBNMBl8+uZrOvr/WUx51RCRyVXOe1XMT808fCMU43VTbwpe9LcnvVvP
IqFYdpNWrNfpUfVLOd32oAqORn/hfEUTuQi9l9TZzToaymtwWAXw/ysyo8vHNC2yDpnPwddWaFlt
7fw5CKZn+E5HIRoiQFOlU29z7G9oPmC9nRd65o806kENKJMk+jDnCspupV5BCvOenmiueYxgB5cR
IgnfhFU5+kQGSGNMXl5A8HZSk3MboQ3Ti4TLT8rc9KzOnnYvb7JB0aI6hPtHrRjrDWA3fQElogRm
FFUgjE1f2z08KGxRk5RNV5IHnlP/+rrMluRmhXunRMCthzlX3eCjY9KXBtzKswJSRE/Bv4iHE2Hu
JAK3mQ/M5982H/w2i0kRr5noShkXfkZICQXcMAZf8TxtlgVJfOiOsvi42cZzaNAXoMtDQkLmwzr4
Q0AlpUsD4BnoxHTt95IMbtnrnNLug1Eh4crkqXAMCFG7OcEV0CpOzukH+7NQ3NoqyYDfGozXVIWN
XZhfEecxlW6pQuPHaITkYrPwGbx9FTCFLRc6er0TW6BOVuoHGsGZ7l/jeWTcq22vjzgGlFJMxpiL
SKBg/tRuNuyJQN8XL4Ki19GjdF62JHLnGHu73UFgClFZfA+5E84b/sU7CSe9QfGnkaqFzSEBF090
ZYH6JqUSuRdU5ZTLAOUjoA3fWt9I49zH0lDRd7IQ9gnMUzOg5d87BdeIQwvuQMc/LhXPZj4lM6ys
OvqXrPY7KoOjKPGt8QxsmG3xU43HtwupquQqTXr+sq4wuUO/3evxmPY8TCCKiVpaVCMxIAOyzHdW
xUEfii5CVoqh/tk976NdAcdISU0Cv2C9Zwfw+QFllmkxHFDGLauudjodVMatmJ5vlMlBRkgC2zzw
FMUHyrF1SGwF3pnpY7kHzDpmR19cKDrLmjXlJvSEfxoiS37LcLU1tqpWd15rbQLIM1O7SH7Py9Ab
+/XhohxkjL+B0QXhxgd2c8vGCZFpeGEzg2T25EKLlrDMw4I8EU3q36tP+RW7mtzLCmg4UQmgiDwQ
VpqPeT+GhY91up9q9xnqlOGE+wb3S1A3ENYgyeFFW8lKGWMrzPb73Sz2QviBQw1wfJsgAq2Xpb7k
kYfQK1Mj86H/F8SM6FbZMWevk9BpVSwz+H5nSCuMvIiRjTX1N1wsxMxudk9lm/g+h0H8YCOcgsAt
cQ4V2tljB7fuwbJvMIl1d8dj+M81l4WahSaIy/qSMJYuGTRr7hAuuXG/tZINigGrHlqSAGEAxvZA
MGVNKuBAbeak2i6fD4JZ4PEJ6z1C+dFrjc6ISJt7YRf73VqvOJHyLpADVnexOSQlEjDez6uxusVl
It0/t9kcNM2gzsrSSJCLjC3VFSyfFCGfPhKfDLMzJtKhiImlP3RH+NRkLC5q/yjORcNztxH6Sf1/
E7O3htAA9o0luwBTyomE0xX1iNAUPI3RxMGNN1hUtKzJCEZJ1JNhV3xQSAq0p35OrJg+Z/3c2fGd
wDHeOWD30ZIaX8ezjSwrB9VtTgXLxAnmz1AH9ZoEffmuJGK6KY762G6HkifKPqL9+FRXJ4Q4AXel
w0QfYHveg1Z5f2MOoUdjpRB54/7iqFHRYedLezYXonYRb3Xo2NAUnGmhmccgDWAxLRKAZYOpwez6
nRlVbGUcW7inm9e4el4ocGHUbXXlH0hsy+0m2i+46nuqcUqjn6PbuCtfN4SK+hmhaF+VfqgJFL6E
3LsN30q1lX1nKfvYw+oWzVp6wzhLaBIG6vweb5KnBg3SDL2OJsSNsX7R1GxEnlctawz6/hllJL6F
103ZZssYZj+pXwOCMFxOn0cQCYMqZfjYQ23eBB6/n/7qM6z2lmPGI+R1SvHG79tnsX7gkdywSSZ/
pgdr1UJomQ0hmPilYoBX9On3XxPglZZG+UfzEC6pA2zgA6blQEfrYeczM/io9mc0/9I9FWcaim89
t+B3M3hNmpRIYyyAAUpm6eRFyjUECAwVgIsMBezu0puZonkbZEVGOq0YsiDJ0ou/nEmAV1eSOWZE
LDraGsKsIAbl9rwoy8IF1UIBXmkCJuGQ21L15DL+izLnkRe3BsBAEk456BfqqwUMKKXgdVRWc0Y0
sqY7kFOlr/gSLFrIgFzgD2nKAte/9onoKxhBGNpXd+zm9xICrBXZYyWmzfUeM350tYNHdnWFHhex
JPyK7DqFpIx1kvBq+mt9ELUXVbsCcxP+xRcSUxXKqDig9OdAGolM+p2Q9W+rqQInwiCt0qGfq8VR
RZ80rQ/nQeeegpHD4yXlFDOI8FSlIfzFUBs4+obL8rBj0dsYFyk5guHekMUkNTo1bxUS0zSLXxpI
Lxhq+2lakbYUms1fTIH9/VSqr9y096lfqM+WDPF17hKaKZX9SyUHyFOmlXS0forAwGQkSuInLEkP
05OSleoVr/jR46WsfvA57o0zbLuN03+EnACfeJhcilNf6D05fdnKZoMhkwcsfYj6MtmlvUCqdYaL
tutQZ0KMUEcsobC62ul9cLxE94e5zbLdvQLAW8e8NnYRX8952HWNF/KDzJNq0YqgcLc2/52FpR4p
rXBO4V2Ycs8Kc7VbmynV6uCAa8OEXTBG101nkvJRDFzhwpmY0d35khhAmbzYtwwfDswhp14mggFt
s1iVjKsxYAwdSTNR6U94hyJJx+FSjLcEphLtbbtOKJRxFXTdjTauslSiXrJYS5zcJGW6M4ooKL2E
KBDLhiVfInQqS9t+81l5tO0cT+O6z/mskBkD6062I15O7xF81JAu5UodAs2H9m3PBAnxeXQBNmuM
KDsazxdnB7N9QTTZRAWUpESi11ZR33SX7jcSIxgS1gBqssJGZM3XmW7DVMxm7tFwhKoBAB6LvWa3
Sayzz9ogOPUwUh3990CZzj1KzmXRdscJycXUrKuL9OnNDw/zVfyEMWBRDBB7sCMMnEVxCyQZXwaJ
A8luLloMaCqrxrz/oLqPLJw2Z5oWJKXa8Fhau+ksQYPmw5rhDcCJHIjgxjtG7XYPUU2qT/5VIhng
6dITsHhVG+nZyuE9I2BnnxosRlxOy9QN1rzMmk4q7/cMezMq/FBDnygTd8nTTuPVONa8A4XwqxA6
xgZkbdBkBjx6I5cRd0HEpdPEcdZzg5OqjlQ9wfKa2ovyjAtPVWe9Zad10uAtidyr8BnaxTwBnAvb
Vuq5tjRoT18ktwa6aCAjWk1SjuiqZcJbIzPdTMM7/BEfHKm65pNTEdIiT1g1KiuAdiNBOdKnHgvB
C5sb+CNV+2CPBUyJuXQpSSVvdPgorMrd6rFbS/pdGfLnvm+PVgsN6zb1z/TnjDRtd7Cz3UCc5gDS
MBA8RVLe8leSLP5KQqAE3f8epP4uK0/KAPDUbP7rvhmNzjxxX8JGEMHmtDVOLBhhPYe9I7ABwJH1
BiCmylO9PE3mnnhAvoLhcET6RKLN2nuWDsTiZrkldi+ODWIJlxMekoVxucNyJ2kljyFRkqaDimIc
oLY8aQDEpybVw3iqInvTz1SembJhkdm2XQ+UyVGF8Tw8Qu1K1GendDrcJSYSINgT6l/FCdF46e1l
IZcYODeA9/CQ6eWb9O8NM2IbVec7J9nymNxsE7FoPtCiMCnhAa84iF9rLMQ6/8L5fJi45D9KONkV
5rR4zXkZlWeiKe4BVjK6xcGtelBRMU3Qdp9hfsL3un/U6hoEIRGbpC8qOJYwzBHnhZZlzaKYWHQA
7d+zzraMWVeyY6DwWM6aD9eoUYTIinF+rQd4cj7hi/yxQgRGHj2PdSuoSweOOQa/CLesF+oV7G5W
h2UWYoweOTFdMrp8w9BRu4Wrg1+oOXg1eYVdHFsZpRXikQajWrFa+o4jZPHrEvTfFhBXA78fTH4L
A3Y5el0FnasA4/v7TY2aVQlYl5g9BK1R4i6GNsjNhlGyup5G28onjGfgkZKSMjG7zKPEZ5FWsEad
YK0gg0mY9SdHXpe9otmkNtp8iOrhoPoYLGaxSykvbtZr6I4Rwm87nEIJl7dd2WcpxHZkRPwzD9Ky
gvEM345GIqp3oh0jwseks6rWDKvbnf+y97gb2GpTrW8NH+M9ZE9KdzUlWxsoCo3Qa65yPbBYkjOn
viOcRbZF2z6AymgdIE0IkluSHK4a2M4DIlPtC+40lIKUm8HdDHNHDR1LBjUk4qWNeQxOIr7yymh8
12p6xj+cuZTAv+gIZjrGN9yMfB9Ao82wOhLDjUjDOrnkQU9p+obI5kr4OBUeWe3QoXshKTXek+hR
9jaJ1eLOowyDBdXbrg/QRZBoUqgjyxsiylQyqCg0dxAGPa5cRD69yv2mZw/r0xgkvD5zcdr1EDVT
2x6HnVlp3wT4I3YGtIva0+3fdyezrdqRdxa8E3DkHIpYsMga803D6iWmayk2v8CWyxInCL+TKA27
PEtvCdDmrnjg1Fbk9iexGksQPDW4wlDTRCO/fHH0XuLYJZ8jKYDOb1zPdndMeb/RxV8iLPc8lqyN
9Ci8vSfXag8lreR1goPUC7nZ+0seuNeTZfLbO/sisSfO71Hvdy+y2KxPIhI0gxwrjP2/lJ4hW3n/
kwr+sYhpA1PddVC3keMHfF466ek6Jk2qppQme1Vqkvzc3Zgon9wfF5uPMRICe2/yslOud4QV6teT
omsGq5ksB5J3drVoPvqENYQ0AbLYMlrr5JmeZF3C0m0Rlta3/C+QQQc/RZPJ+1Gfp4VSpj61qWzW
oTR/+wlJHfzQsqRdOew+VsmIBsy9oUXOsJ8BmWFmjlbMLuC0wiO9MJkBPMK0yB88mwE3ndA9Hppj
JcmJ0aVrey47DqUW2tWAfgQYEok8X+dlNmF0tR7pkR0Pf21kJgqw+XpgRlkcwsjguCPp27OKcWrq
3lJliekGajes85crmVGBMpPt0mZ7oFqZAqLtp5J6YXHT79cQDer96MjUogh0UmV6Sur1Tl2kQdG4
L/vmcJynUHBBW3XgWnFQd4DM3ztvER/oReHNRvhhs+Ar0wxK/K5oG8tAaqVzfyu0izK8IVku1XrG
+pVVmbZuIeAwL7AswVLLjYhXvqNXyQpjoNtBh0Mb0YNpw1l83jO/JGTEkueSQY7FUXqoY8JX4Jqa
ui6YdZcRUVvSDAkC8t29YuvkXH81WMxLNu2/oWMR+76DewPSjNBs9PA2C8O0frbwLMo7jOhL1GsD
b4D41kvXY3KU9S7D4OCuSjW0Zzp2OjhHhVZF6jZZy4YzcrrpnGcqbmanZfauhxlifeyY/AbrzrRb
gVIsOCIF+LVTnr+b7M+1jappeuUZDEtKMrNZSuhPipLTLL/2Q0xSOS/fYYLX+QTTuCbVUiAyfUp6
oXi36L6XZ8+g7DcThoca+T3ykYl7N8bblD2aN3EaLCvPwsOf7j2UYfUP4ef/PNwXzLBqIP71zGrB
dsYT4Sb4qA9Oglqxjqdz8+Xv6yCD7wfyPANS7GwjP25w3lOvixzKaZS7aHDCP21XKmDl1hs9t2Or
j6JiRyk+S7PEIbGKAl9+oA6D6QQVv/v9XlKHIfqZrSzj8dXZ0yZ8kQkR1JnuaQsSABvon/KEGqdL
dAKWYplyQsDx8lak9752DDPN3uPLz5nbKFTto13Gi+Y8RBnUyOGtvGZlnhzjOAeU2XX8iijNVBRO
PaR/qNx1ibyDnaiFVCMMGaAcpwFhsCfvqgKNj57H6CBW//Ts/pBxR8Ic4QrvhhLHlx4YkbmbyL1W
3nBQzKY+5ipaMBfYNwt6SCsT606gSHR9OzxKpymRR3IBIHww19pCr3a4vpEfVI7ouLMxW4EKjAQ/
KDcKmgUiDimEsqOwH+GS6BLEGP+ILahTGn4m9U6lCZaQ9vVnS41d4IvCv48MJQ2W7O5Atk2OxSin
OeWTWO4rcIWLFO83Bn/6EP5gHqNbQ0ghBn7S2lh7O5FK8xUjudpJfHRw0j6dKtirPjCTz+zYwSjO
MK64lr3U2T+CABl0l0buVSSwuMjpGAU+2vy2fSNGDGSiG573rvNPIvkDOZggYjwPl4fGud/WQoAI
Ti1/SsoDqjWTasDgvuyQPJyHbmf59kuAP7Q8sc7ydajvVckHZwXFCu/NUYtKleacLoSqEszF3Gow
ZXmnGt0QRCv2M2r8AMMYg0MlkCyXDoNblc2exSOm27cJ5NoHfiIpWmLyESBKqU1rtCmZbUskXs0z
2q1XR6DgB3ELkP8BfTbKiZtifGkSq1L4L1nl/kmC04OE0ydJ95aAFHgKDb83tXOfcs22ad+Inkhi
65HEIPVCF66Sz9I/6mFoZiBSXAqz3SeUsm0xE0DPbLApIRrLGF5HtkrqF8yUlVQ4eDVTT/MIW7q4
bkPhkiVyFcHxPksbJfpXfCSLX34PrAirDqSMpASyTyVN4I2QkNAyPEZiOwbyXagKamUzEG2flKpD
sMOv+lwJ9SwvYtA9A4DfqFdNC89ujCF9pmA5UQL5GV5ISAeorOCJUIv+89ivCSyJKZb9vcZreBPI
EUpfULLySZDKHqm4r/4PQ08/92uIwRjFXPaFYSP1jBIvRakhyI8mMJw94pJVF4rpsv1jDjkguHLR
b/IgwGW/0Su84u/bPDK+cDAIjJHcBPzKtOsAeVEH+CFv6m4YEYombQGguLc660RgwbkBJqxQHR1T
jZq0MrK5Q5aCyd5Cuon2qBejqMemx+zQrpft3f6i2FfbW0nO2TRCGNu/fpCsYEofE4HvG8sQdLnW
7N3tmKfHvRa9+A2gLzedyWDs/3MEBxzMF/2cGwCBWaWfRFyoUjDCv9UrQ7B9oYa5bymHjQNsRt5p
TSQ0piyH6jAH2ZGvS0Cu9D8KdrHG9v9/J4HxmIbd7VuA5wpvU6zUR/FnBA9PSnopJDXJD430+4VY
9HV65nq54kVgML/MGBqYqcsXSC1VsKHcyRZYMbFAgiZJmRCEHHYRrgcRj4BTRbQMxr0tF5xB3uAB
HZ8QAUCujTzOPudrEVISzXjmCWoiyiK4yzht7NBlUM8VFzivSkgQl+vI5exfkPYDBhcUwJmauZdk
ippfi5ARXUC2ugbjpD/CZg4ivdEY8bnx5Q3eQyTJoGE4WvbQ0gYYb/YT5bm65q89fz15s8yb8LAa
XgE3v3E6npkv6wld6y87+E39wAM7Xyxgbh8bVZt06AIXTkDDtXqrhYB6EOs7tIFPUpV2O9ou53nm
OkkZZkxIXsIx2OuX3hyDQ6qYTNhni5hojJfTQRmmjKkxU+N92uFER7fuYmse8kV6ppHGlUM+cA6d
XenapeoMH2G6KNjYr1AsoGGeS7vPXQKxEoXrGkRy0C3/BtyYDBLO/AL/5iBLK+lOKEkPbMLN03dG
kfAa5/W7b9ucaOZSxcXJtSZjSrwkp7cNiSMrsCPzRq/PX90U2midsIdXJpygnS+9lwInuM3iqBoI
NOMgruCRoSqTHLYzr/YcMchyvgOwtVZLyKOTTB+HA6qLwXor3+2ppGo1T3pqX90W/dPTNy4jvBTQ
vEGibvr18xkytBJAQXBWDKFVApOz1FueEn6lN2T4qysC436FsORNz85ABDOf8+FHhe938IhSq98l
jOV+TIDNjMxpHaMhwVothaxzLoARXqMPJAQU6s/NnJA9M+eEVDXbePZ/fyRaIZYG0mFmLtk4TiaP
/2Hwqhvp0hlGSlVQWnXszP7yQAXtshkiGQM5qVju9Uciv5PiwHEPsZCKfXuePFrtVg55g0zYBHAZ
BcFwkL86XFJi3KQG0zP8y5VUH7v1aoKV8lai6U/w6ClwoaqYXVp+L3Iy4sz+CN+6b5pQ9GXRCwkV
7M2Vk0S1qz7N2xN8WtQaCPb5Ae1hAtVUKoFMIZj6k8D9PGFgwLdhK3xezfjBn+PWa6JOTdssharj
QQ==
`protect end_protected
