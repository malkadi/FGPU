../../../../../VHDL_Files/V3/CU.vhd