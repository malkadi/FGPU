../../../../../VHDL_Files/V3/init_alu_en_ram.vhd