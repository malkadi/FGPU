../../../../../RTL/FGPU_simulation_pkg.vhd