../../../../../RTL/float_units.vhd