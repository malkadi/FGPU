../../../../../VHDL_Files/V3/gmem_cntrl.vhd