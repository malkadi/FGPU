../../../../../RTL/gmem_cntrl.vhd