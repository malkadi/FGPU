`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
cQDd3XIPPlgRDhqULvYHvwCty2ZrVwzfefmANvx1dZIylIMC/SlAcj88wfYJOEUSOPC1U3p3rRJH
cF/G+RPdfg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
hcwXqOGXIKp1yMXglvtwKNDD2csTguI/218BbAfP1Qe5YaY7t7J14bh3PN4/sY8v5SUfs5PPhYYF
AVoQ7+Y8KyIAkFOjVjl8Q3cizlaMAyaX6UCc4wmflvCCOjy7mkT0VJKPELyiFH5OE1gTiKu4NfqY
cLpas2QiSAVn/xZw83g=

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
JJiSVarYWytdLFzHp3wkrD5+jxEb6zxCxwIxMuHES7X4vO/81ppoMZmSB67P59pBX5Chyu0EswKT
bCRha6XDZljqkcBWrrqj3cLRE57UCaEr1RVpDNBMw7hjNrwCb9eTELEwb3X0mZPKBqVrRNroBMN5
Mb9o7SPJ2GKhIDEDF5Q=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
x9rjekK3vn0E248BFQkRU8rm2REs1XV6NiMfscimCVnt3moe1QOgVJzTLPCcPYvThLcZJXwVyFUX
J1k2lVxuHKaC3FNNToKLX7girUcVANbS6jS2AjaAfdpYmQXF6epSjXy+KOWM7AfrGv2r7XNIcV6T
P4He3ZDDIABlWanBaDiVD6NYtB9SspFXaifjJ2faT9Et8gWmYJogYQ4BjXl960BUcxWS5faBudWm
MidcfsfVFpzH5bJ9L+thBkdIh/P3Rjr9ssCSzEagp+1l0DsZGX583KqMaKiaZiIsR+KyQ8Hrld0H
vh5k+kh3k9z7ewkJNwM0LCpa2Y0qGSJOxIauzg==

`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
bMGW+/GNxe7XIGxZQsPwYg9NhBUySelE4d3DawPwcsMkcAefxMJ1JdlslSvSp+VjxIobQhkauqfs
plGQEEjRkhr+3m8iz7uiwT6s+TtBZQ509t+m12KAHsziCshi0m7JEPgqnpkYUxS5ZbKQCRgudms0
J1TIIpIIdBJiHjiJWPFKhl2FSk46olekE0MQ/LvS36IE6UC8sP+H2MLZpAxpzqHuZ9TNFvVcyr9C
pc7viw1i7pElJF0USsLWRjDFrkLdXdznJwKPhjmDvq2WWhH0UZss4B7FZEDrUrjB/HO8EjVy2Hj1
fpw3eQ84VC/StEBHWhh2/ovbE1xsoAsXeBE8Tw==

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
pp8HZNaXt/evJqKzoiOa8A1cmkUh/1mQf/2Vkpam3N+hCoX7wAAqGU/zZVMPYP16RpMjeC5zeSin
YvUeVcdgv5x+e+joKUcjexTi2LwQorDqPIl0bCwYx4LccUexnWG6I9/pSM85Q6QNP03F3dTfZ+nY
q8I48HLVTNxhG5xD9+JTBp8D7rjXe9TJGi+hVikOsYhuY2PrwtvuAWhuicAfJnsIE23LJrp0i1cL
6oyVsfKsx+68L6qOWniySUGZ5yDe5zDF3WoQ1oHIZl8/tfnTJcGPsIRyeo3fpk/6/w5zWnz1pHuZ
HvGPaU9zIF3KNoE/3qKTDNhAcVbvP4+ohJfKxw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4784)
`protect data_block
nXe51dT9MNW1tnj96BZVcWp2ckUbi7OzZWOeu7JA4JZfny71Z/Ro9WFaR0keWyoYgodZ0HXcSq+l
A6/ETZ4V96mml7+ETYwNJ2+OyYRXXP2P8XaSeh65Fzo8b3Ft84w4c9rpqXlv/Kxnx4dGTLP5zQiD
zbLZfQHY5Q1wrVeiWpIvwOLFQVK2n0TOsBv+MdK2zhqKTcukuKtlyzCU92qQ0BMPZMPBdMJ1f6bt
wunfN0uX8sPBwWzgW1IyBtymXpnZ+YJ7txXQtuAKlk66+YE/49Vhp3bw2wgFj62F/yqXoVLqvgiG
E/xmWKyktNGAWht5JB88KHar7BY8prfsfZPsqaTkN4XmY/kYzO1NPfmcYexvUPRwTP5Ck7Rk8ZGw
tan4D3CNJfI/p5aA+WOLM2lpTpyQlJDzEraJA8+UmUA+aCjgNLdAXEzgF7zs4Jv/BEAPA/UhrNfY
71GiujCxm8gaVpc+6A8yLaclSKnxfRNQAx7e8BR4U+XuxFLAh6+RXBwRIXvzwrbXAgg2I14CQG0H
SlM3bjAWHSIm1VUa2m5OXqGk6IaIg57El5FwS9EJ2tlb1dWaCA32LcannUlWf529nWOHIsC7G54q
QC/QaKJVR+mgO3aqMolqYEOcBBNl5HBSqj/rWvqyOys1BbwY0/qoufgbV7TV5UsH3CcLobELHEG/
aN5YH+vn9UALNY4UFP+suwi/HHahKg+a4dRcjSB7JI0VRrHlzC1Ba5rvGJuAXiqusTxwEHkGuDCZ
11l2MUhX4HUjThFYEcfaN9HZ4geaxI8yJb1sBVsxKhgT+8tDiQKQk8f2sz5RgOmlRiSZ2j7j8OcO
7OuSUpCrY9QAQ66rL9cz20LMLLx8ainHlX0omQwehM06uT7b97pkp9kJYpiDRh6cuYPBWpyF3KFG
PWbA/EDbA5sWU4nBQYC1mynFGtwaOoCjnPGPj6eki2uve8Rq6KHMuCPsgDsl2E4BIoMF0nWPSaAS
0S8uYIP34GUh/4d36uJ5aKTEO0+yWayUDoOU4e8tMQReWzmQ7xmVVJfLaE2s7uuiTse0LFiGZwb9
2aC5mM1tp5JOS1XDtUlOqb0qY5wvm1PpgGCcUmeAfQ9Xawi4Vzbwny5udtMkYy1Pe4e2H7NGoVP7
KnADBiml2oFhENZYCXVBykKauJOqOqgY3iV2a4EVlX1X2Bl4QVDqivh6YJSHlEE9G1g31ow5dFP1
Iy/q6pmzNdlAPOCwl4ZT+nqtwDvxsJDKP5SvsF3kNgIuE40DfWeGlElNe3+hWJte0lv4zyCLZqdR
e4iU8jH7qxfeLJLOWUsQpr4Fl01WK3BdZl9hqXu9XTVZUcFOK6fDX7tbqNUjzRI+1MTQvHNL7zd2
7rM0ZmjgE7rb8tUQvo0iLTwgLFR4UqW7wuJ9m38KQwQYby4iF26TegKr5RWQYTZZ4m+h8Dj8NvZe
DoyAReXr1CVbPf+Qm2R4k/HM8EHaF6j2KV5Wv4GJERbhpz4h/g1h95YLToOyQMomALpJTOfmvq/g
7GbX5hprbK9h6eIuv4Lb0Z9znsCJJ9vUB8iPsSyRy0+vhS9/7W0xOgr3QtKOnYd8H8dIfJBi9EMv
Yo21oCXP8ZEHHfwFGDCCWKoP/9pe5q6vyKSqIE5gl3+tOjXwmTBWqj3X4BFD4rWq61RAdJZaC4pJ
EVO+cQ0IaJCvkv4jD6Xn1p3Tv5rWoe1sF36v/w9g7ZaqeT0jxIVoLXpBfgcHJYfUl4W04GM32/5i
QHsFnh8s7a563ZlnZIDi5YggZ8NLAqR9JRQw+uza3W/rrYS8gSd0K5y8T2LEAou0ekif08INgm9g
YCM9dXXiyecZ5Kbr46FSbMB7NW5rk2Z2QdIrdC+7tXEoQXc45nCX5yZe8ESbuOiXPzD3HwpitEkw
XUMcX8TQPUB132a8GuEsiGd1QjHitn9D3YWdwzSCDJ7SsmdDLPp9Hre9jnnryQ/N5gM45ugOT+4S
6iPpdybhZW5kfh3xC1k6ZekZ7peTE4s2t6zn2PaxGgybfnO/dzBxKJjsyBY+wAYcxMjmRZEfYKmQ
q/rfs28FVr8KPc0mwanN0RTd3xSUj8neaLAev7nvEvllQ/N7E1Lmung2aIH6H2kXikArP8jn14CV
s08PYpgUA6XdXIydplox1BB0pxv54Va5kazxLFWxRoZ17t1raDog5RhJryUEhrzWuiyGN0bVOWgi
n2vWsmywcsnq7WJwA6FpjSTvh+r2B/83Z+UQPZZH2StT79DyDhjYuJttmPjFTCvI5uYalwK6BqYD
pKWLFn8l1bWuuHR4gQ5xXyNJEs4vFteL0nVOuQlcEWhmDPu/YhwAxjoKg7T6aHdfrmyAChda58Er
GZR8pvl1G6N16eA/xyM0SrlFHm1siP587UlLXvDsXYFB1vvu08nRLsRZPCfZqHozFzSKySGT244H
cPEymALbxnF4hk0D9n6haZaAhtWDDMCYFDgZKI7bNkfiFBv4xjVuLnn4hRducfGPRjGKYICgGp0v
J5fEt3xBUyLU5xmIsOGBjTKQ4Z3kX/tQDtBME9yAfY+W+wqEEpfCNcPoO/l2leKgDBU31stLwJmP
OZY6LFlOrqQ6IjjEVGCgYVEss6Q0TBLP3r8Cj6PVXAcGVQtEaKUAeLLOMoSOUCXwnbWZe7WfT1RT
Ip7FH4b6l/XoKzrweiXCqP3v3eijyNmu/ec6fOxpoZV5czP4LPLga5O8SiSEdghvDIM80TQcvxKN
SutyDv4K75em7Sdm8gDr5BLwyOHVuKEw92E6hjoMbuSZHqfcM5GPAHi7oD1fHzwo3Ya9YGsbV6Y4
sNL6GNzUMBs0NQIRtrWLBJjbozM4D8HoKbZcqEPz9x7qr/sm03nLw9YWSkHHiPWHDAQbUO+lSu6M
AJsRZnH1Qof49hosV4isjrn8su/Q7IqtUV1H3M2VNLN6niMVe1OITFw0otPlR9vqFyoC2/KngtjJ
lMnOOzAJqfpjm2M1mk0ajpJ+eQLjyNhYXbzoMxyaXAJztqqYjqmQCqF7grJW+1G7Ic3vplqMdHbo
cx5ZHfPYJKgQNz2GyPsANGbETcBbIPTrTA0JIrRehCvuOW+5m7H0cJRp+PCmqo8TrOomeUXg8iSH
uGSlvLAMzP4GHcbcuRJeiGtTqrVFk8CsQod/ufqSZWrfaLBHicwCb+F/0UAHB4/ly5aG6BWcDhne
dGw5IaR7/b34PfR1x7FMnnehwT+qLSBrqW1JI21u7EakisS3cRgdWAqJsu6LWJer/Spiv7lmh63L
74L3MfuCIQ8vcHneHgPtYMoyy9Shuy/ogOkKGiXRWlYmFY6DDAZWVk3F9jQpKyMs04ii/iHKfw14
TfCEDpcaQd6ThAtm27DK0eSZMqtseN20TY6+S9BQy4npQSYer85G7M1WdklXwQ0gaKCtMduxCoMP
mEeexdUzy/mYJI1M2bd273I/3lT2lvNVXvHj/6mA84K9jgFH9RMiZJZ4Z/zzxsRNbohzu3/LWKfA
f9O1/oDde/QdxpY5aBWyREv41NiHNA2PE2Jaqy16Dxs1k1gexcJIno0CJ6b40NIL0IklK7XT8Kp4
wNq+K5fXp3ZtinXh5h3xJyVyl1VwI+WWfxLBOGwiC5rHCWWbmcsHt1h7IWT2Tznlveo+5SJu4/uh
mREBftrKQKq864vAZOc/L6AbvL7LwdkJfh+h8GJ85hyTBfOdscSMv3cUu5Z6OkpY4jYUp7D7k+56
GTZ8aDPG85q43U9WgHuCRxR0xF9MLgKZ6qsP4y39FW+9wCBcMwX3NXlZhddZDeWxNw5nIxkMRRJn
YbCiXZZKXWNOu84kh+Q7+ex+7NO0xGyUcPM8Yj1/9WCogbfWf1Zx2RC/ntczZxFdmwWURIaNEYwu
evG+LYj4sXw3+HR3XdHyyWF8Af6dNxiMNb0h6QrTMYyTJ2Q+ArLK3leJpoKPEaIDXTUzIt0vp8XK
FIaWrTWdUXkHzI8maeRcOSaMVzO6niuJoJZTgYTwYXJKMyXvuX1CR79pxIaDMKdlnS5Wi/npI1M/
uaSzU6wlAvv2APxO0dodo9SlKAPWA44iiXafeHMBtHMvC4MPFD3rYwV0pWHV12KuLGlfnmqo4Meu
KP+nbIaOtin8kYgCOAvG9aMVAh6tH6XO6sPaNLnWqQwJSsmTAsvYXYxRRWvBIcnKAWGB64t0BGkY
B7fHku/jth8a4U7vAzA32yMFQqWaraIOcgdC1DRTPFIFajbu5tiwtKayEO613tzd6+dzZl9pDKE4
lXTdo9ivBEjvDauX35jNnmWJcj4Jf1vZJWFoiEn9P4L41s8Dw9egXpj9vXQbIWzN/UFsclbwi6eW
ISYW5K8EbeOqoVgMmcdGeXTiWFoa2nb/xkrULWYzYVpuUBneKFPrfaqnT7I85DzliIvPwjBXHGQZ
ZoBPbwnj0iP1/g2qokTMT0cuoIBB7BHAXla+JzNpGhsd5cn/7afGPjy42f0lo7b63dHnzHQlftY6
dCL8ypn+BfhR58JnuDeRnBO6PJnO/APFCJb8v7x6iLIhPAMKdle5kiLIHMo5fRAPi3qIjLn4ssh7
hi4ZVnWjKRr1To63ZSZ9wym00pq79R3kXG0TIgJ3yqL6BzOXgvtVdESGFlXA9YJXcvdzc9iWxPV3
TizRbIuoKKrji7q7S9WcpYdSYz8w9KeY4TuozGXZDUMik5U91QlOXjhYF8dAN7nl/Fv/QeOPtzAE
xylzJ1XtPd2HB6Qucm97+NsAhwNbQIIX1gXbplvSwsh33hPVvTYNXYKm07vzIxHXj5bD0/Bq1SjM
8NN8zhPgPGkhUwY/CT3SeI5QnKN6VGSqdjHw9TOvLYu7SCu43N48CLLfSBb4yr0NXIbdur3N1FBX
f1DZ5JpQjgMtxMje/ySp5yQA2cBZcaGYROgqWCO48dKUj8/uClLQjDU2iSee8hNmn4WTBAqxcf+4
lWSc5wjYbNES/7Y9tvo2W1wIm/lrpPaic7HlrkqqVvzruik4Dd0xFgq6tlMvtOYRn2nmhmF+M6cJ
6/sP85fb9io1YZOzXRt9fNxVfR9u/Xctokhh5mWJL2mMFAG9EkiWovvAM3V/QEOpJOmMHYV6Vqr7
4kwD1ZL6y3wlHuQsecwAC6KSdlPGpbZyqK3IlJF65Whv6y2ngCqVlXUGTHprMGyCvbC1L5h7yIP6
k+mvmbPK+UtQb4pK7OxFz/umxSLQWTpdsCtnFa+uQGnVRmGTeRLEpp0lI7w1lD8jsBlZF1WVRC5l
PXj+3sDvnrX7CC0yrlrvOSRGa1xmvdvmWXs9hCfl22dIDGE5AUrxMQnei54fHxfRWW151Yv3b2ue
ikftF04MWjU7PrwiI3zmqjnrSD71T2IhRwG96MXniuNpGBv8PKG7OVwHcO9DcfRWpvSnWRA20HrL
5KjZKrsLSzQRnN8d+LtJj8Wj70yP8yl7tXyyc3Z+a6tUrLxZkzczyd2cNHG3N3Eibba7gKFfCHUa
QN46Z8b/3+pgEWlBJqDetyqNFNrnfayPQC8qRxuoUUWYJPr2EXHIxi0OdkCdF5BhjgW286Y5Q+Vg
WAQPFr5N9NrRWWtGfWi231ART/tyV9ZBgsvBGUelmiUD5wlGQAEivdD0nAKhBefZK5xDrrBUVxzM
umzD/yliG2XMGCKpUGWW5C7RKUHxQ2GwuGcqg3ol/tZPZxWRHhrmelm+cB416N7A3eRDJXW55AKU
soT2o/rPToH3URsUs1lfLo2sfuqJuTT6fw5IgDysyLKBmxmRzU5d1mjyRErzP8eN6ot1cFN7MLAS
dei0UwpfnfTyKo+J+SPPo2yaL0vNzfC/5DewHHIxCsjPEhVGEnYH0I++FnfVRYuQADTKq86tULQy
YAyhpfzbYNkA3c3sHx7v6+3Zlq+oH+DLTAjjiQoJWjGM31gVWDhjoWQ+pfvhzPc9Cnr1bqdZzOZD
1614W7+f6ghUX7FklzZo/wrFAmoChJrjvjNrZF2zFlYyBpemv1XProjV+xOdXwrVp/hWMv/Umb2b
DMgGxww52tJSaodfpva9p08ZXa4uCjeN9sf2r7Gie+odVsgm4gLD8y9SYFA+AbUtUV/JTQJqpXfe
u/y2M9Hu1CZWcKvzGAsSgk15mouvHsbJCFF5qRTMUr464Xr7UpdNkPIUHI20Xole5xh+G5fX/YkY
Wl/vvnn6EeyPuWYvWeUwukBLYfw0NE0MwGnZ7Tfn6+6e5oxgvA6AI3ql1+WFcc0UKjNeDzUyz5CS
37RyaNW1aW028X7RuKA+yR+LHoX6q7IFssXAMdWxg2/QFwU7rNsSsytCeaO+k9e798PCQOJt1Cw9
yLtwGuHoj7ut0owXErtQynVt6H086sHLQ3SuE5bX0kui3IY7ZSuiOtS3i+xuqS+vaqNFCbE=
`protect end_protected
