../../../../../VHDL_Files/V3/gmem_atomics.vhd