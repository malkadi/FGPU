../../../../../RTL/CU.vhd