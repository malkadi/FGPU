../../../../../RTL/init_alu_en_ram.vhd