`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
HZg7J1eicTLULECaPz6ctaw8y1kpWgApgtfn3Q+zYY0GMZZHrstjvvtt0rjShEIyHEmHswkTon9F
uInqopAFVg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
L2/HzTdtpI+DDWwQZLtw6a20VAniDvlrZ5k0iYB4G3h22Zth0ONh9GaVxdnh5RvsADtDStl24FLn
89acqSnMq2//5lAdWAp/jsSUiUTqUuq3s51XcviRecb87oOU+8iTczHYM6EqTAd3Utr3aKQ7HiMo
3WL0mQVpCBOpCQUD6jI=

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
OUJeS1bwtebGQThLvBFH3PwBsgx/p0nU2VJ+e9SC+Hrio/pbJwz4o2xpS2Z63xJ7QN7VhCBN12gu
ZFY5Ng2Sgl6wTkLeA9Vhfi5uJY35hY1D9sWB0j7MhUUJxRIFWIWs+H/FElpBvWn/H5UtcrDSuhP2
nLymA6ruYrGfx7a8Iq4=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
AkdqgHhBI+1kEGsbiaO9eH2SWpUOBQkGBwaPxgDJYtBsJdOF2T3rxHzMH8aRRo4rOV4wq7F5qDYZ
2bRKyZlKyXwxOIrgHQ/aFSyCdbfrrJedXNOvayf3bMLKWGvmkeKTZFG4ie8bYq1NlzxjEK5tXh5u
do6EoDDl64fqmvjtPSKx4xrYKjkfDGC1J+lF3Ws5x3iNXrNkIqRirBHfL2nwSIIbCGtaZ+SRJZcG
6fOBaI5sglgjVMndkM1UDvQGQg1m7SekmV1gNbuTjfVG4yDcoHwJCq9TChQTCfG05c2xR2kyrVm4
vPlYfKMD9L7sptBiihT7k+285Lhb3gyxkn+LZA==

`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
kU/KxTFv88aIggtPFaqaw71mguuPJV+CvKI8SqHLyiEfFwnEl2rRaQjfKPPKVY+a9ar3+m1VrJZq
XyAytb5FrHwHwKJ8PWa7bc9KeMqYCg0WQyqVAR20oTRysvr0JW9ZU5xcZQIfn1WQOAidCGjGERXk
D8J1Mok2babDuVuQ1k1BLyAGty6ATMVk3dUAR5LIplcmY2dcgXHhvtTjcDGgu02ufeeeQgDtYdEr
XxPaZ/IuZu3RKlqS+LyaN7GLtQ1sl1FVJL4oxiYEefZ24cov5R/2KmrDI47bvcitqcxarcKhbIwt
EegxbadS43xqD9JDNFUAaaCu542z6SRuS0zC4g==

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
k6DApHKykfoAVe03+cLJSaTvIyV2mgyg0ee9r8sDTCqvO5kwFuomMl0B0cjUO/4j7+8GeD0YVUGW
M2t6DJMbIxuNlNctJRXzSjxwlBu2lOTLqWCd5V9OOHutCH8JEU8ndSXTE8ecj8B3ICDoE/uYntN5
p9eeS5YN3Awwuuf7vpsiQrcsy5iqvO8GW2b0InrBhe5m2bb+CK00dsnS6RTA0bU4RH+b9zcISWyN
JJFEeDryWX5A5kyBX+Em8sHpW9ssoOlBZUuAR6sGhqbdC9endcp3vkYasFpW89RPhQcAE2DOJVLu
qXK6y8bpxJSgUq7bdln2TJUwnHb0mgJEbAKlHg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 114672)
`protect data_block
b6F/qiQzl30/hekDCqOp579uiF5hd01/VS8ZycjN4pZrZ1CvLjWYG4jiNmL2+ysgQhB4w7jI4kTb
g4vuyOENhEbrKwVN1P8c6gPiCyO4nAkJiVYQNzxHe88JtN0UKyp2EdkuHzHzT6d1kFZc4gOi5j/h
0WD2dlkVRhoPxDk7OXjKmjgmcAW0dnQ7zbQJK9VgtQUOybyF0Tdqv2DbbiRPHa05tzER1013tfHC
qC0IFhe1xBQ1/H9Xuw+fjSmKSj+gv73WuJeL3p7c86GLkJiQqI1i/FX4UI2nIsm+yGZvQKOGEkuh
dgZmZJ00CsRDsuz+Zx1MaaotSyJX515hD4IMndWoG6hYKO/8qxVxOramP15ni5atC+OIMxnsn1c+
lcyH1OaCCBZbbedOFzujGKhX3SeKgOe5S0vJ9j5Rcj4eQ7rEg0UY9RMePkPGP0bD91lMhmopiHjR
heafQwoOjqanHYBDdzneLEWaMU8Jm6rJGzRcXYP6nWt7jwhYEbc9MtsoMhFd5nH+BprbDeEU0zcI
CAOm/K9S3Cc9JyzXZbfg6yUZgAK3ZtODQx4PQMykEftR1Xpw6hD+bL6EiGiKpcBHxlO7UiKOmOyB
urUtbaFde8NvIibKkI6ZxU4OiONq0pYrhEMeR871T040euXvnUPfZjco/+0RbhLNWseEoi/xY1Z8
o9T8+QVPTPOIXU3g24Whx+cFcwkda1n75kzn+s9oC3PlbMMZvVRSBDtIC29KSXmH+7Y9IH3by/DT
LWkgbSFmI4rcseHl8uzINnKReJlwLapJ8JvJenRA26OQlIXjzukbxn+JyJL0MuihXI8YfJZyq/Y+
IqVQWDGxyHvsEIICPsq6h75gfAhUCE/IJf6UAHr3AIg6tFHgeBubE75Kp54hagVR79u7Wl0bszC5
rXyziYJtcCmTfF8e3b4033tnaBtoO/iU52pud+l8Uui3zd+OnHEiW0eiOdCRhvYTyTIIFYnVzCTB
jpJ3sH6McErapEBgE54v3omKrT/5PQ7O0E5DwbOnGgjOSLNo7oT+OOeOG2n5lhgbZikNbXxPDt+I
kCIO1Eu6MkTj144hQDEgGNvedgMc2eiGnhU9D4RQufwJC9w1FhYz4HP3zC3iXZN/OyBcEIi172Y+
NBLIe7Mp8f+Ad71ShMkSCa5qavfkpDN7E7ZFLwS+HXG6/3I2FA+CShPppctLmb3hseKYdEdVd9n5
fIKawwoDZnWWjLX0VloWqzsuOI7GDKvxQdee1gbNx7lBUNXbRxFLcE9RnXADUF8kPo7VV5lwPH9W
rxwDsV59F6aRVWBivXTlsODxxi2YQRE/PtXWjtl4HT4EJ+BUOIyQjExjcM45lc2gFL2RVGSIOeBh
TbKKj5BBhmY+CsyV6W2SKsq152c8lkfkXnixdmsLWbP6m1itnPthki0RfOrY9zTmfpzqlIVpOIqF
P2ZWEkPUNPrVOY5WJh9dw6kiKlgXTe4uUC+VrkCUDz1rls8vflovKMauk8Uoib5H8n0eHtDiUIjy
Rb5ltrWawGZMS1f7ZKCDMYwA0yb306mFUJwk69sZMsnONXw8nJsMo/SDDHZTATcGH2/eVNIi6CWR
vZTDkrOLA85b3vZwh2Z3Dk8PFD7/D/aIH1wdaszzQ2gyhe+dXvl+N3j0KGK1l8H2kmHFCOqbObDJ
p6PKSgs+CZu2Amiv1cZaQ7GRNzCzoIoG3zWWp+uFtJFT9j3VrOwZMkNc9b71rHdZq6s8Gon4J4oG
skPPjF0hpw5RtXocAQ9D9xPrlKmcsZYbVwAUSAOy1xiBhE5B7b8KyCoyL3W3qp4k3SJtpWPqENAY
QClbNYSWdNTNFViv3OVrtUoo7G3VvNTv/HroiubNe4S2vnQBJbxIVrcnbp8XqmoRdBVm5Mg47rjH
AdIJrMxa463N73dmrh4fdl5/gbHVPXUItopAi3p2NujKJpJPKf1uJrgJDIJS0gAPgAU1ZX7ECgv2
Zw/oVdP6ez6Lf6V1wEe3OQbh4x0qHsB22NJ0qlVqW7lqr/dnMXbde0V9lsPGxsfWzZsuseZalh0o
nI7DIrdk2EOWN8Be7giV6S3pubQe3Urqy+1+6OkquE/2zlqZe6b4gEPJ3sKrel+zlAlABUW3IdRA
VDX2uGCEgDI6P0a7YVMMNms5pwL10qTMgMswhEZeaR39K2JaiHclOza8iMTxf39/9dYiVDDWuG7M
4XlLtpoBOPjy9gqZiADfgONEFvlYRAZutu493U3O8oAx5RhZpJfNbhttw8kblr2JDWOXf83P6rzB
jTENJKXHYTtI0JNwn1mVPfcr5SM5Q1CtzyQsASQ/gHhmC5QUjAfzvXoBV2KhdwAFVbPQJYpLR/RU
4zo+g/ydijB/7k/bIErgNN4lYTA82S9wpf0LBshVRedaMfMehDJOYy1B3X3+Hl1GSUzsK8lKZILB
CSRGzIAtQBOFJ5JT3njf86qRWcy6WmxsZRL7kelWdkQp0y4VP9gsrX/9bSOD5B72YDvdHjGu3gp2
AXF0mBzhEDxFKiAvjlv+E/G77qmYxt/hewWJDk1xovoN1GPsWSDB/HVvNJeoD9WCwKjyMgn6SIaX
epwUh8P5hMml86igahvEfNMpE/b49BjtXZ2LfzCyNWQR7XV4l2jZpwP4K/M47NNrZ9lKJIG6w2cE
lXL1DrK9ylYeZngzi9JbQOhqkc1BlHKD2iFn2O4tqZCXo+QVEfVX1hE49R+YnVIA/ymePj7DJNxX
XVuPOCAydmMsEo4DbGHoHxMZQ3QFKRSdkk9FKlCsmSPpcakY7MEIJFOoiYq0B4O/VrXfbR+bgmOs
nCN3Lz7sPstaQJ//I8o8K1Lw+yPYpYSocpjYoAgQp6yD4ikwTEVwZdeA22BT0M+EZrhXlRaj+kPE
BKHGJOWTBzl/8ffvGonXzWZfDmLmvR2DpsVgkhyjhKfbfiU56SSjuWN5hCQdKojtfL2HpOmx0S7e
rvUHW9GsYg6CqCmDDcJ9erlhzFo1F1qViqqAbXLNyfmvQiTFONvU8bU/JCftslX/QuloLt44Ac70
iXJuH9NhbjHA6XIqc6zkuD/QvU59eUx40LusPYgY90LnAR5fSvLM+eNpr6ehccNW9BlwmCJ9QHrW
x3tWB16Ic9SS261rBVbR3HzniX28TcpIwqcOoJKSbLNv73paCcNT73g/n8zwuzboyUAqRR50bQIl
8l60RDTAHw5asx/Xd9wxyUHDNFy/ifMszAXfHQvTviv1FKcaw5OFX4fCPWj/i9S2t2uwpiXRG6R3
ARCcgBNHiTuO1MI7qa3h48EVKRVNa/MLUrW73TmWMzHDgN7EYaP1HkdeFgb1pGBYm2To3GrXUz1V
J79ohYIbIVjJKYL3aXqrGekxlKCBfeWneBEll8nFMLhlpahdR3hdvLTtTImb7FY2aHttcbT92arJ
Pjx3tbm9SRMCRP9B/nf3Cwjev8NnSiekUrW8g8wmNnv9Wm+NfAcEVB88t87GFoft3lQNyq7wa8lO
GSgXF+mU03y7+fDhsaKDY6/kH1zUE0WRC/JNohP3asLvDUA/uO33eA8LVichM1owO65KWcrasZSq
+lt7Rm0t22bFcR2eEtUiAJm760WtayvrXfms05hfhHTyMPPgUzEPR8uA0INEL/xDq6Ium4yOFgn/
2ZlEE1WKJOX2vFPBkIiqEvHURuG/GH9j05orzOLznaRqrCK2xRnMLqGlU+lJHZofqe3yOdS0AfRf
eb27rJ1vz4reOa6HxLieOaJlVY62+fsBfxuEH8Xc2i8McV4fliyRFVRqf5AANiwvmJX7gR+kkMeO
MDzcJQQ4NHPH/btw4tG4qsbLbojd5ENNyc795bUFIyGslIyf3EF18s/eeuXbvN4OiljcjqUcD097
/xcSoBK/+BDNloMf7lfiNyveBN3MNLYAnubzskmElTAXZn4OcQUAIK12LcPiq+mOUmnPzrbgyW30
ARWcoc74DOT7MQHDrgWb8wmQF6FjOLyqSfVsCugPTSzup/OE2GIOX3XtxDwX1FmEgxE1W48cs1ny
XioCZJRA6HY8aZo25QdWZwTxfS5gu4jedbXJNeAqzxDLMsBsn7qLX81ojWhjw6sFRsdniA85nzkz
dUlWQPASVTJ8sQx2+FzF2DN+FS4VXrsjuCWsGSE0dPbv5hAvS5kuZXS4E1YnZMKL4sMJWa/vDcKv
dO9QNcd4AsZSPYbAc2Vtaq3CRAHZhwKs2xsMkJEC92DjiMkllpXvwyudJSQ1UV4WKvwiqUuxoJ/I
HsEc5d7X/jGALAwDsDDswtVlqfQPW7lZ29tj1882/ICUIDiPmqtmioWq4r+nAhBn2slUpCy4OJie
9Z/q8LrnC7utwhN9IEI5jfIcCffYtnsuqgjwYNZYqe/erwotHTbCwW238i68OhQBXAcAP0nfUpL8
EmQtINDnFen3qKU0Ljsp+NZzqjqyWxNYXH3cd0YbNvdESdTP+9k6e+9J/yPV2zC+FJTuqOm3M/2A
j+OBxm/0fSoYhvxBVeCW/6iWaNokprpemzF1DVNiigbFwY/2Ja0Vgf5BoqH3gc8Pk9SDT5MtT7hm
MTQlHj2VOvy7/ICknRikDgiMC89oBkjZSOfvbsjZXshvFnshY7iXLA8auFvVfxzFWMOKch1DQ/ur
VUXvWkMV8IV1UX98dEYRffOcRy+i2bxCAtdcUkIbOQFLI7y4oZnc3CwgiRlTGgdbJBA/w8emwEXH
yjcmfAKUU83PmCOzoLHqRJSp5wlXBOvO52wQOzMQkSIKG1uQUWxAUSbtFblqetfDqRPm19X0oKG0
Dwm6lcq9G9RkP52eLhHyZrm5i08Gm1D43l/vwmn55YlvtLUPqAIs+pdggDm1/WkX7r+pIhPjV/GR
ZCY034fN46+DeAjj777DPb4nv4vpzkjG21wdQ0GFTUqFMOmfi8a5tOPcmrQRbOqw3Xv/QqUWHyX9
NCKtznbkIJ8MHTepu+4xZsZ8VrDiDG+nNSRYunGv+CRxUo55KE+CPfx0icxm6GAc3UnhHWT3YCS3
tdwMn83uL00ncvwmDkRQPZvtW57ib1DfUaI+FU3ve1YZRAztnv+LL0q92Xxtm9uBD5S0s2VujTQK
jUinCl/jtaFBJVC7Xt8SySKse+upMV4uDlL6+JjKawDQ3hqiXk35SWG9A5qpHA0Z3gYYdGYkXoKb
b24Td/Kv+WjSdnwr+EhkxJ7VUPHZ+oT0ujJ5ZBLoA1PKU8c7QjbYrkcZpO09yWdJS9ilRqoykpt0
yRVrwNWbW1kt4x7IELmPssvn+GLDPZryFjqgy+fxFZaaLoywBnwhV/QHJ6XUguXOJtp2RzP9gFbI
fLGZeRQTHIfxQa9EClBq6BckwNZThHpMbjHrhQvoYBM4hxcCVaP3MOlT07m8GRmsxJmjTjYmdd4l
+nVKijaGNXZnfZkGykH2EpUQiFqwgr9Pi/uy72v5sRnsbS8N3rxzRU6kK8T1OC+WcY5mVzqAmOTD
pmFHiJ86QovRKQpba1DoOWwpVbNdL+J47PM4p4W9/prL9AHBZ4HwUzJitLRzfd1s/6Z22tHzoyoO
eBD2vN/sdDFZb5RmfvdpecaseKx/gsy7HuMiH6fdBgfHKWZdwYrv/DBjSFr0aQbFXsOuSvKytMBx
IbyukFzPx/KifJr2i8sk6eHeT8GbTQ7+xUaB5q+Aml1VOPip/EClw92hRzC2Rm8GtT4aQOCKVJ8W
JFuJD24VY4GOocR7+uE3tXhmxou543T6WLPHMZegYOJ5Q7/ozH33L4R2kKIzMuW72MzfywgrjFMP
0nOyjay38DVAGRF0fPyC/oGYAlJfrrU6mfpMtTt1h8D/2vdbVxWQNpFSqEe3BRsN+ndIt7B3nlz5
j1hoMpJmEW4q91cdXLfYjJJSyJwH5v4P2zc61zccD03AV+cp/asof/tkFi56ro/MX/RzcVwaFTia
VEixNC8FTfJ+Zr3SJ734xfH5vvsR/vDG1xnmy5Z3Dg0EFwkehTYJfxhE8lb7YTKs1qQjyOCSonkf
bkqKCSp9ZeTGJrFs6UeCdwkfBjJ2rExmsMCbyckqQfEZ4pi0DMowbpUDsok+pVNyqZ9i5Nh4Z7cK
hHblbO8VuNZAjoYro9RN+Nbjg4AGMXL0k2OAwFjjzOPlUkkE1c0zMsA+p0AubXbKQF0pGrKX+W8m
2b4ho2nSr3rwELksLlmz7SgUhXAJncrpowU3+H8vOBsrfO/josEFMdf8v+JyMG/WMHt4xSV1tCP/
VbTPapRRL1MNJBpemWxWOaKUd2Epta10PmjT7WmHu1Nom0fBTFsTTjM0H6rdFH3K4vP3eP/Wh0eA
3n9ZuLpqa7TbKE4VeDtV+t+LmflBdjPufZn1VKXRTLzUKFZkh8DJD9Lc2jkdiPfRiudtsVqaDsh1
mDEPdsnvyNhw9lZY3jbRD1Z7wGFjQPtgTaPB5ijmDdP+6O8d/O69RcPsZo44NXviQm+GqAJYwZKF
c9qY4bb3KYjNVQtCWpiL7cs4/j2fthfeqmS+H+iEvjai6h4d5QB4lJQ3PFwQKJfmUDMJo9goZK7u
efgYb+aELlPVlvob8lbXLADDEYquuHpKdSFzsXCE9pe0SvXEnTa/29+GORTAB6Dxzrj99S3vgYm+
FOHdObaRFxJzow/vjaXsoSOWE6Uk/IXJ+5wDvFxFiNykZnYrcVAn7MzAIb7EoqrXBsNGu1hnfZnH
CG9uTM1eFSANr0+7rbZg4x62bPWzWj1H0/9/4VJ+KBF6UszTYI6BRh0xmwNKZCrOndwKc3VxA1eD
Z3jeU0U5UHkEtbSgMe4ahcilveYhQoBl9sIhLt8KXQ8d0UXQp3t3nayhhNH3YatsZc89Gyhi4kly
jwE4vq0hn53/I+IUjocsZ5g/dZwuU8kJVTbcqzH2wo5y0P0A7r/a1iWGAM8bbRnK5CcuVrmlGaCW
qyI3FGBf5qOWibWeXho6UyJTJxjs8Uv8HgjVYYmQpf6oVWrTZ6Re72xFiDN82yc33hSTiUxEXxh1
ziqUahTP7V1iQbj4glbCXCT5Kjs4f5CX4dzZx2szj72o3U48YAZoan9lSmZp8hSsguit/OUkcXxA
AK+ntS2W/dCaNJcpIcm8rWAIs40JAH+oLJOgn/k7VkexIoShMioGyiwgYdIoq32smXCQ17i60eyH
8khYY/kqli3jS0GCeKS8Dqjj75nBkoe7slalGjVNurKgzU3NhoYR6pSqCiXgSiAk4B0wAbJqYHVk
wsTpneeEqDcQPT1lpfe6XCfGRlwhYoh3o/ZqN29nNo6wWpCHQEdHah3LZCLJyn+ZaKyXfiDbqEEU
NvS65xpcsukIBAEKMQXrFzIUuaizIO1e4OsvMS3/3NHbaNoUaZK3jSDYsFMFJcShun+8X3UXEMuU
My9901BL9yhYJsu64PB/g0mRVz5ctumPl4We7djhGKIFvcR9HgAYy2og/aZDpeI1BLfKbJ6e8RCt
ydHkeqrB0vgog3/Sk12gsOLgfr36I4dqEuY2rxK5mu24PPXf/jyn2MyVEV3IDL0WZK2ErmRvGZ5N
GEzGhsgvx33H4LgrJtGCl+Y/+KkMAHD3UEyEJPULmM8aNhYDR11n1jxZpsRfy69KmvJsXivLZlfn
uKh9HNUohIsCSM/2+Kvq9HnrqqNJdmjtRQ+N3Cmvw3JQBHEfSNwvqlu2dP+mlkBgqVVBFeYXSFCC
T3olI6OdWJRTNxQclwd0ewINMCSjFbb6KypO1F1PfGfnl6t12dR/BuKkI+kfFwM++L52Ci4tfYYE
7HgyGtkSE31OWKp1u3c6l99qHdOE7WSKPz3Pu/AYWsiX+sO6PfD+g4sdjezdhYuVVLAn/0iVyNT7
7854tEVm13go0ctXvwtIpqEoXfaF5cBHCyXpTrmMlWqh90+u2IRCD2VJETDt2Sf8c9tEagr7Rh8/
0GiSWfqmPwmfRgyrf4B5F1R4Xo1443gBQyCYxgXF7u4eVlg3pkwSHA9A6mLs4uBZ8VWLQ6AmlGUm
XBG1W+hbsLp0NoR8A0cSB44IeXWC2De5mqrOCaRAIZmfKO92VCaz6jmVcWPQIQGPS3dsc+XJlGJ8
8PQiJldzdRLy3xJkrfXFzWDdulSmMpIATOFydAoGAwR5JwdpZg5RoQyMUJ88J4aX0iHj5GFWSYJ1
guZttfra+HmdMPQaSJVBnGeg24bFLUaxVZVIp7MH+ii4cOTkrMzYToHpfpSuai76QREPWqae3amh
rY3kq/RP9YzusG1Q8pjgvgiriiTxHCyFHVQsMIhtZbLl9K8lAxU1vdgnVNkVi5Ss7/n3Ye8wOy0U
mKlUyBkrQTtN4XCEr2K4qBVyq2EG8WzOFK1rov4vYHnkTGe3WgPkj2OHqyeIubXiCDk53iR1yo9K
W60aSHq2YuudMLXtqrZx1gtYvO03pWAmFSj/xwz05/C3N7wg8MQa3095hC9pHKSp3oYCIaMiYmZN
zcD7aPQQWaqOSeox1G9VY0zJBNsvY6Phq2Y+mA7PLY55Aal5NU91jT2NPULvEVgjuQffRzXs4qbj
AjBVTR/QJ6sag5ThdJ0nRXQDBxQJiQdtGS59SRxWF6Z6fkGaEqTwik3uTZ/L+RUeCye8T+G6OMmm
oDPR9W78UykbAgXEAmf9cIacLc9Bwytr9SXc4faBlbQZUecpnNtfzo6zLfuG3KKqQP8LIxbekE7C
K6BlskVSDJSzdQ8zW4TBtezb9x5o2JbZyACvF8JVM7pr2QtaoPrs4Q+jDeB0W1VxsILFWc7gtU5x
UuxNYipn2/WKFZHY6AY2KwGN+6czKp2FE6NxqDSK+RO3H9LpsRrYAzre8ZgbXWlgQ/1/HHgM7XJf
PHvGZZSSA0+nrdfMj4ISXunCVuqwP3p3wMUyNpqOcd50ay3GOGZEXcbdJ/bkaHny8vqSlHlaKSKI
sbvUo/3w/Vrw5P7CRG87N1nHJet68OBCxynJGkrCxl9tvCd5A/kJFZxral+hQ4mJgLZkUoG3aIpJ
v8EBPntUKvkykASDsWTPed8p9svjQSym5ieTPPTZ2N4lvuI6k+5kWtQqYt2CLqwwWHMf+p+qIuqJ
FU4kTaO9MRODd0e3gYtpMZEcSappCuQR/iDkvX/hrbneA45vvJN5ZBvTc/GHjoMROWYy99zTmGnB
KTBMI9nqD06v51lRPbE1c+VR8y08zIvtGRMMlu68tAgVNHJ3/oVVPit6JZ3a/ssTWIKEKwX9CQAJ
C1SdmUrYcvi52B1WhhINEhf318Mz7O5wmkRTbmjp0UrnnEAWbr+unOJVBD3oy2EMEVOGM6hAr8Ej
KgJV47GvKIlr2kyvcv04Aw0Z+0heEa+gzExSkcN4PUOjsMK9WtqFSV+hJidvI5dBcNn1OOvpwB/8
XfUoWhksQ7dpgbBXLmR/hWbldyERP4aeibDLxQGQMJP3gDjPeK50oL3PCY3F9iKmTU5gAyDYezci
jYOoT7cGRr8pGugvYEtfLa1fx2Oc/j+qy2Fj37q5Hqg5ZY1KYVLNj7jSbSpSyZ85MACg7goMeTQt
mtWNpYdjbc4cp2RgSlSXyQRbuBT9TwXvdxkWmZMuRMU0hYJ0EhoUse/n3bt1rlkMMaQN5zQy+UDe
FWpoMYOy4kOo+rRjzMy0X0ixFElLGqqODfmXFFtY3aW6OVwZn4DQhuCu+y+miu26BdvhMaSX4MzE
ajj/f1/yFSAHjUH1MAzRrydDzWBl8GZPpTk1zn9W0LWsnyNC9nbsTPKjhjZPeEoykFHnNk+CJzT5
vo3a1dslXmWxiMRnJiVgmdYSzFls/vKAhTn2ZJ8I9CUFAq1fwww2CghAjLlFa5h0XnR4pFSG9xi0
zd18+CU1zaIw6LAFcX11szP8R+fR+8EVU89v+0BvoLyda3I9aHCIcTNXT6b8KKKPrr3z11XCdLul
Vg3MjHXhZ0uvKcrrWVnamUk5ueK0Mn1AkEzwZy3ZqT/9y8Fd+j0gUaJyArTYsi+voooNFWdlbDQP
UxWjB8+Q7dzLMdCJgKPBNj5T4+LYdregp2qa9HfLKhhwpb9LGzbYcLJBKeAYiGIm/U0Tch2POlz/
ZI4zhElC5MAB6doVvA0EPILaQtpg2tQ6JNP+7U3DsJxZKTaOAks12Kjv0Q1rSUTUNTyQZboI9/Gc
Wb8bhpu0ENSw313envW9gKZMPvjW+n502jrqIYlOrlB44pTm0ErATjzH7aR8plg4HJxQ+OjGfoPa
orilzf8CFKGM71h+7hXueF6mBJiEHEkQaUd4iFjYw8LepYuLsKW3WgOaUoE43N0iIb3xyOSp6p6W
9NzDshVIfDPwFWbqiIXC608MuZh7/D7XZIrpqzDSCqQ/vLYImRwhVoTD5jRjcTal2H1x2R4/2+us
cWYIdZ6ZLXhLC6HJIN27hj3se7cKo7BI6besDshUVOXK7nLuaP0hx2zzJixIeZtXLIwnJ4snGdio
ntpccfCopQzENRUQBZp1U6VngD8JIxsbF5FJ7EfipEuYmIVbKrMXtGCJjT3Dy0ZeszPtffPSablE
Mo75Fgnjn5Iit3SIockDHAy3EAUZjfUfVNVQL7WTC6IEpaOOrgV74DYxbZf9EO4BqpBvGvpLLfOt
dJ9X0nL3GOOdb+0DS7XbjJTlj7gLkSp0L9DuhE8wD8mUNYx/aqrcR7/Qw3Z5P2LpBUZfzcK5IP3h
TuDZr0PrdygRIzmxFo20wm9dl0v3hu8vj01JhKFh6jTYKLFi/P3j0XBhhv0COgENmfEbj7pIo/2C
1vj2LMVGdhXXNNvjkJiSlGbla3+DWwUqrqZvVHUkL12Vn/sCW4MgnCbN9x+5sajqhzT9A7idR7LG
iE+fg1NDUsDcsnPZgYfBvsA0FPG2OU8iAsZ9OR1O8p8vTj5Bv+T3+KJ5FENfOHmf+lTtwO9+tXjL
RdX4PmLwn/9bGzLXS2iCxTGqLZXBQL692PKLGLtJKNX+okBVtEkvpSxK9Bi2N9QkAHD8ej5S3sK6
d8PPeExRfEOQzihkVQMSUke86J43cJbXiAiroiil9LwQoGTshGBSZEizuwNHBKRMZ9t4Klvtf6Vp
uVbST617UpF50tqAsepsdcP1fy4NSxoxzDTvX/EhKjt/A2Nj8wsoDygk5iKqrElEHznP3RGAY1ZN
2zMBrHV0XaKgSzsR/0H2BpXGV1GY7sId/XhNAMYGcDwaO21LthDHVC/jLVuHm1Z0V//dE5mW5BcX
dYtCVqTXw/vGpu+rgWC+JIo7RSAxhBWHiNE2ByZc65YHM07zwfpnmGREsP5SqQQJxD+NB89tIaTO
8fjq4jQ2CO277lbSPQeJpCboTJTmrH5b4f6XYGhNOPvrNBNH8sub0GElG2f1GuTAf6MI7YdyHtRu
KgeqS1KcA+vlf4qLEH1bvlyDeSAGgmLg9C9y7/ukm1IEbN0O3TsigBLYIhn22X71Wi17LunYn7R8
UF+u1cqnOV5ZMBIYcCIzCXwqOkL73VCN0T9S/kgfRvOvmr3+65OfEDrgB+c8CYtHqUAcgDqbvmey
NN1HUb1pd5D2Y26ALFnJjKveX8aEmaurwxp7Ni6k7+kV3f6/WEp4Jqv9xvZlJrcRQWyWaz+WngMG
r/oU5ades5V9gTnmHVj096O57ESt0lnPjKKnFqzjiIG/ZmgJQR9ianVf/5nziqh8ksDed87+alXf
DRAxA1ua766TblDpLdb7sd7HfkT4KT7Bnr3nhWz3WPWPXKgi8yoE7vkpXQaUnMuHnodbajyff2CF
Gem0xk+ztqq/8j1KUkpWXuFAuVnrCxVfmA2GIIJ/ay4wHYhuMSGlyrnJh38afq4Uh1mAiTDjmpVQ
aEHMgufX2GDtVGN1T1E5xoGJFlE7ld8mM45Gxp6FhpQYOt6HF1bc/bw+K1/HMjdNQsdfCjeHoAK/
PUbZLLtVhG62Ic4r2elvs2yF9zDZ11MzFta2Wq/TN5aUPYTm17zsbaNSOQ088hSyT7ZD4o4crfAH
/Wa6qFXwpM5vPTfpnUByGQFAYjY+du/S0WpQS1oD7Ppi5oUR9A+I1Cn90XLS0pWVXuOcLRScq6nI
4wFNQry/QJEeC9oVhMc31EohOtscRo4dbDWR2gE9TEpkBR2qkWyySdSZKQZD9QPqXmJdwC5nYQpo
P6j9bjNv77YeUpcyJdWXJwamoVfBY7U+f3xmj4i18S+hB1Ki8iVElMR4Sk0WMTfo5aPvEXQn+iiS
fnYGEBjclbSaGv57Ur1k/LOWcTUv59JjQhYFURBpZ+aunYPij8jqvWCZ8E7Gy1Gm9duK5I2EZcss
DZES8QcdJNTR6bl5uAL783cfREQj4TrWgf8EKxHn/dvBtR05XCsZSu0IOTvrmBROFgl+yrXW6iCM
3RDffBJGRKeaG9AAlgP7VOdOrV8tsSwP/Sop79cBTP2fVo59V4a9efcq1a3u8IbdIw9BRa3SE4nr
GQKqz3CaACuz+GBVoivM2iu8iw6YhtM3mJNzbufFdG4/xRVXiPLsIK0LaXg5jHKIxknP7nlvJFrK
RvVRlICiyLhTho2lm7k/y7kjCAcQdf5hWOJXArjvKVF9kEwTY1abTN0Rh1ZlaT7qSc0V7Ej0xQ7o
QU2lbeHUMEKV9vy2l2rq6uLevy64uLwL0LnHNwWsLaDp6OmGZHkkXnFK9RpXslmkeguntOALi7W4
zncD7rJU+tx9MzTGqjL+kYSlI4nZlh3y0+J53bSanr2aoY/xKu5211OlfoqINBLdxdLV130CjpX9
fY6pvHl020TdhltwezvDHQlSr8duLOiSMPERuh8han80Wfk/BjG91HSAYeErekSJaGZQYO/Gymz+
0xHR3DT3kcrqsHw6rWJn5O0+fibHJN9OwwJ9B5IRgQWjhjyWqKlWvkyZvDm1FMoZOhypYSROh8jk
UXoiYqx1lQjr/97laqTSx3nYwsxnIwlvy0M/0fq99Gldn/mZICwlUC4vDIKoV/jhBP8uQXdm8KHK
7mUNfsSBTLmuO3QWgWU9DuZJPdZ8fVRs1sbVHfukswDFjfTNi73dGiHeQkNdu6DWzrVX42wLIyDq
EI3yoh4KQca+O4one6BUJcplp7eQkiobf7pFHn/Aa/tbL2YWeuu63b3QTTnn31PIScFXYzxpHB88
OWXxphIqLGLoM+maKBI6s+sIYKTmEbVCYNhzSGGmop+ei73RXiguPkd9ypnGb4wO+n5cjFAk4v+F
aZv4AewaBYtNh4BMtKkxI1xyEmK6HIjRft1ezOdwv6p2WuinIaqctYbADsiB3ZL8n2jgwnf8JOTY
pbrqH9lmKB5q4cCxUYWXrnw9tEKaIJjLRXmxYNrida7tBoOQnR05L2NF1i3u57WykwZSIySUoR3h
LF7XZANuZxJ0s2yNMMRYLZxgXLOLz+elGv/mYIgtG36TnAyX+T8ogGKEV9sVCTNH+Rsv0lOxdsek
KbOd8iVWely6AZZE7yvDxAIwnJLYBz5QjZiR6xrk8UTVSKYcJAWLTbaunBA+NlPGnfFhDyCzVTiZ
3ZdlQZzXUK2bR5H8OF98Hu/LHy5bY3u7L6sUHG7QmLYWjpPrSEhf1o3QPGTWvAdUt0hFmxesJGwk
0PDSzynaV+LarnmWc6qs3DXwWwD8nqHODj3FvdMuN6uAW+dd9bob/Ieg+dgPewvzKM5Ygiuckd0/
vkDCk14sFusPKquONprezsT7F4ZKl9RI7f/AdFO+r/J35GtQudgnf4bdEadrPYJam5ZuUuuAvZVD
X00vHTLltJFGM8EizZi5K+a4swE3IoxfzvCmlG9BB4h/ozbzKHfFZmRgM4jvObXxm+z+Ie3V9ZCk
UmfFeyMOWhdQmPHO4/3XhfcF0PRhgXVvMXGORf4097S8pUD+ILN9NUGMXfZsA2sFMP+gGRf87TPh
04xnFQINCBfRy7q8gevegWvNVV5r19NtmviEaajWYYD4iNI996S/79SpEeqDShlVuabMsKGqpAFk
nzG5ZU8kmKR9x093AKiCH5AWpkDhETRz2IaDeHGAIRvzNFg16MqEqqIR0UgzmjH7NVxb54+c6Ral
gUOIndetPPA69cp/1JETpjqZYxL6FVgICfkW9mmH0st67lk0evCfA612j+PEL8pfXQ1usvHFNDyu
nSUUs+RHRazAxfmBo83dFF7EUk3FQrt9ZSJRlGHqWjRQVO1YxLC22KvevcA1PtjHhB7VAwAyNYnE
qOwqCFt88JxNve3g3sMglUJUguyv/7k3KhCwMGxIL7sGAdMnu2pvYiOssQ9mUzUK20VDQ16tapQm
HbjVv0F78cbFtQyHPLgX6WPpN1NVrJm8hhJoKe0yRcY5K7cGdRNXMphqra55aA1IObClifHPUF/v
UEVTgWM1oLRDd8q7oUl3nHOL60WSFlb6j9mymRPYIhQnlVlml6bhSkagtYq+jW3ASBlP2/UO2V/O
h6niXOlfDTEHL8r4C2EimIcuhGGcqyy7EZwRO4UEwMNTkW4v1JiS+i5UPcXhLHIvZKGe50YIhoOA
GiQkPDnCjQLl5VZr5eT4W6bDkUT/VPBy+M87UHqdqPXzNyJ4arBK1T1Ggcu+4p0SE/3GsIthiNjS
d5o2baSaJ75/O3Qjtu7uF30G6STe2ZdF2x3VU4ilrBbXxqioB9A66rbNv9T4EIpbavdus9Bavxqj
SBPzPHy6BlMqT6vaGqB1QBYPJWjLPrM1cg38RT2Bfh0pueNo/QzmLldUiDII3o0EF5Aob9NW1J82
DID7ZdUxfticCOf5IdErcev5nsLuHERAFNy85NWcLGu0juoG0YxvHYPIoVshpXnYnQQMVux0I3Sn
6iD2SlOkqHORV7KYXpi40cGwwlMggdCav6VhQ027POkZ5kT6KcxgDvl/IiBSaGA1/QvgiC5Y+qAe
5IgoYrNWMEgHlZ2jfZjOPAw7W/WwQhOOBh9EH2JExPYJV5EdSWjvHgPrABtPZLBuUF6a0ZCnVteB
2hBo4CVHKfZyZqe/ufNBnbZmXA72YmBY1/hOv3rVGHuYvCcKdeFFKStL8My8coHy1WnTLDhG6X1q
qspjddwtinW/WmxhQZgo5YkTHOOm6fscAs75rGCeSX5oBp/1rYrwE1otrMfayod5K0qXf6E8a/Pg
KlXaE21hkbIylPrASDz32NRgHFlfSc+2WbhuMCrEacIbLQuftqJaTi5V/WwE4zxIptfb3pJxDUPi
F6nzRLgZkJPseq3hRyZLUVbjeGIyQ3YdWRw3VjbOFRiaNR/y3x4fo2LaShIut0T5Bray3xLka8Wt
RLeAszIxLkaEy9JiFiyu4pjvv7GD8FCNml6xZyydhar4NRG6JmsIv3jFgHSJGApN4J9IHM+eN5Rw
XPprDeAvHYjxvw70qDhz1U4jb270jvqSkSe1PwueanR3WIecBFhALzrD8i1GfOVoAf0faySk3d6N
pH38t4YLlV6UKQwylA8S62Cqw6ZZpuu6uEZzgWGhcBPSuj08XHC0g280VrnOkK8gmFl+KmyH0f8F
I6NLa2uDcksA9AJUX7l6ralfVCZk0ACHCPeZ4Lkc967mgdIjub3qtTVq9lp3LDLDK18wqfcPfBz5
xpAsEXqa/t9+ZelAwfvZ6DXxoT1Lkkfz42pcuocHrq6idCWDlbOZ5hKkU+9GD5B+Vy2ucYCUAR8f
lraIKpFUiCSTN7bhSaGd90eSM+xsha8teQALVoFafwlQ1t6fPWXTyy4Wxbp9o+XFt+XkVg1O+DV2
pIrQlRWiG9rvY8WtUMcGwp3uiYWlONenQoPyrOGwTwHRZSsCj8uA1MOtpWGNEBTF0/e15jJ1Imn+
9WXx7e0xOSfs9aueoZv4lI2BCP9FZUTbR5bVeDhX9ThjH0cOBd/hT2ubUVKcLjKBCHkx+Ei8dbpa
nzc4m9SitkoyLb/uu5A+Ha5vlln3J7vxT/Xoq31XN54037FWrbPvTeGdboEjwHPLe1cWjpUAvGNV
AojGgIy9rQUQQrnXrcAic1NLbVIgZJ/U5M3LGwR+33Q8wMsVBS5JcFUyQn2Pfot+OA+gWwo/fEoS
7KeXu4hZCeVdQd3SCwewFhF0MAJuOvtu3AE0JU0nf2i35Gfsg7RPYnxlGS3OYij++JFgC6KF3b0D
a7K1hiXf5xRmgUtkDoO0D0BZQljlVqUyJYqk1cQTT0X0IBdmexUBNAXhNoJGC0v6I3Uhp99EE7cB
YSdaut/rmyaAvdgfXYcbTGA8q7TpFK0HnosOUP47SKbz03zLIJweO/jQAKfSVQaWKHrQT0irWnBd
w8zM/tmDO4TIQTRxbMJGogZ2w5iqLRcdLBAjpv8QjKkjqcdPW0bpkcuzLOXZzi58drrZw5D++f4H
anSyiUajol898wx3KZg4mXBRncsiuQsRMs2AO8MjbWqUhDlkFSlZcayrcoxiXSvwPpXWvV/UPjya
TxO8KvQr87GJDG8c1NO8W/GrnPkbLMbpKoNglRzIRuHsOK9EqR7V1BgUif/4hZrYaRH81hEnmPT/
NvJALenmceQPZ5Ln1Qk9dDMXOr5A81+Dclu45dcEzn15GXxJCh4Jy33gxUyDaJ3FK1xXPAYXyF/n
3O9tBADEtk3o97wERMtGFg9uZXXhmCXvEe8CeKXP7w4k1n/pyL0uBewDaEgl/bAilfvbAticQkrS
fd2RE/xSNIVoO/at/ru7THLXA6QeZVPLUKVRz+Lz7NwMNQ5l5S37oaAMdb5r9+Nzy1bONI/scbUB
OkevxfRNrbtTWTbslBUDWd3q2aO4GkA4Zslk5WkfomDvNhu9t7UcvKyOEPjf+5kV78rdVHykxoxf
Oakp/ZI8nF944nxkYSQbuW7dcEYVYdaqnE5NKjK8nuNN/nqprnFIuQfxVzjRZxac8RVT0Nbww+Qb
Ti3IoErPcSHXi79xWqxgrh4CVpp/GtRnmNnvfQXazrywg2+CHZseVifSu6piDbWB1WbaSexznlyi
DjsGatzGrSZjgqfr2/02qRACPyiaT7cWwHcXMIbI8DgcLIDbzgKZNNAhLAvh48ZnPeNyyIp/sRIX
Zu1okBWh/WxTREbU2vxrIOdTy/BeUQhSwI2XTN9kK+diHo9T6g83OlBcx3vCecSzrqOTpG1hde25
xHFmF+YSj7pEoDSbWLJbjpip0+D8z+DB7R8RJEJ7lGulyaoQJQol9JttXzOC5jy9LrlJkgKNret+
q7kqb6FieBaa381RroY2PyEjD5sLzOafT6YCHWhPRnC00RT0TNqMpjThk7TmUpXlirwIZfNryvw2
TUGzKm74yFGQs3XI0Runh3Csr6x2rRI0Kb8D1vSJ5fIOe7qQwEpD14+XG361rTuHV1Ck9CXqsxHM
7+sZaUt/Ox3NA/dMRwEnH4vXIv74Vkh/tVd+tBCcVhrjJK79W0v7K0OSOirxZKu+dtOTZUPhycbL
sB4CaQwQoSJOlfXVVmUjgQpCI3aYfrvI5AIIAfdnmcauhRqBLT7txOoPsQK+K2rOie5Bp0jW2jst
sEqQzKN4Z+yr+Ju/gclwHZij1XrGWyqJRIp1MEVjUGQciJSXKQrRZ3eZSvelL09S1wjdYFJrOXsQ
I6LUMIw/l9pVfT5aYvT0+sX6g3lDZJ2iW/EXpVRBvyiJTS2scVGmHF1Eh19dm3ongPMNmPZmTSEH
z1AKC7vYrsdd31tod8ZDYLFKGIaDVOyc1Qh5+gn1dj/RZidUrWwdRCZoABWcRgmw5FQ4NGk+61J9
41DOyWrcJdF0HS8NRRi2Ae5GO+8u2gM2CVkTZ/cvEvywxFoy7I94E6LRujK247mqx46UMoJHYYEL
ASDxk2UdP95GqNv6vUB2RwI1ryLVYvOaTmiK7LRAGLGYaFfLDnKmyX9Ol5QDpfBOJ1DCSDkiAV7J
h/Chi2BQOdLaML4vaJl+NKOfxP981+DACsncbbWyuo7ie+evNqXwMjuwE7wNHC9mfuEjUi84AmNr
W73LIf5sZshNY6N+SO4G+3+D10KpX2YUsQnwb46+3swdqBfDb97oXo/WjMyyT9NeO3G8c/dhY6h5
z/12nwUk/X77CCIMEfJvrtrzfsH73IlASbFm0HYvhuzf9tq2mkK2uqQM8vGW1bPI+GZG0ALAJAJG
B2HPftrsF7dA/tu3fbFq0q3WM1WpdS/V/nc17TRWMkImdbPrHbfibBzH++lv7k5QvZwXI26/8n6D
IzHnP0icymSmMOWkQieTnAa377mHT4QfslCboThV3wWsT8i7fAsWg4QMl0kDpaPfRUvGBf8LFwvC
MiauW/xBlxYeGW3I4ob7Ck10/EmGtbLW6VwjdmW7r0BD704O0AbLQ8X9pFn/xC7RdNbn5RcAkcwr
F+muUkoB9xyCEGnJE94WU3hZRtCa9KksvHWNm0KWFvov1u+HGMYLn4+QHuSlGf8kCfP41OcFPY1L
GCjWj++f9SmBHbs+dTy5Grc9Fa+PaerYK9EQAP0pO/06Ti/8oIsq5loL08vPqLYyt8o12yD+WhGi
SXwQIMHRdVR6gV4dulUubjmQj6uh9kks6sIS0SPiwgxMsploaBlWCJ9yTM/8/IInHEhczRHtvAwg
T3/kmunoWjW5wuQB7jHiq5In6EY8ZGlhScndkZpj5fZSqX3xds37IY82ErcKYc5aaQDF9kmITBPk
tWqbmBDn1zyI1N0fP+cB83go/UsWv+W1UUuGdNsMHTGkMpgEr/HGZi3RuMwV5tX6E4cGyv+w96hn
vzMAhcVdZ/cYmIRbge7j3llTt+p/OMa+/14ufHLazifkT4JS9DZ6+H0txeXRhA98aOYQwWfOtetT
Bm3nHH1Q9gmA6VcSGMSIOoXuigH+RCpkqfvfm9qY3QGpz/ZSWeUcC/ihWkP0OAfNAWqWimzXXL9A
d07SuwzA8ncrF4XXRmnd2OnO3oh9rXKbleYyFL5ev1R3co7aSua7Aqy/IpV42+MXVjnKnstOlXZN
sPci7GXHZYU0uCq50AjbMiamqkd0y+C/gihMrrr4WkvjRytLWou2PrTlUYGOf8seROXHPhsj2sEI
V+UE8dX7urDSlbTHnXLJVDMd7ZKT63tjtyNZtYNZXuakdpHBY/kVw4N7QtmEvSka6bkZU++Q459Z
df5Mc7xrGuY7UM5r+k3nh/wtN3wvhpREB7MxTkkCTd0d/Yk1/bgUiExmPlmBQYZ7Dz5NLKD28PR6
4p7HyhYP/IQRqKoi66VFVZcZ/twW1wpPCcVGghQI524yKw6pNzrqWIly6BPBK22cqzzDkUstvwk8
MOGWfBbjh3Jms0DpEPLQsQ+p6qp8P5vultcwKDScJzOWME9jeZ+H42IE+z2TVZAQ3Sq8DVy6mbKQ
gyAOWsP4SFZM++V9BV244n36qxHXUcIXkGOOL7uh/GYQe7bSBHZ/bHSDgUb622VLE81FkpNMaWqk
8QxyFiIGGudlhsxJeINrP1ekdglabSFV5s4qs/6eEr49V2PoH+Z8A7k2GiidbkqLVZ/5ZWQUG3xI
N+Mw5/Wr/m9xEQ5uQXLc+W6yDTcoqNkZU8Fx2gg0ZYvzIejSVpWfi+rVJCNVVsrC7SQhpApeigdI
ueyMT2czK8L/MPBgFYT9GV2B5W5Rgsx4eHHtvFexYnumQ7/41xKSgkbaXfFVcvX15C1j7976fKy3
5NRc1iPxc/KMkHdydq5nQygmRSIXoIVUYB5r78o0VIkJ62oqkQ+3m8PVUZKV/WsXXQbUxpoMrhyn
bvnnS6xb7T/MVI5F4TAE77KMIYHecgcw6huw5sGPHGbY1pepc5/Ahn43LCLhBQPwskZlLx4UY9pg
35LIn0/gyM4CtKQxxou/zNDlNEFM7ZI1HV52V2JBhHIhDyChCaIjfOwgfsF+ngN47Yk3oG+W/ljX
V3mm1CmRh/RsOB0o6gWbS9jqMqcA6bTDK3qFndywfBqV/78GKEtgJFtlsikcTNF1X/OUpyMTRmzO
/iGwTFSLEspikcrrySKiX3+muatBI0JSvslOcP7KZRkPnAgvuGLMvB7SkIoZLobLjv73vZEOh3qg
xOKgnHNg4ZxSDjhnSm7RhCzSywixrcx2r6ONNBGJ9rWNu9AU/Auy+Pmv2JQIQmEEpTh43glKYE2o
uCDHC9kNWbW/zbWc0FMg8vDpVhkeMIGXwXqk2rsb69QJq0HbTS3UkVBdyg7ZrS6gLvXqeQLC638D
mIw64b9FgDzqj6YusG4CCDL3IeNYAZzkprxpvSzQk8luSBqCfqsp+Lfj55Vs8xCTx0fuwx7IiGmC
13l++toVFPboIo37JUMohEX/vrw5qBzRS1WI5A+NPU+vLcFR/M8D7lSi+7wdPq8P9E6hShOROti7
7vWoAweBNJbkj9QXlfV1aETVOtBCAQf+WiOf7lK6aZR2B5+miBCqv39wxugGC17LJ5SVtXCe4343
bJG6zFlPWFcUdWDdguSusdTcsfkES8+glNZdGJS2/bJFtYQz+7MYi81tObZlH+bNa7zqf41Bfy2l
8/Xpy/SzNHyDyF8uqmusJh8VNj/MbgLbIMuGEG/1AEOComAT7p0c3n2YiQD+u5WvYZ7fWhIJ3W3m
O8nzD+E6IR6wJy2fHcpkDN9WuHoCejRIsLptLFfORrGB2rzr7GhLJr51yAOUZb4LHM5V1CQ67Oa4
p9bwBrsU5BAw8KKsR91m9VU2hAFX/PUZ8W75YtTCcG2junatTzxiTik6gndfcCaZ3HJCKmsuV7K1
YHdy7264mQ8iWeBBUC3z4Cl+eALsL7sDUeskBy1mXYxf+ykq0NwRHzqwrENNwcg7oRMDhKoFM7zC
Eppb3EGDkZpRS7akktihiMp1LB+GiwPs4cd001aE20SVZyy4uOrvOdr8EEjdMBoz8H+EwWl+JVD0
/E7unaQg1D0HaeGJsvBwsvG22WsZDUgtKTzo7AFF7etzqU+BECsWV0aRw58ixqBJopllLNhFn/7P
pir6Scm+ay8WAS/meLE+Ubguk4fXNuVtFwGRdEpEdnXW64RVQbjDS3kTM/orlELJgAETeUkEvuNv
O6P7cumxjy90f/rjZizM6yDiqcpDKwZL1GrGxG6MiL37w9RnZ4w3xofQP3+Eoht6fl/uTuPYG80y
rOTFidKTnqpxUuHVWcuYGAgHC6eXYyba1IevWGDFTrR5SyLB7pFm5jrU4H/zfEuOQJLTMK/fRmad
tGfny4wHGoObTK/HGaO/qimM8nOh6xnHxLMUmi0LFm7f+sdqTO1sZAPqA1uXMS7t2On3+tPkTGUL
jy4KpfRCpxlMgdV3L4/OGiZdHFtK8MtHV+Nc0K5e1okzVCfNmu1vu+GWXbzBOnCQkGNtyOMdwgcp
NGQ/3eZ1yoUFGZy1Cjd5xI9CrCn/94GtIZFhXiUyXJOJ1WxRnzwRvCqQQcrEOqn8lDlPkuRwzwgq
zn52trwW/V58QmMoqrlB+EicZTYiL75ku21/o6vF9XobLHDTpSWSfFtRLjwIEyZqmAScsLqCTaRm
Kfx9EowWzT3fNsNcOtfh5BJI1Og3U6CHivH6jMi0vc2NB/Fs1o/TMP+H41AycggCvUp9xIeMtwtV
p92XuxpEzC4LVK3fv0yCK2FoHUINSgoRFgJNcWfcqMoZrFXynAKt37QZ84YG0V4e07y+s6KGEXux
y7ud3ArUlkactFgDKPnFcMVUfTIF6zgtYTFK+sN7c3CKIMd111tu1AI+dO2me6aP+wMX//0RRRep
8UFePVKdtdrpxLdqUZm61+g7VMHIfh3wjDI88hj0pj0iFIDJD4Ki7vUj0TDnkPXSFzFS6Tw/GIc5
koDtCIJPyJ1Ygsy7y11V8e6cnTmc8Qyg8ntGv4VsCgnaJ3NxPT8/UO96HZQx+tpFdy/30VbG/oXm
es8oxJDkRdix+irdp+nX2aP1rMedJMa0bRV0dxjbRiuEpHk49W427QYa9+OGVMrIaJG3wwAz3L5I
GMyHpnp8yDXvMwJvJMkpz21UeysoNGVe0FrDyso0WuOoiJlD9sufLUsObmbDX5ptWSVglfDVyTdy
n06R09uGvhwPACEnmMPe9BPsSnV5+Bug6vDaIoXpyU9r3MoSVDpPViCOsT7yi/JpacMAKoW2LNFU
KnvEdrrnV1G8uiHlObm+ydD/2LL7+iEBkqkyNXaALZr1f1YZtmG+Z4bDWx3RJrxR1lB5TF/NcrES
daaXtVoK6caJx/YR3OamsVGovyycs+avpD5cmx8j/0SyJLfXZ7OcTaKJXwwJmPTmzrcbt+TjceuX
U5Dg9kvXlSg7d0qdEphUbKC9dPfSfP94ZPWLYhh+vMQfEXrExy0a6kHA8kWAgbc2yHyFo19p6T68
lx07kRTmPWdjWtOUdl0xnB1UtNhi92s9PjjbXezq5ehQRW9J8Y59ISGovo0NHZ8vXCAaDP186iOp
Mp1km29w4GAIyVF4ukKu5i7KODXEAZoGGi3Kfx8Jhj8viNs/QWn+3i/Bu5kDYkqZ3kMhJ2SvTakH
Cyr3koCnziPah206tFe5EezDZFXTdYarDYvsXBvANQ3gU0VsnKkpIcOneIwJNGC5Jwro8izE4WtD
Xcx+fBE8jfkckHGNsDEx9ZHt+tOnthFYTddGPwyLbh55mkQZVpmY2W+l+wf3YDT7QcfEt/ygvxax
bMhebo12XHb3PDpY3atSBjlYe6MoJ0GiQroBTdLV1NsUaz6jNqwmmsjqTcYSHoy9S7znrwRb7i6V
iZkoIDy6akxZc8Pabj+JhS+0/SKl8uAS/UBQNW9bKwBR5++aVNOy5ogcHXatqykwpP+aAuDjPOD+
0zpj5uZo2C2NzqKuxp2o2HOpX5mrHLsTJD2cG20ySq4cI9HeY9gz+gHPWDgSdBFta1+2joTXCR+1
8f+dAs9rMrrQ2uvhY1NB+iuXTZ3TxAfl3P9rTE811JSvY4096bVohSyzT4mROST6AC339rJOKV7/
zSXQSqD5XZjPy+V0vPBEqh8KzTi/f7HuzV4sN3IlxdPADWHHSHDEonrdCtIaPNwB84Zu7nj/gAvc
AvHKHYakgveF3Z/izKEXi4mSymGe/uy0bHTmTKeeRJfA+qAlx38/HCVbrm2pnkU5Y40A14CBjpn3
MhZXfcvW+jLev8xCCciYuVi25a4UciYd0TKE9E8U4c8qm+uPFOAIKCmg65lV32nOWgAtKsKnBTIH
v44tmT/PJOes/ocFlIAM7OtDKXms/gDT57mIt3eXouy1ESsd8ZtdMOYByg6cij7gGLGCQH4oYQh1
FJGJLNbRt/nXT1EUPO0B/ntxaBr0MLvcfLQopCp4+WIgYuso0gV/3UqtlOuMKkg5wuvZeb2to/g5
NDYAW9iHwNtxkzrQVKjpt+amVfE+K0Hu97bkda3/RF0aPJz0dTA4pB4Wf/ndc68ds//5SME7MQue
i5r7evI2BiZ37eCEDZdCKXidbGXWsOzjNLpVpm2Q6O1/4wiJjviAnME4jWcTj3SLTLACfMWrfv5D
y0E8uNdVtu4CTUqlk61QeTjj64jn0UohiyqZnzQe1DpKF5D682Bjtj022HXypGJKQQIJsQh0qgz/
EdndCC5nj1mzh7tBbFA15eyOF7aId6et1qXIdm1GDPR22ZOvFT7xr6kVbmju+psy7ZsUou9XdpFb
/cX0cGmfDv6TCHB4Sqp8QVCfW1CAPHtIyrlTmtTRsxxdIixGTapQfCD0CkE8PxMogHWJ6l8BvX9c
FW5OFBSUU3EL1GHQGN2si1PVs6d8COtUzsrctxoi3JO5EJN55xGo7ZKgV90EdH6KKRzvosKBG21k
++TW4Qa3EJ+Yec3JVOvFGeww3S0EyFQU5pCpZXZ+wymQa3WSkujeMRO8A2FPiiQGjIHF3sbLdmRM
qt+Evu3GsY1zWXHG21nuFfmZUPweKXbp8OcRe8bvLsgvk23bJFU3UjvFVLVzV5BFgIkLJKR/PI4S
DT9Nc/A5TPzjBcbq9kI4kCXLETACyGqJVJ4EG4rGqoG1Cd/7roUOJBuTka+Qhq0rXZjob7dCOr97
s/aaNZjjoT2v+Gpe7aMoeROEQhPbIxHlCnhkXAVu/dK3nlKdzHjY7YHeiBR7m66ZPGm5Q2pr1BeN
DH2MsRInQ0tcZOXixWVp/6V6JEvKckyORs+g2X94SoUHtzDduXlmUlYTeb3T60Gk5MhfTKQTW4jP
wAediO6TwsKGky7T+A41tmQxx2dklok52Z5GUtuRo8xhUcTwNwGeiiq8w051APEJU5gYCqMQXNuV
xLH4EGA+rAHYVjNf56q3p/1BhmeOt351L343gQIrfF+fMZU4eRRloP/eU0ncvCVGkjSzdnvxUNZz
j0hCxE/Ni6ZhFvtmmrwcG2KSrodAHli7CIk1IY82KDE30NI6Mw7TCxwUi+CtsMGrIS4sFRBWhZXe
OBj5dgGFH3QNBqnLNeRZVhBIcjWoj7DC2C3WCubphnxcaXg38QCC0Mup7H0yVk9BroUgCEeBsPd7
6vq3/2Bwt/AfdF1C7zLpIqhBs3XfYIg8uB6mi38RyEUA+1N+aY0kL7wpg8X9149Kzls7+IqxILYJ
hdMh6AbkEKtyQreTLiip/ExAPsXb5rvzteMxm9LpfPQqgqypD2gzhUdIXyL7m+abusQSBbfu99th
1ywHSnrgxk/SmFK2A4BdBfOZBTzU96jBkBWdleoLiuLS7lCIqIb9XqWIEWCMLK37Ou27Hj3YvXBb
7FypwRuJRJXZHO5aLQgeTociY3PAZxKxyc+r+oTmmX++zldp7SjPokivUkRFs9zzJ/HnfgUTqqQI
PGxhYGTcWXN6nNGrUMTSbHQvyN79fqZVFo03Hpb2zmUGM6I+aIpANGJc+vyEQxIkeZTXMRJpNQxt
0Oot4LzttU2NXrt/dsyapM4yV+EmgsfqN5kgCP9zsasO+s0roFV+Lhr9cY0XDL3XW4hpycuChRBS
sdUHOOAJoDxdNOYqfyHLDIeoJ7wMsKWdQB4YljDoivStn8oNOIPy6YYQvyCuRiGkzyckgDn9iAQr
iItrNiExy1Y15st+0WIgjziudTSzZq6kUnH6o4PzM5EYPDfg43hwBxqf3l+TnCHF9v/ZXsKxDMNk
h283fDw55Yu5aPP49D3gUMLLmQnKIfclNFsZtWEMWLE5LVR8LzqA2MkAK7sODTtXu/RlMVPvgpIQ
EfPLAsb70tC+DrQxmYpONu2Wx1Fj/P6aHKsvfpEdP6mQ5EjKZJhcZ+ijhPqW15Kv54fIVCidNdSW
Q30Y1vvKaQEWn+Gu54q3/rl8f0pvV+dpvgY7OS+oXcmrH0b/T2bT9BI1vqD4r34e41aYYne4Di83
tguxAOulNPg04N+JWyFb8XxR1gu4nFciURgVfRfCL65vJnrVpRXRLFrqh6YWtE0V2QQhz51BGYQ5
d+MFCUHRYsaeHQkHzHsnOFjZ6SNKV+36LO9mR7MqrkiYcuO2dFiDABHemTwz+eRwoT7G21cNKzw8
SRobKgLvNRyYKuQmYZNvT0zNndARrR2QIs2kNA07IS5s2ebOVsi496RQbTQGCNN8nEe+a1HwuWgY
Z6YF5XPagMSkkvsbqLsEhc9RqBaJhazolmvbDsL/4hRDEBeiw+UdaDHfruL+dNNQ7sOdPYVAZdWK
4n2VH7bPKhTvJg6WQhtkpVUJ9QjVTmv5Iv7I51iWM9xCmJ+/iSUqwl3EWp3dX/qVoAWUNMHfp5x/
mLYYVLHqAqR/Nj9+znXj5DXYEYIsajixG9U6+Y4ky4uPTcCoomgnyRI+pNWpfEhUWyzZGyuiS8I4
xSnJDz3wUA25ZoAZL17olWCXw5cAaQEaGA8p/vUtM4eTDJ+ePo8arnnkv1EvCo5Q+NMq9PXKOE5g
NCnxuzQeJPMoZBm8yF7ZEYXVlk1k0oi1DRjh11B8JbXigXyhFowo/EXVmHyuLQ63/efc9aI3cGF5
6HCCF0EfozB3Y6zrC98F3b7j5M9yR8E6npsdogNBSg1FpQjjsvzfNBls1H1AWTYPJzaLA6VC/Btj
0BTOkYVz9X324x1k9ql/zt2YCmqZgkyNux3nLxBElH5FeN82VAWyXwpSvksan0Tnu4iiXhmffnDt
jrtLBChtcsArloUM6GgF42WHy9QSeDvU56vUPivSI41pnEuzoQJgpxFbd3CTqwg2oJ9tqy2ShdP+
B6maSqZhPEanx45AWR+49DeNWykZ54OEKJ1DGc40RlAXjs8szxL6SJBWE8kHCbuaOoFA0HMHhlug
EqFyhjLagVQ0Cb8FhmYF+buu9+AkqxnCTzTTscyG90UT5ftWYLd4HxWP13LSj5YnKRTILQmgL+T6
cHwW8aAYZXzJNlsg/gGRLD9prndk4pTrQ3KtkAY5476mAoeb3CiBuUSCRaVzCbluFswaUKsLAHDC
jdjCA6NNFX5eg62r+61ujgoI6FZe8bKw1ROneSWmmBaoL+2BxUjKfiacly3Q/QjYWdSJ8f27BSLQ
oOOIEP1gz07wPU7QMqJpQoIp21J2xXa3lznKx6t0ZaB99MHslwP+Qcww3j9rXVZE0TR/x2J02gzm
j7SyLLkH+iiKTKX8P6kCoF12YDSe0Bx2/7cEFJlpBER41rBh5O0G5PkdvHJRTDvsZNm+CnEpa4me
nESFoMIGwcXpPXxBJUZ/wFm0z1+HePkLSEeUH3bUV1l2pmNXkrHiHTYjq36KdfUNnsNtaHqFj/SG
sngGnwxEHK98Zs1K2YrIAzhtwBCwuPckKKta3c28y5xJ1RYDwl0Fh3XYRqsb17hcTBKsz+eQpyiJ
k7+RY2U+HOVhT5Jl+vh0F+piHSLA9aLaX1Ru1Fn12ddPNcoZW3HcWtIZuS8sD1cveZ+UThNk9R5e
1HqGKoWN5lxGjMrCpXxkFUj64aNmn5JcLXu5Fzc7WWGRf6k8+QQiVp2b6IfjCH8LJ/FQZWgZWqFe
z0qpx6+lmO7GjXGmcSxGKFlhCfUBCw8zCZk+fa0kBNj+Qb4CS40erukBSa3X52i7gm3kKoQB2yL4
47oA7WTzbhLOALy1KgUMf1Jc7mYTLnONg/MAip49OxNSaH53blh0ehzAlIYEqKkFGSjSOgOPUkPU
Obx6HQaq6t62LZrhmI+0qT3jYuY6856CfvAQ85YRGuDfKmJ8kUokAwaNI1qPPqJYoO4VxXH8NB58
dPZFw0emzRp68q+UrDUsYrPr/m0AHkDbbPfHdGs417Sbrc7cxwVE9TEjJTb/2b11L3RCL/6nAQ3f
hq/IhUQzuJB26Ma0+av9e3j3Wl1G2FKJ6g3RBKzPFLe1zVenJrkoyQJGzsDygy4BxiNCoXHc3nLS
Q/1vaCZxOfSqdh8otYqIV08Ea6kTL5GdPmJeoDXCw2su9YJ4mWbCsJ/Ej2gNzfrsa0N7RmNUma8a
rrWONz63vedpnzexxQwKPVQk1PsKU1M3O0UIxaemcv8FkpUSImLOJ/KzohsByJyInRC9+dh7UejW
Byp3WIg3nNU8PX5njI6eCM8DK3Ol3Nw1d3gj94OMacH46T9bfGb9GXoFlF79yEZEH4m8ru4OE2vg
nSKYISA2/9xy7kl9O/VZsv1u1t7qsF9rrzIsYlTHfd40ewjWvAPLoHz3uYGRrj13ZMWj87DmrwN+
xy1N+RfGKUd25zWf5KMoj76s0Xpz7YYTQ/BPvoxxC0wV6OOHDp9mIQuo2pjv7i0/nEWD6otEoh6P
HqZD4wCXk2HqVkOhJp25duACdCFXljsJJM8X42X43HEVzusiUJ29NYkNQq2Z9IQowDjbuqMlfdhy
nW6oedfjXCtUn3CAfppw6yOFjILaOGJktzBa5XymjlE1sWjEIutf6LD2292ISUyf6BT/eYqea1Fp
6RnHy9exFvGAccADNd1lQ8xBmjB0otiszhHW1td0fgtj+1iFt0WLfc5dmsE6WcNeR7Vd0V9M5eR9
zUwFaQRhyqL6QA05AzSiD9ewO2FNPZuRMi7UI18eXdXFt1mMFZZK4gYsnLZQqhbNIBukUKnt1Lqk
9pz8PknvEh2Z5bp5g48nsOsC7ymIE6CfqJzPoWwcTTda4d9qmFDP7osddJC2aPQy9JrlWgSxJz0r
v2JjWnesQ0UegezM212kx8mFnq3AXKBIzlIjQY7Fxb7+JELF6r/MuNLxE71lk9kilowOmIWemZmR
bUMiPJqoExZy2x7pFp/LXDdwPGG1+VHYFkop6Nlpz9IFQllGvwyh19VYX7bZbK29isuV8DJX9FRg
hL3qXtupIKvepGtRI7ikkqJLq+1pDejGX070MD2kyf1MxdmJp7BUCMtWOT7xKCggg0WkGaJZ4s3z
2CAAbCGrgilQKaa4C7BmnoreKrbdii9wjCBzVkE/rhbtq9rl/GaFavw3iEzax20s9zPlWELDbLS1
uc2j0ssZaPV720O0yJnnZs6cc2mgzM1C5hLVYi/iRFZ/1fEwp21t0MLVqZwbyESBIM3886eXNA7B
82rCl8bk38O9CxafK40hY/ThWn5NvB842e35m48wha3fu0hM7KNiKwchI8gvA/yTHzrcheKBUWdz
+9VgVi0+byyVarIijuKOuimH2AqeBS8dOlIQDT5x3Tx3Kv8PHzKB6jR8P9mo+xASyRA8LlvwGpro
2zRtMijSb7XJLZmj4snQlqU2aVy7IOboTTA/kkNoZKBRKTTSy4eMPgrWnzEMaywZROmZOCGi2WTX
0P/TcuwNJP52LxvdkETqNLqIe3VpyKH0JwSURqnFlkCX9DyqP9wkT9id3Xw64T0NfKi/BX+8Tgus
NzZUy0PbEeAL+lM8RvYBUDp4Dt/HbLhh+d632/UJofteF9h1ubZEvqi9cqiiFN+fMMwe5WsI987+
YFSeXkS79pDn8DaPrQPNbpb5Ukq1g9jTW+kIDiX5MsQOgghIv6CwaM5ybhoBYpLX3hlvvdz7HSDY
q9PFxtgnrb0zSeRvzg+YDAzHV79NcnFDOsH4Odbak91/ba0x1lmEJl7Ku52a4uFnvQA/9XLnAdt0
M8IKjsJoKUE6ltaW3NaacIfMfxKkkS+NSlxSPbjL1h355XNbGS1/7TyZbBs972XzJczpA9p4gHyt
AKZtKcsOgfIz8WH/RqbgG7GwMmYA/yEyEQjrPsvuiFwfNT15DATWp7mUI9B2CEUEcXr5g44349Iq
nt/EhPUc8ZYmE3enUtuMhLfdJkHVmXYRrZ1BUg30LUEgyiHLNnQhrqWv76bcdsbGgoln90iWU17F
HpXGcPAOCdtA7c3YEdz17W5Y3QU99LwyZbyZip73YTS0uUrs2xT6hsVqbsBMECacJfrpTlWYaRDT
cdtce1npjk3Qwx+sTgu0mlzKC5CF+lNqVxZedCYdnm9yz0DNIJ/ZqwtrtPG6hP65nZhrMBYe6F46
DxfK+4Eqk3bQw5L40d4hwJ5Inmi7HWJTA0I+5RNTSl3L4pyvmEt8zpJnzwewUK6ggHsfH6LGiy7o
dlJsYW8rV4AUThSSJny4qU3T2JpEBU6Pa0pk0Ako4rdQbGfi8GCTv6lvwFOe+H2E4tQhjkZ/KiDk
lGzodoQXGvS3rmBpqAoWrpFpVQt95uootSQ+5kWKGsfeIz0/swfUdYZi8aIkZQA17TuTISfWodF4
asL2HkgY/akn7cz5muCJL56EaOtvlgLBDzP29JKF0xITbsAHTe9q0IrZ4YdYEYHAqnGmfwCH7y+T
R9SDZUzKXfzJ+MtIOqn6Q5gV+d9O+Wc5oI/k/5qaA95J3+p0Lc7nX8cUTw/fJKWzdPZcC+bwMWp3
EcMOow7HjNIBkuG8/aMmQgkpyWWtyi3rb75Hn0ib8ntjcHCbE43rfVz84tEk0m13QiIgl5pkM5lo
raK44IzE7AEsZ6E6LRjdqQ10WmM7S0S/ObZSqrZ/3tRUJE5fbh0jgsqTMk1gSsY91f82Oli3WM5w
f9CmLausf4lTttJTmMCQJqOpO11306AUeZTGIzGey3aAh3G8aFYJxd6HgAJXui4Bnomd1a8/N1n1
gtHpy7/eS925QSY4AaKaIZX9feXi8MObB4G5XqB2tYellqXk8Ei3lYAMrhmgy0rxd0Ou6BaVmI0e
1i4M/jqf1EaIFowM4en/c4o82erDFiBv7tddgs687PNCXSR/LEIbULXCWeHL6raBek7ULOfcTdeW
Xir5Ajz9xsv8atre6hKddqfqrqGbaFk7OU8ZCG5XMJqm4hUYDNbWaOVO8E5A7oYfa9CpB+8uu36B
iEZCEN5jDzlWRLOZSDXT+MTIY/wCtdzGaRogAxqwSYHArburoLj2H8E+QXZFX9HjwCLBxKQQskOV
2j9n7iMbBeGFGKRA2qZWs8PTXrw8Upe8p26tL5lIw3x2GFiy+Q+fkduChx0hFRk0rggJ1DtY6kB0
L0GEnlK15n2srGkbrLDhmNVZo5pjSnhpSQZKyklToiVT2Nrr3Vjb9hUgbXuBBhUXHaJDwrqQG7FQ
b2l2MIthBmwP+RGmOg+kTp9m4kvS0ORW83FX7V5kZIHOgI68yM91eYZ81NS/ljlATV8UOVbLxA0r
aillWMH7m5VHocLDzdjWwq2Jz/jIzk/hyUNRH9B0T89oj0AexwbGwp+c/IROwN1/WEIz0TKwO9FT
DukFE2jOkB2qka+lv21mRWnNjWGdXCcWe1Ede8BOuYwYxeT9FdRZFMkjRM3FHuKSWYFfkoBf0dk9
F6+zfWymqTDPo6EFTqqDVz+wLLKpWa6H5MyLqFb/5cfbKiQ1llhz9fpc+MwND4cCs7mtZsFn//dM
tSzDJG0kzvwbMsVVw2ig6FjBWiojvg1GddsRv4CjWaSFzuhxLA+6/OxtIe/LnTn8kixQT32jLDHh
nYZXaFJU1rCeMvJs+stcd7boKTIR9qOD5DUE2mAoiUUDV/5BN6bSG37/12Oe3YDbDlh9zkd6ei4M
JYWVn8rJUDYA2g9fBYm4YfczNdh6yyDymC2217UsbzxEYCj/B4t2+tXvjH7B1BFVuAPY+11H0BFs
zHFA4+skz57yVG3PVXRl+vbfHhjd1qbWm1FPm2cN9DyF/qJ6KVTSSvaOAFq1ZwqsEhqUmmZIcOwn
Qi94eLIi8U9neAcTVjnSWWWLF9+TdvKLqvyGTYNIqIsH5OqRziap4VCKC0T2aB6NG6GY3rAiGMBa
e22UDi2J9mW6KK89ZFyTGnzCcgAO5EYHVsc2aR7v11GL+JFJQEw9cYeNdbtlwYA4qK+Ag3dkVsNk
r2S4iODkpI4jjEAmTyNWoE4Yh2U60bppdwyGtlhJ8maI+asrkAuZKpqb5E0IAsmBPC6BHnkdL8/b
+V+Fs0gY98QYPSJJwsyY2FIYk4zHYwbPpVnx1VEZiIM4Io8RJARcK3He+74GS9lDnSlynAYUk03d
jf0oKi9dSjDj3EilyGSkpGu5nzAR0z90DAXOG+tbAuN164ZoJu1FiVkYCzKjw9xIBH2O58xdLTXg
gVCt++7qiSKB6cXD7U2x+muF0SLGQkrsNHv9ZuCGlyI1KBV70w8b2WUZKJtvzb/Yx6NWM2vuIaoi
4Nu+fFnK9gI7+gtBxmBfDu2pKY+vL2BOu2c5irtgEve90Qqvq27lqS0qEzLzliL92bB+gJdryujA
T1eceYaCDciDd8lDLV73a+yTCvcUg+tVPywKYHRv/LfEtoWK7wzk5WNQb7fSvg/mbUIeZmSIYMXW
q4XJR+R1WjRmBlyBDEEhRKtek6baqWuFbJZ0yG8/n/qC5JYlTHzXu6lZE3ifJX+zA4kz+kMYvnZi
GY+Jn9CjTmsgvNYIVdsLVtv2PACtcZoxHQLjMTV6rvneqjGVfms0FzOq9yFphN/D1We2YRbbad5c
BW6Tq9f6PtT00TDwkuBa8hnofCF/DctjdjGbsc7LDCpHKpKl708XynZ4E8iDDLdGrmxPHJYRJ/x+
A52YgcrjVmaEdEWP7MVmEQVR3l+LnMp4zySRCzpkTj9MnKFXGFvr2k4hX26sCtDqPYDMvKWGm/ru
njWAUIHKrot2LnnlxI1Ndz9XBatQYAK2QSu1lHFuqnGSh4h4Z2k6tAJ2ukLQYuY0g8hkxabyS8ve
VR3OOSZ6zXjs8qgXTAiQSv2bQ07khJvDwaRy2Vxl8hgQ9bVLjsQp8vOWPTYSTP72Cez3SLbP/KGD
NT/cQBxF8NBPI8Iz+IBp644aeVyqoO5k9uNT7o1vF51usce2JjxUM1jK3CWJDe8AnTKXu6/Md5A7
7MTr+87C4lr1gO8F7mJDI2YFDRGQBLfxeSeqAcgvY7wO9tcLVDVu+iYPcnAUIZz/nO9fsmtkZ8nR
L2yNdIvaLK7wvQjJ1JuV3vViFanzz/5I/4pKwlElnZhN2TinRcMb2dFlE/wj2otVJTw/P1L0lw08
8YT3bsiLCCPV96yNRdT8/T20NPIbBHjUwm7KmD384wGjDPZCqtuHPDvDFGnNWZuVPLC/llsR0+LP
UpDW0Kd0LgBunNkp8lU1ZP1rIQjV6G264m++GbKP0+awqEU1MYhAYaUiBy6z2u5ac7Rd5vIDlZ7T
DPkqp4f4sxn/uHdTYx+toX1lb25POP2TWW//WAimZiDtVFxdaan9L6tvdchtWzztxUVhP4MdiwXv
FyB9+TyVM1x35iFGz+kJ+cMxxv3VRxFOv/q2E8V6P3d4Pm3cJtay3Om6XDiYGqfT+crwea6MGUfF
BZz3cRMe3cqEzPNtSLOkZQPzGAyLdU3cudIGYPjJPQFbV7DsdjvsW/B0b9DInc2TrIj/WEznej1y
ozk0CD0GtGPZPuT3/0vwiTsYC2XdorOp5WtLcAYqCwyd+xM87qkQDY3ijE6iv7ifEVGG/lhSBeRH
mjnV5M5UjcxKaiGWKwUk3cXvmv8/ky0tKpC7jOoDP5AmlrO0SAU7uvuMmOO8qaFmwH+vefh1juIA
Eo1NTKT5JsjpOO3BBMCXh2A+UkqLKJD+R0NyMyDm12AbVMpdj514Jd9ajPAY0+GCWwG38Tf0o3ER
P4Y1CGCjCJQmg0M5nrks4LWgCE1soz2t9s6xCU/68Oc1kkj7fCll5i/OyPKjUX3mE0tBY47kaN8P
/oBLWTtviwAccw42ykNNifmyLXfJJMhX0Sc5VWLXGCVD0YLTXgNWiLubkQ+elE4TJMJlid953yIa
XxhqEaen3pgOgFIe5LeGegtoj36jAmlpjQg8dbrG1ZVSJRC68q8/8YguybjsOlexS70UH8tUKEz2
fN1ERyGGM1L8bU0Ozg3JMGNpc0pDMb5bCcxPzxWHNMHRWdASumabz/X/q6Z//ruBjSJEAOOZ4TW6
m7hcBB7XQ3yqL1//kZaQ5d1NQLdDcHN2pPgrkovNtOB3upZhv5M+9p3g5CTNzEVlCfE+aDedAt/G
dyGzItzWqJ29GpVUw7B3AIOw+hpXVTgKZeHN6IoxL2D5URQ5oX/rjSjYIpelZfCCBWKdOs/4WJag
pI8uaLXKTPY7+Jc9zhwz6vHVTfMgYEDotA0+lCRWzBoEHVZef+OwpH1NRyB+yhyIcpwb8cpeDMQm
w5dFIxzWGLOGLRBHO79gwwiuDWSF6o2z34ySSyi0US+6IFWqa+YHzS5StEI+9HbtftPOid0cKkVO
a+RRV7nQSu0j5yDMELpsRVg4+FpO1wYM1eqMn0B5X/W9aH+NOrH5Ck+3stVvvj8qp1eF4CS8k7XO
zk8IBODIIcqW+6BGnyKzAEpSzrx/5IYlWse6FI1n9r1lVu2FaMkLgiHRb8zMCiR9PXTHGPeWLeaZ
6LyBl9KJNcOLE/ZltX1AjS4KHWa2r3REVOcfEIA4TDHM7PqVaoAFPW0xaqYmVCvCDkyq/iqPg9H7
KDZYj55o5epIfFr89FtRw3YbA3q0w/4WYpCDAPSEMPk9eaTVqmDa0vdJbmG66rGx+0flrcoLZzr+
iiT+FI+c2YlcofvZsZRWAnAxYqgPqOP1FjYXgJZ5uqyMDzJY0qWwgHlFda7Fhva2A5rWF0U9Afo9
PZGG1h+YO+YVi36VetJYQ+unvzmS6LadcBOSmzAHkovTbppTb8hHfn62fm4LojeSIPsXZz8bzgzX
uyt+RVbeaoGTlEtc2anJCzPUI8we9E/6pQjHAIj9HVfNhzbWG/T4Hvb7a0zkoeMzJn0uEftPN3KB
m7l1qThqNdAfFfNrysXf/NmvW8r48ggNW4imQdFRohv6ZI4pKuvswgED/gy0KDO/WvCBhpQNWimT
JNv1hhkBa04nxlooNF0CyUh3zknum/7c0gak0TNJTUKEwS695ViN89dEXdjU5PI2wXvxXBFo/DCh
1VS/Wh47E1UxTAracwB+fMuhegf4GWJAXTCqKOwcbFcbcr8s/ReRSBeyeMUCTPrUqttukGJptaA5
e72omf7IySq3rxN2W7kMALu3LxnVjeCKAp4+i7zEauxsQfJ8/zh+oDsGCy0Nb9/4A4qokyCMCWYV
FLCk/QnYuJmZI31h0YjqcnL7+te9ksVGOtFCQNz8dRct/YsficcNeOzNsGJb4JbERROVRhqavlJH
+2/+vHMEn1TUC2sKZakmgYjv6CXsczVfmA9Fu0bA2m9Ki7d/3N3A8hy7Q/53aSt28eZP7Sf3/Dsf
udbgt22aBnJzPu74Q/oR780/uVBUgMI2UhDLR1lhz/oKtwMYlgQELPRHsywvgQJtJdNfFaD5rO0t
b2aXvh/pjhoUwO8MIqqCb5Zm98em7Qt/7VnJn3+792AsmGmClpBYlfc2vQRb6a1hOIKvC8eKbYl3
pcH1xJih/AnErSJAK6bQM4lGRgRFpLrj+5ekI8JkdwaWyTdWg7Z93HkGoyxCzBTJ5xJOdd85ODRj
lr7Yutj1BlMs++tUcyu7tIONs8EASKzz92XRM8kTjgIbmv219x96LpdtP/cJM0+9wB2RdtE/NgwA
pBNInlYZraPDg9eEMLXoUO60Gxp4OXY2uWhQ3i3MkMfFKVLXofNcyFFPMay3vrU09GGhoBeyeoRN
zoFeISi55AkiWq11Beo0oprv1eBKRAo1G3uWnJuprZ6JKx10mxrNwlFkOyubvGDQmTPoIoIvit4k
n0ZMw73uz1k8BFXRRIS3JCUJ6RPvPoI2PcmcXTtgZX9mHYW1C9W5js1rH8lhIQwsqXp7xgGT2KGX
xVg/jakYPc4+dyFIaFzeWu9VqF0cSru4TBKaztH/A47+37jqwy815MmBwvj1Ke30/NpLCtfoPUZ1
SRu1hcTfkV+TSqVP83XWK9r9GpmwAy/RKeWfDJYO/1Ol/Yu04BWQvclgDP21T9vj3o83upzm1GMG
jvELm698fFo4T2Ccy1jbu2TZGGDzLyKgBJj9MZczGBtFXwRbkw4pdLpLCqL4duJtUtlQyfbFRjWq
T6QBESd+NvOBKtczKGmwxsqiQRhQtWuJoEw1UMvP0Xpu6mxvo8cBttYSfDs0p8y2muZUD23/ed46
AkLHYe7u1yzJCd8pO/GI2wkxtw1+2LT3T5OyzhBNKmqBrn2ru/7srJ4CvrMCoY3xs9J+ZwJTEoDA
ZqqWX0h1ENxi3ypNa9q4vEN43i98ISbhRJXgpXmNPIjd+AwgFvPd1wPVgL01Cp9mSrrx1du54iO0
kJOe3HuaI25kgSPpNcxownFA7+DPC0quVIK6KSauJBTXekZcxgWWGeIk9lEAIdgyxeHDyFxjl3Cp
JTRgYTU8NkEypawsETXTy4CCM2IuN0oElBYHa1+dgeaSfeJehg3GhjDFOyZN/6E+SwMDhyK4OxT6
c8/P3di9j9U/xRTt3gTSUOkCJRNR9/yF3Ajj33IrknngCc7aOoVIqTsJHupKFeqNodLhlAGDTe5H
62W2X0gOjHb7lpeTfPCnHQh4TGqVA18WZRLG2DbT64W+rj6f5oIftCyAM+ZQ6ytcY8u7GCk3qajE
r43W6RZu0uWID46ma9h5V4qatjiFeXguMxUP82PJErMwvmwXtXCLSHf2d6GzkhaoldNaqEvD6mi2
u5uzpPlYAd21zalOF5tMI1drb8o7gZYloWUym36UejgilCNiqQ3q9GjgDcbBczF+pgEUV6wM4D5Q
ei6vuWD3QlMuPurQxHBIiY2Sq5nFm8e1UaOmhCnlnPHAfx9l7sk5RQVWCz1qWoM7jL+QTzqbyWOz
jQR/e227J+tn9lCMRbx0AXOoziLvDl00FgRQlyNUfiHohMfsb34gsKZ5JjBSZGIucLP/IWN7QkYi
EhlpISI6L31+fb+nL2k9Voc6B3PqWalDXt1U9dKeyPTdUWFgG2YWy10wgVDZtaQGPk74NnMUIwnk
eMSaost/k3ZvookLPDeoOp79FQAYCTpMMiTTGMJGVDZL1KzxAWV53TIQbRWDug8sZH3RFPcWhqGl
ExQIt1pNWGcn94Z532jOWn+MZqO7BKw/CnFtbjZbcK1hToxhut1cLk05gsewIB7xM3OZcbfJTqq/
2tQ2Paa6VZhMahD2VAX7k6rFWlW7B5pdX5AQlTJSpaQaO4gyj9+ZkgynuOfLYYBRLBUUYEl70z74
BgCr2EGya9gMvGapBE/HeH8XpJx/95Qrt+r+ZBG0+v3NGL+utsowfnL9Tie8jJyFpjjst86BuE+T
K9iFOOynA2uVcm84U8T3C/BOBywvW0V/65K5hW1DTJh/FCPmhgV9ytQlhvIFcF3qAlL+x0E+isrf
TnX7vjdbtrbGjRWqgzeOccLkaK8DSVUetR175rx1UECNzmpdVJDvjMjFmhvkJZEYkCZjLW0iHJ0P
+pk6loHd9Hd+kTJbY09wlMqKsKp+bYbbZa9+3dpzXKpoTqAc75GpWlJ+tZEdm5Z+FC4va1ttFNzG
fArah6Gdv3lcSPNRmodIVkAmc4GyIFk+yT7LFk9Debo1kLCO0GzUJxeSl4pLQhwN5B0FwttSxELk
QJPeV5W43CSfKGwRiFBQQAd7G8wns+Fyss6a3VohO7J58Acn+yjwrqnCLAca2vUZCRWV2rI+x4XA
pAjcPiaE7gon5gzwUjyOpkMfcBZO7bI7wDPlCp6Wkd9V6SjnpZ3fBczXDvJxrUELiWIhZXxBZEup
2ZnMZPStR/nRFdqKzz2tGfLuJub+t/xAzVx7Mq0kM+6evdIxJaePrBgnUrhdLhm7hHoxf6T7vt4X
bWnYnQnT89JCSWtnYA0hrVqoePqTqwwLDAtydgJy9/VbKmmrSraELQq9CZr1VxwPsPQELHdf0MtS
l/xC8nZePD/bfxu8Cbn+nR1/kMFKYXagUdVoioYrxe+8NAVHjgcTC1HHLB+slYzVHHh9vNMJK2BX
/LBk5L6Db4EuxZDjgTN6KNDSoFDEMbLp0CxIt82nvzPUOD78R0bdGgtDhUnIOZ3tI/yYpW1/TswA
5OvrfqW85Bg7lNeto4i89+tvhEWXv/2u122Wce/H0nY24nzxuvEJTECmdG7HdBtboyx/UCZ4p8mi
DjvkztqnFBr/18HUuf9pVtBMpRi0tqL45itdYyW+spiDc2Hs9HbaxekuxCyrgTHiZOqCxGGjYeKb
ZGv/U7X31uh8fR2doWdOo573xeVwdShnxv4r3ULkoHr8BUMaaLcTKx0891D3w/VsRsU8CMV7T9DG
TSFkGJ1CGcrkAy9qf+/ea7gJr7sc2HXRgeuhxHek0DXO7lVxhe8QFuOjMprbM9GDj1Wu04iRZF89
LgfarjDaxlgg/pAAlMw2c9BVHaLE+W66gXCbiRwVFZ5l57Sz9PnsZEdJqDUHIbfGQTx0UQ0IK7bk
HjfTkVH/NpEguQIwM5SrdMR0dMBAxpQqEOSFLRIW/rmrdS4Zp49hxis5goOlQPOpw7xpTTmkqykV
dnrB9T9Kkk2gRo9p1rtnaElpzqv51LkDsiJEDwUl8QNOOZaTqLZXeX7mOd5UdyT3aJlsy1dtIBJE
ZdqeeVOQS4UtaUNBEMq3wIgqeZ8ZryGO8crJCDlpw54onR0Wt0Dub0ofb7Kce8hUREKH5XKrGfb/
lSIxyR9ApkawAGD30BWsPCe9j9AcN+Wdj9iLp+1xOloQhBPsGR+zvar6Yq+GeLgayiwSTHLP66QJ
O15eRt+vv7JJ04ok+anhPz3Bb8vzKMfSM+d3FM06qm2DQbIb3S9Y07x8mF2wkcksZd7Zy87TdwaC
BoF5ilO3Xxk9UhUR+nGb08soNBoU4w0TT6VAWLAMNm7+lBhxyEubF3MhEsmX2o8V4+u1kzwuFTR3
+c2mc/EQiQFKSAJVl5te5CnU+GK+/2Hr+S1XjOGkgauqw2vgN9oeFt7ITeRwNtxvWYRsIJ2QNRad
Relulfwzt2/KbQzoYWur+6ELTzhb5cBhzijwsawOlx8uIC9Uk0TmJUTwPSWPnEUGBYUO5QHsM5rc
MyqaOajwoX2/HqDciAdVzhAWG0UkgFurTOY28iHw3+2HZ6gF+29y7qXrbhM1VKtAsnk8yhof2DZy
lx3ugv9ljQkRJoa3kabXZRN2+oSecsJvg/w0PnGmhoVXIqlOgPmHbE2ZdQajTO93DijJEUWcxFnp
3qM5SsMSpYTmF2WHwZXLfrSEEzKVBZcvRp+mYOQfmtyIpWLq9mgj3/io5Hn7VtPqe/SRprF9gcHR
8IC5Otf6fcBNd+77pG9D0Q83Y/kJ2jmpcEkaiVwxn0MCPyGemDj1Ov7BT5zD5R4TX6lWFLLHf1rA
fPyoH5HEox7qKIx72t66cYLoGGR7USaSkns6gSHm03uKua7V+66/7dEPPcFmtPYXuf4x624L/tWU
tYj4qU0DyrgizIIvGkvRI8yiH6PG+hvKkMuM+CUtKwWejcjr8DBVVdX2Rdcpw6rT57ryDHqVg4+J
IreR/M1qc5FawDdZNj+djBBNUuzJjsgfZFRTOrA00Fop1Qplu7ASKG9+Vl1DvhD5ESqKPWK5IoGX
OO0UuAMFxpkX9aSvXNqNT5sgMQyNNs2LTe7jfDBzm2LWRIXMKGw1Q0NdCjv0gIENnuTRaTp+RPOf
yfQPjuIzLcwdrO66sHFVEcCn4Bvfa/u3RE2SUJH3fxNXmceBDyuAkn/7bFeEZEyCV5k+fGl2UwbZ
PB2ms/Zbk08iE++RxEmVJU/oGP9Yb8Oq5dHWqtbsE8lBqFzTZcDm3PYzh15xnuCC3UWdEBFORgRi
YtcMI+e5kRpIFFI1JM2zTsuuBnDaRYC1wjk9cpCIOt2OkTsT5Piy88dF+UQv6zaPKIO41RcK9GkO
C++Xz03a1wKaYSCshbX4+uP6kifm7bBNr+5Wn2rw/R2aR8TMg8QP6S9S5f0RYQAUZT+pkXExna/E
G+qiy9smezVQR4K+5iwhUetmsmWPKvw+ruYPORaNMZWFmkQVA5j29iEOyEd4hJsJpZPXiY22i/ZG
HXerhEP9df8yiIdVBZH8u3V/IVAoUVyVpOd9eLjrw5rY5q2sohtyS7LS4NAOub7sDmBfaVD5TB9V
m5t4p4TRTizpEoFZgVstLRBsc7felSy6p1gFjcWgb5tbufPjup/3Xv1B6s2tihvp279kKR23beR7
3kVJq/A/RMs/a5Ym4boDT04Xlpgiru/OSuJL3A3ZZSQB45x5KprJ/DsPEP8rcPc6dkt6MGks1sYL
xw5q5GlRQVfB7BgYPS6HwWUlx+xUrcfiM5OyJREdIV+Qga5iDWM+yLHmjbhE6A6468cYNptf+LnE
IjH+9ySLUIgNwop17AYZTJVyX1vS9ZM/dgEV9Y3i1ufskoT9JM5F7T0dCtc/Se9/dQucisXUFMhV
Sc8HtrkWKr/q2Noc1cv6I92XKAhskpktLCQiZYMOB/au4b7+lmYiLpBOGdVKknzEEJJ+Ls31lglm
ECwifSX7S/FGQk5oK6xYpmASGoOV4arZtgBoBv39u8UWiuURXo6V/+8s5RzRxhKpGFGGiW+AFoPl
0P0k/zVJWeFVKxRUl5gIRaV2oe161GID2BoOoOXKFZq1+PwLRPp7to62UKk7bReatc2uKqvbt6+h
8SIOjqnHMwXMwSUmj6lLnM6qTiugXk7gtizai7MVnJrm6IwshLGrRQb0la3wGT7plBJwsk6TTl9/
0RsiQUyGoTbMMbPX2KzpeyHYGxJNRFDvJN+tPDYHRPEOVGs6v/cEpFQGo5ENAHTkj6XcVPuuEH2N
+Y4EdVZGugs/WwhicX/CJm48CYncKkECWD8hEUcDQlZdoD+v+NY58KvHH0Wi3/q9axI3mpjeTHT2
aX9PeFZTmKmHp5k7lSw9mJ8BDS9miA+t5fiM0meXLd8QRWmLN8QEj4QpHAjQqIFNsfB5v72Nl8K2
VvU+z18GH1bQ6Y1QwDr06m0DZVMBaGcbIDAWUi6248q22eNcw2dl/wdbD2SiLaWAjNg/EKALBK2b
cEfkSfMtKwyqPWUtOeYX/T5cfcY3Zwpxq0TC1uIe2aQwmqFM5ynGxdBWlo94rTkY0+XqoLUCDkPn
C0VvYnZQOwTWcDPD35Htvu/7j2V1i/1NxFmG4LrrMERouWZO6ASxPo9gBeLv7CLvVGIOUegWIt00
oEXMNgVfmDkxiy5sIocrSu0fcUKCpSr/h+ndDOsNv4XKTVFiF23xJP8haltg8Crlg2AjrXmOuynC
1D0M5k4B8knsnEBMRmdg/t+UpUFtzH3DWJnw2dz/y0r01ijD0YPl7ePyG8DFNqhcWAO+BGCLXd/H
j05teemj0UC0fIUkPRVbxt2z4p7MIl/cpjsJll05DKWWODw3rDK8eg2Zt7TBYyD1SBWONGazSOxJ
t0SjhF9T+u86lXMel6Bch0onna/ByEyxk9VhembIavJ0KRcEpef7Fs2xMTy4ZvtAwPHNF4gvgfhG
2tiGjPu/vCwT/UDxCkyLfeFI6dHz4Nbp0TEG6GsaSFs7ksxyQh9U7caJ5qmwCpoyDj6KPOLWwhkm
+sTQVOUcYJ8xs+J9KtlLuw3umYC0PYxih+QYOMPkRh592FfLa61IKG4LuEek2f6bQhjjmXDZAdjo
tq8bSqyDM/L1vDmIJUmGW8XhQtpQA0znXTpHwSinqQcemHAT9yOkVZBzE9b+kHZEmXomReDTE0c2
r3HtMoJSz3BENOlu7UTNq/SROYDB2+uATMoMxxIIms24/kb6um9xKnERV6BBnj9PeXf9+EaodOUJ
KqZq6AlJzFcAX3hVfCQhKID2ZQUuD5J0Ye35qOUDqslLVRKxvoJvPe64rgMQTfQDUVO0OtYDvzIY
nbR+/U8+0e6p2E8X5S0/e0uhr5lzL/plSADkQMtvMrCcGcTbvRqNTM4UPVxnhs7q1SwlqNRkaO+p
C9J9+oha9S7udfsVS2Rm4uWP7u+G+rcrdYOiUVu2uIZZ3NAAG+2zdzlpz7wBhjvAPQj4+BIvpJmO
rLnzCw6X6hrlxf6iRvPQbP/qf8y2Ce0XLqtJE3D5B5OqhFM1tfXMCDeEbyU4GMSuOt3IgyRuqlEg
tLAi9DRHCZWy4iBGTAwO1Tmt96JUTEV1sA0UXaBobBmcb5bBqyqdpju6ylTyBqGI76CkDq+aRpIp
7etvThiKUfAG9LH+YYBj5VDa5ktdHZ9iY1v3qeIRpx9Hn/8XI24QPyoaKF4LHRcA2PrmP0D7i6Lr
lb4rzbCpodnxqyySvmIoWla/SdHRIfT3mMg3HSwb0Pf7AI/1FHLtWL5PIJhxKqdCbAlxJt2lA/6U
UdsKDbi5kXaDVnAbBJiaiHmYRIzj3r5QmktApV5VinK8VcBiVEo7cDGlzgIt/A3ev4F7BAf0pV9M
5Og163jrDsK5SOpDS1pYcUz2iDY3w4rvwitbuoWDa0pR4WQyd6Z8iyA+4xtecITdXYMIn9Q2r1pr
0BxEbftXDCCze6oEeKx+DNPhOA1XjSKNw/BhfxN5emiD28dDLLqsjamth5Oz2H+doTbkZE1JWUbK
4sDBnhbmK+8aRWXNdNKQ+H/A305+k8k15HzG4ytjCMeONqua7DNLMb2ub8IZ/DHH94w00m49hJHa
ELwQl7fRSx8pvRUfOHyXcbHwX34rVAgXVJzZQD3XLv1d6qXZ391aAYpidP7YgU84r9TANMg6SxWo
UZCK0PHEsYigNzh3Q2EeOlryKPZ+t2tNg8A1AP8lJyXVZRv/OSJIRiXhEe0bjW1DFTK66yRiIZWD
SYcOaScdIlzxUolNHyNtEfqLS2LNjU+T0/ewaKZ1YQqEEEr8bkoY8icFZ+ZtMD2ivqbL8ZnGI8nY
wUrTBYE0IM3NGTgSWajcu1MBuFwwbde95rE7HUHmCfL4VZY3qISkFQ4vKyoiaJS/SMCUVFknzvoX
kohHRaoGWbPxxDgt33Xol8kS/duKNU9QnuvvLLOU0zY5nEz+BOEJMG7OR5P6jw0bjEfvYaZuKnAo
1kWFLuPue7IbA1kueRr46/PyXDiuGjfCG58BNxn71fqF09LdR3Agc9OuTpCcdtkoTP6SV4tJ6AJh
RH0nKrWv71Lo0SQqvlKIbpAJ0/4hlO+R3V8RJ9K6KG7JLeV3Pdg0Xw9yITyqJS39/d4vnDiYzMPn
eh8ycdfF/6/bMOdWS9J9fctOUaM/yMs2hC3xQ4/4RZVtsuTtbt5W+AsNGvRVP5LM2kNRXmG1927o
d3BpItyYFhxNNHicx02NwZYXQcphkBrMX3lO4wXMa+pnoVAHfqB1hIOJAzs15C1rNC2HuGQ94oIE
LGrL9nEv8xLac6LinTF8EK5QSYoPw9RRE64PdbiOEU7uhRFEPMfUtOfC1++jbXZcJ7Vzc6B4RJab
l7zugd3jmRY6Ide7vWlsVoZRhkWEwWcKmNE639fb2OMoDtUZJl2KS35kIekgkyGuP3BKwWDQbBnE
yHVUzOPCGYXVkBWj6cypzZ1fMvxV9jgobXmy1gqhugaQWh6RYuPdlJpwEso1gR6eP5os/csTrjah
zwemx97UL2Yms7JHCCIYmQwzgMI/OuQEGZXsSewHBaSCsem0VCQxuV/qLWdcT3er5PPquYyqxir9
XzvtOJt5QWCFJfwKoyKQfK+7kWtOQ1p7OfWFu07IafqlFTkcEi2W6BJuo1sEOsOMaIq0TChDaPKJ
1B0mxY1mu7+y9We8QdCHDmUEg2Tae5W1AV+KYTGiFCrqqv9MUgDnQfVZgTgZ0awhqUDWPJ2kIF8x
gh7sD2Xp8ub6eJvopuHfTMoCGXzntloWHg5Q1r6tHB7rSG/bmdUhWf9ISItPaK1sx2hIvdoroT5A
OrBLgaBIHS2UyfaaNPjrs6/7c72AvzwtWGFIjbBrqT1RqNNgpTKSc/LKhVrbsjC9Bf3QZMcMjK5W
JAq7TGJab5xQ4PXMUjC4x6dswS64dNcX9n057B2DPTrse4lZ952xXWicDACISbp+7WMCYkv1fKxL
xT8kAJBMMKi+GykKpBFid8bC90YJmxi2Wr8UUsj2KnuQ5P48oP2tdNNTdODz5oI5UXfolsxuLxMp
vKKFpIBvdIstxObatM5kwxgOZr4SOohNBZmHB54dVXsJi+2PuIrMnyAYxroQ8rTLz1NC8hu1pyvi
XBPiJL5OxSGLPbnz5fVI6Bi3A1M1c/MgTQdruOuyKIyGuj3AtrMG/lImX0Lqa7j13pC3pMbFcRT0
41g2zG8uN1GqF0gW/FDexgi1p9Vw75JcTCnZFQVnNkwOWSB6OsiuBliWHRAk/lxX+uBhq3rAGxdx
gep8Bh4iPyMvTvSYqm6+OwoEHuwsGbvYIOBGzQ79qg2D42HKokVIwSLJ0ZSu0nkBWMdW7AtzO2eb
+kv7/fecqDOayvTTismM2vuTMziT3a4ylZJkhgS2RAyty1mqa7WtfN+QdlkrUsKXs+1ztJj+0PaS
DC2h80ThsCnx/eddwgpdRW6tCX32gIJJAK+YHPwR9QStNlsCLg453AMWgRuCDYw1hza4mvtpHf8B
8P3zQH/cq2f6hZZE0z1XbySRuU1SzTZDuFo7mdeo636eY8HH3WVWhkE2tQEie7FmbUrncGsCXAlD
aMt1NNwyheohBkufyCmIBIsQ7MFEKBJr+gE2umUCB6NfX/UcUb/+fglLoJzY2LKg7kCgGXgujQIw
bktr4Xs1TA6V8h102yRYMA5PgnYsAxqzoGtGiq8z7bArnjoZcyadPzKbuIJYYeQAT7NPuwCZN6k2
w7GGPmRVorXwHlLvsdPxmX+VzjsaG7E3mnv7z5uul50FDkvZRGlF1qcFCqcDc6fkMam8Sjicaqoo
X3goX9zTWLZrAYkVVYHPZD4edN37T7Hz7adhXSx198YSXUtWJnCJEJacQr3uRokiJrLug0vFcDaY
+WfAyLxdceIO7a6kxc7jI2XsATYmZszdYPClnXo1nBETKWgjJYARoKRJ6hTQyDYcyErMThiu3sVC
ui+qGwZ1jkBFzIDAxb+jWL8csgRYNGOrbb5k2+kATtSwLTUIJcA6WNifKVKJY8TryLkjKdPDgwcq
HkjOqzd4Iq2VjrHLwQLmdaxFfFRGrgUbj/nhAWEPvWvdYnnrbE29kdZpxwUF1eYQJfWPZSsezlFj
IVOCU/ZizoGZDUYof9QahpYRLPiHCVNwv9SXSLhbyKYLOTs0ypFripK0JBaSGUmgcsj99CokTkXS
KDSPU6qH+VepIT5zBR4sc4qh7e1CC9JsTZvYZoI9CRTZqSMCQff3OKGoDFL8xCkFL0ft8F5MK62i
vSJoq7PQ+YjhQlhmRAM91qeddujMwBpUnT83kN/AxmBSjZ8FNvgqh7mK83xYQLWhRaS5mWuAaHne
GbZK5/vRlKtRamK+I1rpsCtL5s4dljDRLD1Gpj0t65NyDaLjLz5vQU/gFL4SNXAORr12Qk81jLyi
UVYTDJbAvcysN9UHrpRUXfRCAQW1RwGVqptrLBQp1btUU2g/7taf8+taHTOe3yEM09WDnRDKWR6g
5aN767G0Ww1Wwpe8RdPAuYdkF16nOu4fDxX33qk1aTiSuod+YRT9fgEsB3e8FxhrOhgEm4uYOQNP
VzR6CLbnMVPxTncSfDCgUXKe5II5O10WiHpUAe6Il8XAptXeT299Ro2/rDkcteEfni9wEvMMxq48
JyGxdox+/OOOYHWIzCbk8TNvuas9+7wRBUiIfPRvUt0pnI9lKnQUwCikIuLJFjkQAIkcGQA7r064
Se94s+SP4qT8CAZcbJYzVU/bcMVcA6/aKnJREItTZK/cNGkkO62GSBxlx1bXDqD1wPFa10nKMShy
tjm8+5c5Pc5IqVUK+UfKXzSEoRvhypPTwfWhUMWH6EePQZa1U5YQAem6Oa7Skg8BpC59UBJHtFZm
wOfq4m0Lxb0H6bM/7eOdHPhxPjuGEs3msA3EyWWTaFgHsRrUP1m67bjhTia5eWZoDxci1mDeY9NZ
RWarh9oSPHNZMewLBPKh8U33CNC3JtDUnOohjnpOF6mLekz9oLiHqvZ5csH1ZsjJYlDiaktOc390
K4ASPP0oXxbwa0qb3CgVdH+d485MWZSV6bTxyyJn/p+qfQULfY8ni+UcyQIiNyrTj2/hWjXsXoM4
hg1wav2qDgyy09y+gCq2nGjlhdsKtQbVrmT0Wm9BOr5CzPrav11/uNTEvIX3jQPqBWP+aE2ZcVPx
jXsGyms+ZHX6Va6mplC8wL2SCg9qgnPRPUCznWuTDVIMDyCScdFVw6hPvPGonMvCGySRLd0y63h1
/bfm3lFckdaUYFjol0p2pF63O/sN43Xs56znTzAn/XYkzfQNNj3QTLmUJxthMYzf1idxwSunjt+4
o1vY6KI7Jga1Q7r0RTWTaMroqT7GXo8Nr1y5WOG0dqLmRHvc8lnIxAi9nDVYtcRhKlQIuqScP+nB
jVQDTe64K4/UYCoYWLWpaETB8IQ1DVi+rclIvlJa3UiY0x+S8PbkX7Gt2BP6YV7eDc5Q1Hb2ggrw
MqK3cwwu4dG92QVTrbxz8l7nfjsOBxMsqyWhaFFqcnXsLKUJ6ZBdnTWouwcWeWnRpFPtISITOB5p
ReMkK38GfHez7oB9sVk7IKnwIEKG1PGi09VmmEnzaUWCWB8mAsA3l1kHvrxeiEeM0bRhl9IZo9ku
nMbluBnwtLzHYCE2eiXOQASixyEOBxqgTrlmCmj3NwDub8KGLIzu5PJAYYIxtN1h+twH0z1YckgQ
RfC/0EY9Cc2UTygKZxLJ+ZknSwX2JhO//M3GDd1UoLxO+Cl5tiMdxg+G0za5aheBme7Di6FrHAQM
eu6DM/XXQeRrNhafmXPCyMZ/AvW67o/nQ4/NTjGkJ3yVtE7jlr5T1r2yF6jO3Okbju3ghm6nVh1w
OXbM0MXhL+0DfoqBtMxXae4aPib57euwCpcVkgPDPyVVxWLXONvrx+imXywOyj3ltve3VZw8pOxs
rrAS5xKrg6zwxI/UyBWsQYfvccSncErKd0Rh0hDXfaII+TmiSkDG3iUqZFwyaYQx6NzZlZeJTELk
OargidHe4ac/GvLl8zJEaD7zMw1oBajBPA8+fgKkRlX/rpUSo6shK8Ate7BEfIPyOII+aSvNHBap
fUci/PUShkCajzTXaUz2wH/mfGvPeHJBzWArs+gn4z3aUWlsmDatEQCObJheC9wDIegsD2qWqQWL
tzw1mCaXg5y/0OHllvOh3pCoYchjJRYge8X/bou6YjFPUl6kpITCEoOXjgbONiX9SYneJ0jq6+zp
DUJfNd9pg75VUMqxPsUrUnZFdUpK3Iu44OWy28Mr4s6DRRoIWT0oi9CLHRlqT4wHC4/wpvIeEx9F
3hBORli+Ysalb+cjAs0vSo7V4okiiu60hM5SMy9nyupK3Nz0x8esPsfACrr1aC+bhfVYRFLV7ZEl
pgKOroYLlfHUC3pKXyskZMkqLq6OMkRhbmSmuNuKrHWpd/loFvC8IHocgCB+7cPtOMAtjFI220ic
docH8EUM77IueetC3M2MdksttR83cS2WuYhOni1jn7S5J37GT2qkY0iwDoJP1SDF698u5IU3Omt3
PLSERi2hzYgJTwjY9s+d+7UBe6gyBApwAMi+SCq5OWLrCNyPXdhfCMg4IYDIYxKedMlp5ykHPwWH
Mdpjc2DBWe2YaHrk0WG7hyebGZG4gluoDQfOs3kK0yXdpFE46BR/+0j5fyyoSaxC01uDyshujsTM
sLF3pK36UA/7sdje1l71gKPg0jWBGzhpvztKYJthtiTV5ZgVOoVSSi4e2AtKm7s7iIFATCiFYACy
cf10Zvj+Cj5HyR74l3DpKPL09AR4RnSDAtor0mywSCI/8H9aMiiU5GqUQ5y99Zp+zp8AFJyliZZl
bIoPhnp4BSJvkUikRoOiNRhC5iaNSwmzfoLLu8C9JKjrj/HhcBz2ey7RjcMdOZicWkxhDmdeo8no
ZUMfKXf7hPE0PIX8Lo5mtZ/AzlBoEIdyKaoXlAV80Xj/WrPpq1oJYhEgclnmMq6PEQ6iblHni9FW
07XcjHQT21h/rPsxiGxyJihijiuXDmCh+eGPV7NHXzRmqRZODbrjVAEAUtnEjiqBg8STXyhH1tru
pXF9CiT+IS3H+ecrRBFkaaFJt34Ef3rkeIbwxE1kFEd50qUEP4HWpoEWa72q830fmCn2mVrF+OFG
oiVTn0RwqdOO/nAB3bHOm60nARUjZPso1+E4ixZiD44v7bQT/NldYrdWngBYdXK1lbmo+8hwwkZ/
dzzmFpQs2Qx0L+wZyQxVx65JZ5XnDXLg3xEEzBvSTVeFbXQLAdmceTJW3aPgPVUGU9wgwZ5kezQQ
ha24Bxd3nGnHBglK/34HZhPmQDIHzySIRUe7qEQxddAZaUVSYFYosVBUdjSaNZf1SJDTyP0qq4nt
kpvRW69nahhU56bA5CySYw9SRJuJELHcvUO1nNpZSGODR4YWyyFfr8MHjHVymjLjGcVto0NhdZFE
KPOlwYOnbhsYbCjUK9g/TylQ20UTy8EO6r18b9NhzfCuHk6PuxMa9s3b35QNCmMVLa+zTLlOhV5G
u7IHqj6eSGvPZrlg3U6XpfQdv/1SbCHC5KCdR3aFVSowBQ4TPGcDlR632XDNwyHSF0SAJauNHJPn
ScrBkfqYbXeojjx6ur3ShQS7u3pmkTaeQOhCzF/ApElh+tkKlLDZu7wa1ELqqmBgbyWAtw9FYeOA
iubQQNnQd8bsW6RYXftI34wJlBbIWtNGDgN83zAhceoEpZG0p35FgPEmtDw7q0t4EBVlQbLgoFNN
WTCMs1L//q/v/nYt5ldWmYBEwfZOKpEZjURyPK9wSeBsx/DVhgx8qIKMUm7r9pdKbYBHVhWwlxmq
A0FVFemYb42c3TrR13mJG+Zn/pe5u5BuUXb05l3wAspPrn6rzEZRJR/VBNaq17S3hJfH3TyL2+BF
Hz3mOMU1OyqmxvCUhDd/TalV5iKOdA8pKKahagc7aTjW/l5qxIaNHfRNcIk3iw0aDj5TIOWqyYKu
NPDBddIDeVPRLqwqnGYejBXKbVgLxI3YbcwUopd3QQec2PNIMxNyJYKbG1uJSpopLwlFzd5+d0Oa
f/GTb4doTfPyxfycfn4JiFtAF1H3HILnWRX72ushnQZ17mBG701rn9NrmmJiV8g/xRWcUob51Ufv
oaQj/rF76hDtLDnTskfXVkYGsaLIcW7X3IK3WUIwI8c2Fmg2Z2LzYtjMrGycW9q23ovJM0HFif7U
MgaHcKSVGmnQyOZSt0rDX/Z0vWAJ/orQgHUtHgcm4hn3iEF0rN32Go3H5fKALfynd9ebzAPfcSUu
Xm0SMgY9UYK88PllJJ2djxbIVMZmP+Cp06TjfpYirUg4myOwLCl2ctXWh+OcBReJJC+D/3hhfWpz
N9UeEi2oeXqFYXfJsUNfnmtIz/YFkOYnzRWXlmdmpB0TY/ijs4eEEIeVqXnyAy3sqogPtZdVMTHX
2k7KfnzxL4sFXk/o2BfuPVF4LAZa2r1r9rFbUm4+phP6mpRghiQDBVNBOHa/ookgnLLtrt0c7WiS
ECe6/WnP8sC69rr1KhSpSLai9b8hFduWMJ2vankv+/6c0dldQEiNvtZoL+8JvadfrBTwhRvYiA+7
Xl08mSaCiEd4e7Oc1wfK/Ue3yzYUiHEB975thG6wS+G6lm+eV1sl3al16L5KCH8bZ7Sk02ibKrqG
wQHwlj6DgMGSfOSHlM85wcathZk7w77szHtsz0BbM1rASkkACyUGR2wZ2Crwze3OIbTnh8Aj7e0l
Y0vYU0K7oC9dVIiMLsl7jw9rWmc5/Y+JnoP6qoEhoDjZGx/Z7ihtlKlkj8gR/SpY+C9gaSO7QoFL
KyagNLtpC3+whKawiRWmNUjPohxyv5VYO+h0ht2pczwMKkiXTNjNzmYmILcuD6X8Eo2wHewRdciJ
hK7sBbY4TRUitkTl4xuyrrrnvms2xmzkQQhyFKBcXLOXplxy8UNXJTIUitgXFHZHpWCdeT6hJ8zN
2pimiHH/XQdy50CuwfPqKMMPLXA0Kgxwyarqjqlo0OVyLlszF5CaPSDshuaf3KL7CImroIY1MEbu
Jq3peqr4rNN9+j+pQtaTWym7+6blhXkE71AlykRQLd3EQYa1+l0Q2lmsEcbm2iy3q2D5OaMv8CA3
sqkCg4sOGaFl6C74dBUHY5d9oaQw8R4NonBR6w5wnaB/q9k3kbrTMpHEbLEYRBTxXs78N1zImr2E
MbKH0pebz+vbtYV3D3GnTZYrlT6gt14lodcuG0xcgq4aZActFAUKcolYo7rQB5GVhctvRyc7bCxY
pMRydnx7dkFrcSc47WKKt2MVdZ8AwEmcUTwQK+nX71IsOSnA5qQFd5AbDJdVJZX5Mc9OL6g+P75W
Ytz7aZ5BUI6zdTPk6Pm5LVbAFhKbYgOCbSb9KDMyFHvBqWx8E7PgLm5eGADtPbl8ss19pYHqLD83
ui/k+oSIlrvI0lPI14BQpql2a4u0O2DOgyPtfFcB8qffvCwt+VXyhCH27otoin+c8pLheSPR2OcP
wh88vHNbZOs9NSaY/wofm0ZSLGYH8O+ZVKJcW60osqMm3aAdY/pS4t2TiQKVJYYMrgoSZZrXUOgb
3Wo3yjXqsBqVF7vK3MNyYpj8MRT+9r7zosO1UqiDZ9/gPWj0wLX7e+TLeyQ+MyUqwL9SDvh+wmHZ
ZVy6Xy3tM9nuxVuYbvmHtGqxy4OlxCW3IcDd4Pxorlz11L3jUJm3ZSbXR0Es1iS1uqmro/4xUEDD
UlfxhQiWh9gQMkHiObibj9wD3hR3SsdT2CRG9w95Fou7wc4LXaDxtkQn0oVoN5wtVDLbSQ07UFJx
p/CfZ5fOKrB05ZtjcqrivDWAohQJu3CU1Mwo/tI+T5dSFHAQCP9titaWhvbwbCjHfigzTF79ormW
FLOCuSNKDma4ZLR99HDoF8AI+JGpB0J1Ck74crBCw7/9saI5NdiSl2ky14rTDy6BWIL+sRLyze/L
/CVl2OaNULVwKHZ3bPCekdB5jbhOQpOloG/h32Gw9REUU78dQz9hgn+ZVhyS424p5WR8DJBHonap
XQ0g2dVZRR2Hy3XiU98DkZpwIAHsOYplycObaNXhdWSyrQpzXZaHuER0xFq7CF5tfR+bf3cGDzCj
sMA0PoujG9dG00JXt+YRqIYxUYdmvUc3TtWsrr+uCF2NVisKDHj+2RnjF1YrhoJYLcAHTtSFLGUq
CtPXKURP0mizwe5AlV544I9iuw4K1FjIf8Z8qYybLonL8vOb2uqSLD3ncLLgjzcvokWv/bGYhyIy
YCotHlAqaAPsetDgmgprg1+jVRuFFbyOzagYwsfAC5WoKWdZ9qDhE6X79xe1G5wTva69b0WLU/9W
Gvqp/eVLC6xUHx4r9t6SSGgX3iYPIX50a+S9gSgSAlQLdm6qzjLdLHP5f1Iul6gYlAjLxrwk5PN9
EYdOnfUXbCdsfcUMdh0FyRugSZkTW/anD2rizDNEOu7V0lXR+r6ejtKnc1aThnmFN4hk5cvt+Qu4
gGEvwlEiXxPPKvdo4MMc9pns6ZBlwHuphklYSkNEZ+EeN7My3MHHao5mSv9FpEX26+E7HJ5Cvs9Y
kpBeQdWLyjpcyz3FZhaO6A26HrajX69YdpPPtL+EfcqhQcd5QpB5jekJ4MSCh7cAdaSs/XTohcTt
VwUIY9i28/+QXHeubfOeRJO+q2hUb4CYhTBPh8A6jQ5jaL40huHvUo2JDElRrx04avBf03EFrXKV
WIPgMT+soK+JXjCaNtoezqyg6r0vwZZx8qJZYsb3fNR6+ZnEf52vLr0QiRSdgofEgUstOoRwCYI1
oD67SY09RrLjs/FZ+riLFtxCYwgg101ikVvQvth2Sf1dP0ltNk/c/hHiA6LEbesCQ+5tkVnuv/L+
NNRJhfAOgHxPIFZClsdYsi/GAuIijQSoY5mTihwkljsbNHylJBKfSovHynnqdLX72xKbx44+JwVx
UhTiDicPkNbLb+7SjDGhT7KqRU1Zy+nG/sPw7PeN2nLMDo4ndiuSEpYbmoyb8bAunJjaWHUP7zJC
dhy1hU6EXEodj0+1prYqYtWJ1wpDWbwOeb6emmkV870Z2lvGxi9j/vmyjO+HUbpoS0Q58zV9SF7i
0QpzCnMB95Dw4nd5JSCTZIMuFt5ExyiEHJhSE2oqH/XHryHeJyjwnXwZ/Hf6peDJ2ADOiOy+WYFU
9GUpj+9hyzNbNQlC1tbTxDz524KzcKX4CwvZNOVuGoSBP0hpq9tw2FDq3caIQxSxa4pjlwJVeYwT
fRk15blkD/Yb0f9qfD4dG6vNs8kiHq4hmMEDCV1ExhSUmqzct83Mp+ps32/d4cu2nqLYzXwx4Q9/
wTfpTebv1ilr77FRjMCOdc2RYgeaqtPjsyv9MlIwtenIVDE+oR67/FGEapQmZmpfQo1bEFBwwfQK
7pdzTMfH5l7hxSS/tkjvG3au4JQdM2Tik9YkXrCadLMXrLS2OeGXa+IOeob4rAr+0VK3wowZe5ot
Xgt/lAflsmVV9OTberwmI1OhuL4Hw0+TZca5AOiZm1ik2359JkwKBTNoi98URx7GEaMBRNOxiE+V
L3fTvRBcZp77Oddzxhji01PbLbyuTXGn4JTY723yHHiy5H1eY1EQCMP8YbJza8E8VkqonJpOOb5l
MItLSRKSHY2oR0eMXagvRmvW13VeiFPXQ0/zETrZIo1P3gDBbIOuxCRIvLFDiy6dgkNd8vxEf5UP
8PUvTrgEl7WGpZVgeWkLBlkeq1nshG2V0ZOO5cSGjfltZa8l7i303r7nQP4Jn4JOWODHKLEiqMb1
yVuurlBaVYfYNRuu7V1+PZQ9FdraGnFTtOu5oG715WKKUwSTYfIRq/hZbKkdPXEljp3Q0PfsoniY
MbTtXElz4jsHdLPTeC5flMoQV3JGs4rPuM0FAR/B1t47VdEDiOOfJj/j4p8u3tNnGU/05qXnHf5G
KcaLn2eVX9J0J1eXUEnjNpi/z4RV3pu8Qxa8HzbvUGSoz/Fl07EL1i268FXdWMNR5RWLt+bdYR/O
FpwWN2JSon5KuBvCtw8Os7377yJ4ecVNJWCy0T2kcYch+wXBDHjZ8Xy2FBwaMoiiMkXsvxz0jkxQ
tGrvN6BJWiG0Zne+56c6m4393Dbt/CKRydX4zLyTrhyMJ4fRGnaIcW5IIAZNceDCvb8Gc5eOv4bT
eIZGLzvE9eVEnmxzO52TisaTOgtrJg0ESeGGmEsOsnaGs1jsSUj28LOIz5X3+69C2IBCWDxam+fF
Opmd8yEHcgoO59IPUQMl6n2nPd8v2EZPIfpoWTXIsZ1yGS0BlH76NalC3cX0AIRW4OOlKXaMMh+X
tdCkOPKJr1c8UeGMsGV3jOArmVW8eNpmuSv2pqExj7YyhqilShFFTajaDDplPUg3b0/c4g56pgac
qD9FIkecTx+i9rmp/Vu5GaB5yh1SwjkPKa2KLXmSHVQ6d3jCh/GUAwv1ehtkMApMFsvcvyE7Q1qN
mfKVIw94E1Zt2QHU1ffHJ3nBxnd3i4nOVdjYrLJlSn7FEueeCDw708qAby7+oc+KIbJ9kJasZY2Z
6ME0oYzkCUggyDtXNAewLpDPqXTTt3TbKlmOiJM5UnAVPn+H4a5YCivi3aN/iFxpAN889xKTNbNS
poFSZWInxLbl6DhXxocNzYTFAoI1NQZvRegq8uqCWBJLF5XY0H0z/2pXrAexCD1q/lto7z79Q2Nv
6+jir4ZTJ8TWG8714fviJr3Zb/XK6tLBxqzIAwlFFbw8cXNil0/lA1JXCq6J/51OBRVxtYSu1nqe
DM5/BJf+mswQmHR98NESqH1EqzbclNTS9o+LKzce+kY0I3W2Py0+O3zitdCar3NGMO34jLoo9HU3
zS3LfSi7QRlENpnN7i+BC3u9D3d9mTtfWFtK2irbNtrlJ0/fjKmeCY6GnMBB8M4XKOzs7bAWdWjX
h4xlJJ4hsrTuexQ1/VpysTr421r/QCtQr+MNuEzVfL/NmZ7VC32iZeY+8QLQXuc231A+0XEypx0y
xc+2F/pzg/f2szJA22MEr1LJpAP3StVL39YBYsq6BwCslfipY/l1aAcCa6XPYHBE5baEyz7G+DMA
do3fpgjCu34l6GytBnL/0Cu46u83ruJUzG+r0JyRNtm9VZ0XtibXaZUmk0tSoAkfP5gi+AdSQq6V
5C4001YkpOMRL6qTR4Eg77/1lMjzPMCFtZbYSUnOI6RVUbd/mGlTYsvvpRKCN2ODGoHL3DlGincj
lv/CWZA4kmr33I3LCVC1HuolrGV5gHNeMZI11Vaw7PGWceAk6h1ll2mo5TqI4furSSbVLmqqHGgV
5XSq6Cb0amVGC6NQ13Of142LrNXiRy+qDPFedhafbv9YkJOCa1tkUybvYmWmMRn9STbuqfgGlyTo
XDZKi/ChfSSP5g1TKSdp7yXe8VBgDYEhj5EWoN6BC+N6MzhfaaDTRk74gH6ihXoZ3PAqu114ETPP
JIcMa9TPsvaI8973s6Tytd9yRdU6NOhbcZzPyYXyCwlkwm6f+6UW6z71tQaVvTLpgI7HRn8xdpu7
obH0rhVQkmzzOljEGbCwW7FBd+Gu0oB95spOJz3+7JtTW8ZtsTAF4N6RxFwFBOrbbKctgYPomzI8
RSNhSnDsPg6PZb2ZV07Ef/g7vugkDVdtM19pnFmvvHy8ccIamm+ItEJPhVBqxLVRX5Jwv+pfxDWj
tmH0oNEwo494kXzpOm+0PDQm12YJBoRok8HOGsgkZ4fhhyEknCHgpZ4FNUPUmGkBztaSmqxYLry3
WFcuaZ/ntZEjf/OhgxQamq07jSt/+FFCWzRo/TY0+Rx+kEwcUdoxJpAbCwnopsr/Xcv6Lh6RvDL5
WlGPMys+jNCa0TPYwJ71z8xwi3wFIjz870OtTLukGVwjAovBl8vCQGXUhIHtgktO3z7r3I1QgiYi
CxcNQe2rSWuvAbRuWxCaX83+FuyD9ef4IbcySfv4JuxkSVD0cbB/VoowROvQAvQG7nmDExZLS43E
+QJfc9NPSrQNTBCa9AVHQtgcmArDYPMWaOJ4sFVqYQXHGORjEdHQU0k4UwE4XMHhkwtmmiMFn7Sn
1oRojv4DgzAeFqXEeGfitgIkFwzPPUfQnrJBI6UK1q59NZ3vnCYnfjzkWsbGcKgK6qalV2C7R96r
wfc9OE2iaWKmrl9AX/IGUofXepVPmDyPxwljRWYmmexdo+WtwLuV9Lk4u5M1td1c6rm4edp7yx9m
DWefey/gsR+BRrLqAVSvtCHJ4ff0U7bX1ooOHjCMh1rsvrwOJguTveh4DCHltKW3e+c0IHBm6in9
Pc1Wcqb6fGcm7zpPAfp9ssrnq5dqQNyq4qqs58ySNlmCUyz7le05MusConN2YUzLg2I1M06+GBGf
Cz51fY3O3v6AMQHtIQglxEDC8rrENLxO/IG4CFWdFUjN9x8PULEl71XM1R9+ER1aQIafGC+2jCIN
fKU6+/jz8dm7jIgDkPTgCGfS46gNQqe2pMNjch1DzJwZQpXYpqSJ2bVR4OZ1GXvD42owyVVV6y4h
fu5JejjRRKXhRmxDy2uAsnysBnq4h3rq8512vJUQmI79VgLQV199e0HGaLxyzfEsul5E4YV3rAB0
vrIXiX6XWVzWi7upJtqWK0ho+S7Unls3UofFJzutCIBhNkhdZvpndDGn6M9vIHp+DpAbi2GK9JSs
ZgtOQ54dkPZF9hNTMAIN9oVEEENW8Y0Xi+oTkzZBR2dDGZSyJABoxG/6w7PHy9U2LA60ATeq7zi4
QB+Co72EdWrABRSRK4avuWbvIJkvzpooRb8s96fUbcbH34rUl3005XNWOPFlrRwK2w4ZBHFdHAmq
k5VCIIQi2DJTIVPCVkXQWUBviVytn9shu+Xh7pLGo0T2X0ddmp5NRbXTu4Txym0whz1H/GojZc7Q
mF7bXkFfxkrPNNm1+e0h8ujgbzcc8rgJxRH1c+rzi1gMbWpTY5oQR02VpePRuc9/gwkG9SoDA7m0
OtaOzvozMvHztpus7lMOLnr3bSzUJ1xhHF6r4qgHJF4D3POrWju5DlOMOSINh4T9jiwmMcP4OtT7
tXl3SQ02ezYzAjLL6Hz/eTX1kaT1Tbz9OvszrNqjmmA4QKMxHn0JG2PF3L3IEgDabC/3jsAoNgbO
Bnd2pWKZ0nlvC46sT24KboSW+kVvKqyrsv3UiI+dCMOdl03Jfu35d+Sjo3uVNHXNbymgjzKdk8PM
3IWASVJPVBMkLsrHRvA4/++LbFFQs3A7zhfuOX0CxnikM+gVXD5meVf31Yke7FammUcYw+aowp9u
4/lvjMsqWKtWZFuRDi98F+hxa3nZdk5onjaa9ER4PEqVkbxQsNGIG4fQ2wz4YhANEBdB0cNBI7+U
0+yCUasih8SOalwPuoUR66MPCkFOV069vA8+RJame+PBkfEdYbJcJuvEkSmthWcs4jsiis+OWa0S
zJ4KHGr0efcusON25J7UUpsMUppNZe3WYdDv6fNsGXOrPWoN3gFEgwsUxWd1qN9hiI2ZuTdq4nTD
KamrlLCdEmxr0zwwiGgBAqm7H5A7BNF70DWZtZf8XCPKkrW+13xU0Gbw7hKbf3j8SaxxEeZDGiNF
SCm526UU/O29OvlntfOmtqAxc0HtXuaFxa79yiXDytNF9DJgTyIEKZhjSOmorFVf8w/2VV43KveP
L1qllmI8EKAiMhSjYZqiFu6CmbvM7HAgpE+CR9vrIFbpvq7F4XxPdPqEXS03ie0TNDPedfOhgH+L
ho80w37rC4vMLK109w/RN1nrxTT2jdr9+AfZ3Gj6u7E8fq9XNqJ6C+zTKGOR2x6WqEPBC5zKrpmM
d1/Cb5jkjA1I62tCrUIJIdFln43r3X7e9oh9Ywo4oD3b5ALfw4p4C8ytZ0Txz3tvfbaMzfB251PU
j6lmbQJrDaucnVBDr4YQBEwZ/kQnX7aDPjj0nYvgwT5wQAvjwgpWoIMccmm97IrKLAkQSsdjbtSx
WxiytguHU2QvViFCwLfLarjpFZFMgQPupsydsY0InOrrwOLdgQMkdaYGZIDayUHn3akWWGAMwP57
IT2HYhNbmjApSNK5EvfUR4G8lA8vpWrYhlo4mm+iK4DS8iXoMyPuaEqZP3Ik+6g8BFOCJc/+S8I7
xNWBzF0qMFRyNONZ2k/3mHbi/jNVN9vDPBbBA8i3KRFzetfYcYuj0TqQSxejBJqOwIdBOscVjopE
v+n90O5eEft9c/dJzBsM361oaHVvmTxmAoeCsqgQO68kKZ9mkImWrhWBDXTsJlEHWeR0If5hsNKp
crYsvbGopn9oAxoiizSsi2p5thFIEFHCbI2JAFj+tfstjX3wzXYX3YiHUfgOdqEUS+ItGs7KzMgT
WeHVoSrOSuoWsZwVE92F26x9uvaV8WA0NYu82nuneUZ7++De0ca+VOY0lso/Xo39RMEJPKAESNMa
Xv74i0hqtCbCx28z3AnZCHTFYqAtgy/A+l4/oVZKFgj6NuCxiuuG4KBYZpPrNMPkGXK9OUpZzC1u
mlmbBtBN3MYYomqC+sHGsaZCkA0WUQPCRQ878/tv6hdlAaXnnhk59en1r8qGZS2NqcMQbgxERcR1
LPKl3X7jE/Mdu/BfiPS/RDdNR1RjV8ZC2KF3+FDC1Of1SXBSX+AP3k2Td/yMeN+G2/yW6OUMZJ2+
vMOmiEI0rT+LZEY8okv/Uez5tn9u5jZfpFAxE9JC4BnAqgrufJzHdnFGiHUCNI8vMDA7i3PyDf+B
do4PMGh38lWid9YfxEyncE11F1+vqpZpivBC1o7gO7RcPbTXMM25vNNgcMPc2opH2vbfk4OZmK1I
nMrlXOGsX6ULjdgTe4EzQEPYypaSL79YM/MYNH0B5MRXTDocuLCQe6ojvpRAP+Ht/dBb98YoxKgd
Plc/RZKeDKPZhlEUThJoeAqV/OqJTLiUUd+gzveZOsp7RWDczvhJGpxRGw8sFzNzXvJGV9FgefJX
kzsc231kkzCLJhlj/dBAg1Gd6IMk542sIAXTws3b5pIqP6SWUKeNPwDapf8NME9r79+UjILj5giN
bGmzz/mmW6tNTqSR5PPMXs1Gxc8LqdrI0pBNET1mzog9CeCDEgkUsE3Eg80orJwFu9IlsMfSSPvT
CvEnzz4suJwq3cAEem0QauSV5VWERPcx41oCra390wNCNhyq5O87WbVShc7N1uFeXIX0DdR8bnin
pOEB4AkdTuXldGLFzep4f8RUsXT73cks/y3Xv3IfhuMSnDkIt8jcjt+n5GoxLskT4Y6znXaxocmk
d7pTh6QXlcbRutYXvN7vIssIoGY9QdTmrDaF8z9z3zvx/sEge0w4+BUIQBeley86y8pjf3OFBbTA
8uU1GzcLI1EOP9GYOBYIUF9eyb0l0TqLEDZLlppB2Z+Je3/xjNss1LAS9u/4HgkcuduhU3KwgvxU
B6jXZRbHkgr+zoij+uYBrB/51s032B4LMTuubqwo1WGzvMmMV5LFshPIZocFSqduD3qMTE4d0Dr9
REx6ORm3vOm1H56ttkdwiq3DPplbDuxHZppHSZo/Ruj6OyzX/w70NFztZWcvHaoFSzNQAoZhhAyN
gwVgjn/yMli8joL43RquLMFMNAVsUFMQ1utc3J+hRtOyKJ2Nwailj61D6inr8sLwVjH3smlbpRZc
S9JkfGVXnRszSRjkXupZ9hOEvk/K8R1YQG7BSMMSz54DaM6KoqTa2Zbnsw7L8I/BUxr+l+HIDyCf
TTkySHg1Z18HzrA+ZXvcD+UIBV7W1J2tqLb9PHHat13eLkhrdUCTLkLmNKdD1D6ydkixDrymWPSE
UPaXqrjlrLhL4OeobBb0lztU8AOvRhbXWLwHxuJP06u/Yp3oaBq0qVExiCHmRJr0PuZXDKFptfx6
OCJfoowQX6tFf3zSBX4YgcffhV7EcumnEEnQVlMTOI6m+NoydypHZGp2wV3YZtfTC0eK0QOyG1y5
xK8S+LpKEeDBIrkYCby654ReoIv9ZTtTg/yIGm3FqOBUSyy4MxoDSXl5NvopSpNP1ZXo4TiHHdc4
LR7+rzHGO7/PIavdrARi3LaqgWyA93+gAsjrta6dbo+oW9aJ3xzfNzCXnU468VULOImfVze80kul
H0XDOWDnnaPjeeEbGtFadOmzHb+poT6hIxFEauhH+uN44yr1EzF3ZL1I7XJS1d501hPVSHzKyrju
kIkirrPFsayoNcDv7PRq6k3SXRjSyKuS1lY2OXo2cym8FghX8MN2N1bxhSk3VGpcH6ra+BixoPsY
9INOQBL5uE49iVxeXPexot+AM1i7OX1YmsZKQBAVKPzDsh9gQq5TLm9mofxQ6VaCRWEtiF+XPZds
I35PsvYmxIr2z8eMbaCrYDzWCSXycqR8m24drXRbZ8o1SYYgTDeJOlK6dVg06c6uWecR+L0uXxM7
X8acCFZZRp+hWxaxS/uXU2YVfigCl83v6qfyEpt9LmtdAMYzU/wlzD26WspWE2UV8dJQL/97k+3l
WTyhtj9ZpVgM0yhg05s+DGAd0l0BWswX44YRPTRXY4+Nd8Q/+bzmwPUfFE9a0mbytrmViItfMvVH
KcL+t2v+Cc6oFBFTYukYlGFDGsaZcNm+sKeCh51LbKswzTLvnHcVITKMSXX6znwwfqJTzeLH8XP9
VK+3XJLfvbPe1phBpqBV30+f26SELz8EwLBUmErgUJUq4vvRtwXMZo9cZgMSGLM0TvYZRQoEwJaX
hyDrrcURPvIrrn98xgat/dDG4Ctx1Pv8MqNw7FRBKwOUi4lfed2h4szQ8yvNWuoqiR90IQnVPGDn
TE4gsbxq7dUDmSq4TloRhgi6hoefuDMfUGh89I1pJ+qAVCq8+vcZTibxdXEjiaKA8bq3RIpI4EMB
KI1RofEbip7tjpmlBHeGCoOSRyMj3c1Wa2BI34yhVnaqXtXanc5JA1gNCs6btRPJlTpgI4MqAVTO
pPr56DRAU5VArxYBylRwW9h0JnV1KmT3nZz5aleT5gwzU4tSbmYMwNxozLcATxG86NGOyW2YXpdR
s4w0UC/h3rF8OGT5EU9mPjdr5x/qyAgkAd+uO/8UZZGQbQUkcExtJRCUQIYFOqD2jGNHtSZM7Jla
0Q7dJXaUPyrs52L7sDbopAt6nz2iZRV8yOjxFB7fRpraD4//RRIgpPH4j9GRZIQ8BLFmhdBCvVVG
4euLg+tv7uFB71K3liy2RPnO74Fyv5+LkDYBJDxNa502dHcqPKrEYeZoSUr1CtLWGbt7ucDkwsox
MuQEajcehVmvfl1Bf19GXQSOnyjTxELhUvjNG4SR7gpwvpd449ntRmMO4eYoGrCvK3JFpxR4HMv3
ECne1e1LV6PgfLIkG4qxzkfN4Bdb83LkkZaEM4gsCFJatZfxCTOucETTYi0ZwxrdfmE//bW9da0t
OL2P7y4f0DMK29dQat6c6Zx4BF24QRxdBSGKELQDPzjPFFohwyLh6F2B23WguZndOSHPKsxgy+ef
dHgsrIx3VBm2q33ytnFw7WIiGfpdxBPD/W8ZCy2cmW/leBM4g2KNlk84JZt/SNKMnCWXiVerKnrB
9jMeizr45PIa9oasCJKEi9xtG9dtGbAvaVb8SzuEE4pYgi44caGI5+2OF7Jzrc3FrXkDq4ThwwoW
614O2cxOwCHdoAe54yRvvnycZMe3LJeyy/8HapwtTtQ3bF5vsa5qGxiXaa4d5KduwFlt4czuA3FV
rHMWBJtxVSnVPb51w/X7khE2vPyqXABKnDx3Qv75lcr8tqG30C1W7sbwbp/FJvY5Hz/u/lqfj5D9
80tCFjdXJHeH1krOLU0dtjnk290S9caqHH03cBviRAliJDlCeh7vrVsxpkH9Rud8DV1gaILBXgL/
yfa35rgNvISru8BwDf/OTk7Z3+JphjQG3NXZnxrwLIN9YjEO2nvxjCdZCHbqXdoRIan/3c4NkOV7
AD6shApPQm+8csXp4FFoaTrWUim20+hRtzikN269Fi3LLKUvma2HmXj68a0yIW6EarMGfEC/jIew
M7Lb6ym3MaIuIV4buYnASBdaElFsc8d3FrdJFL5fp72SwEsjD9YANRqFxNmy5WBFRH8jKmyJM7Pd
X7n4E0HbvsFpCqLe8ewvvf6v2VhZd2ikB2HfVyw5E8TXxAnvMojfX8hdxsVl3C0dam/8DdOQEg48
cT3tNXOH/+FkeSZ6qmWAxnmjMJfT6Ol+Zr//imxQKxYljwf+H5vz7SZQd8aj6YP0JjqpRDUGSwX2
m6/oI19Vdvqu1G8GOvx+8yCU2+00on1MPfGYInGEODr3229CfVI3nTmSa5HsFRNUVnINIzBtmbpk
TP6f50ijBJvpRM5sEV7wqcRMqoOQxnSnEbT/zQNDvfrKl3/MeeEMacgio0Rkx3SkV5FSYGYi9uhW
r/GZnU6T25KSBUK3l0PMZE/c3X3Ln1JalnY6Cd9B8zHC83pPNL/m4b/TtGzsqQ84mSd7GJxE8F2F
0iK7BmK1hunP1fJjSnaGa9grky/LCNle0VbUFP1dF5BWfFZa9YstzmFzKWqYeCqr9KJJI8nPKI5/
Lf0uZ7LZW1/bfU7Q0zw/pwwik7bU6IcFSQCTO+GcXesa3SI1vFjfwBRpy1JYE8le9Fpyoeiu/7El
BsDAWAWMAUMbuiFsJWUcNkKx5FG1cOhAwWna8jF97eZptEVq5LJK0YD/K7bTyxvo1kqXOZrQLxop
QGi4jTpFqWfeiHeHepjiU3bS4IZYW3zKNd5ztJ0WR2Y6yGy0WgWyqR+OJvqI4REZxH83P89vL/Xy
CgVExpKUE8ZTI+sBzySm8gA4IQ24esG7B/VVbNr+AoMeqhLJrwcqntLOqXQT09ZW8qkm22RTs1mm
JNmEV0RkTYXPlSRSECovJ6GzY0xp7xpJ/xc/PCHr1gaV8QhQPGK+fN/10ZZDgw3n7yEOcGRwFwRS
ofTzNcvUM00ac2f0DV3VLdYbIaB0D2d10d63bsN+J9ytpAdLs8+UL7OaJJzBxPR8KnAQ4Xy01cVB
C6UPt97TmKJveDSkHmc2QX26Q7oJCJ7mejtH0qldNRg4A7sy4zULn0xAkODGtvwhStPSNWHmTdYo
Bh8RjiApKnQ9JA1DlDPlr+3QJJEfL5MKeuVrorGcuwePFby3Jh0ank+41by75unxE3W47PBhsuJf
HkScaqxid7DLxAYuC3w6NR7MQtKsb7w1wb1xUA0vtWr4f9a7WkSI6AxMWQXgVK2LyoDqkGmbVaOU
41mhO5nCQl96AW4BPOoB7dnebc1Xi7Idd8SF4pSUrXIiIG6edDO8nHJVbhn8aCq0hfPLvKKM30Rl
2CJG9k0zliaIZDdWLC1yFHmkJaVQSfUhX/KADJZAAr5qBagCsDVB9VnqGFOVp/3JGOOvyyVl4gWO
qM8xO/REGcuogkDG8aXVmKbGrcAH806sUQga4s71gekrXvozhjwvkzQD7C6gauf2W11mIl2V39mO
NbVHCBhtWi2cue05qO8x19C1uGTEjopMGxGh32mezmPv0K7idrbWXA4hOL9FXL/iodZZZqjGlCBH
fK40wlmjJzyyqU4HfPoIlv78JlcEo+f4eDjzTwXwnKuxtLFDtU+UkWs4M3aRxoFi7ZTAyzCrCL0u
ppbfwL50mSL5l/emMT6IKvc0UZbpgwtEC2JjGydt3lCCskxUslMNxWAwK4Y7feWMnRyAIIUFSB9h
Rxgo4sNujxAqC9IthvMkkQWM1vMk9d9UgKOW5+A4KL8xZTYqYFA2ISSeAezdNea2LtuJsPNdiUY0
vkbEC82QvhJhMQna6xcKgh408JtjhiSSOVpYm6SuuurKrwRiu4U+DcqRHBeiaIy5TOwIL6wEn7oO
3GEPuvNoUZcbcxi9sOoRMS4KnaZquCiWlCuZwSUBmN9TL15nyvqi9xY/8aMCbCokBiNsejKo7ouo
jf+bIAMO/F2ANIAffXgzWeRC927isXHfzZ70ibGEY9yh/7XIpvr0GsEmxEWnPHqYL+etIPNALRoR
vNzU/G+swyIxfnweWwA5Xk1/gf5695rY/V1nc5XuQTjjzBY8RsTzoPI2QC4JHVZVfAJQaLHKhnM0
mvaAv3Mt6rqnDp2/g5Jt6PiClC4kUGd8eZOiZnl7bsahNO0d/af/msc7AUZnRGN9/NFE1hQT2GqW
NZhooN8hC6hiJ0Ar0MfxmSX7lkfHac1oTt+q6l8FsngfsWT8QmffcqsyYQzmvQUMx+alKoz6f3nD
U/YcJIVrhWM1X57rcXq6AwQl2GEMtn1/we0oYukKYNhNrYZ4tT9Ls9DifmzO11WN0gOaGFxRuXpX
mApb5sWOGjN7WKIEvJnnkGDNylLWunOV93bLHnEZOa/oPl9hF9Z1/B3VBEHp86RS9BJH3gF0lctg
hJuOsgUF04NG0LEHEoAjF2IRj0sIr2IBD8RnKRG+8fMdKYfX326A8k8ZyIq9oP6qMLbL5pP0HQZw
1AN2b+wt5h3OTzEtXCKW9Ir7c2AeyqS6TfHZnvvigC23VwtkqI5GV/6zdGYyQQwsXL0IIvJe2DeR
2s6evxfWZ+dawqofiGhSYhsz4TXmwj+lkx/cXwkdasP3hD6x+NMPIQRhIwvw6q95PFYBhyyriRag
500EzrhD//mhYG2SvccR01D1LAAOIonzT1gJmNsLTTsXqdpiNm2ns+gAPTSoR4mqZ/+dgWKT0ehc
1I3CPuDAZCVQdmK0g73pTka6bQTqz12d/SiMQAg58F2K2muOqro09hzwEzmgBF9mUsZRe6qr/+pl
jAfqbM+TgIaf0jsR0tYxQZwYpJeFOdJa1+woeYt05Bf1URkCMjuRSjNBuykxeczInoNtWwts0xsJ
xDERztiWqVCAeJKITLEsJhP/MZF6giZ2T7/M3Hm6yU2xE4l1nphoJ3wtSfHc9oMTAoxre8tpYiFr
Eotv4HRDKswTQokm/3IOisr53GvpLZLLDydHXN3gFmWsSJfGi2UwpQPnYvlV+/pDnw6PnxscAuaT
5H49nyCdkURDyAFgJjLhwHrN8cyDCUC5AqYkQHwDkUYZVUy6y4B62SQRLA8dyyjVksZ3VpVqMJb0
VRb0q3TvwqNG6hUY8vUxYDfobblIMCq8OIV1V+N5vWa+jHIE0BmNsvxsIlyYcuREkbzcViiPqxEY
xFRtpJzwNIUqAlFTdvznTq8XG5dz9LFmpe4zPo5Z2Jm6j0umlB67GfCQACbc6ArN/Q9al7SBbSnx
fdaoO4+DHaMkoaqJkfQwGGFRqyFceiwfc1huabP2FJXchYf2xnOA31Xv0RKykjHJDGPbzhCbUvDd
WtAy+v1goVdOCIit6Cw3lxOAjxNTj/KJ+sovQQ0ls2/A8zb6p8U1sYmIqmg9E0R2S+Q2eIw0Xm1Z
/CLtuTK8tEulXntb3Wni0uEb5EaQ9N6JT+c9M8uzELVGzp6Q1Hh/NoC5vJSCc7TDA+Ybfej6kFTy
YcTVZChd0tFSvGPtnqniPzjcEv3IMshvkSR4fLgcdU7H+SPWMZSc9frGJC56YRh/E79Bap1H3fSv
jLblWhKuFjG6F5QLTSYdDMlCrTxNpEvjStV2JJyZ8zhCl9mWJv/7hvKlMgwhOrOQaC8cnc4KYBqe
5TlcoYQ7aspTTS9316sMCwTTPG34VCNAoN4juyKp0NnIMA4c4N6hzwgrfyqQ/SClULmvktNehQ+u
8E4sz57c9bzs65W/vq/4H6ziSln+hIho1S4o2Wp+4B/Ce70ucNx5gF/Mb+4lwfiwP8OoOAUa7w07
/OR17wFyuqFQIHkg3N+t6sCMSXK+xGuLwKg1sTLRyRjzg00G0MpSMGw0UBCxsIS0ACtjWTZvcCsI
w1GbxLrQ8eJxftA4CUsAzuUW5uxrW0mT7WDKdXRHm9qP4kMDgS+m5/zvIBntFVrHFU58RJ0JMeil
dogc+jLsfmLP0f5gg9QrTb/3To53IA0y7CXqC64wYhyIKF7xS+D40722f5aXtBzrH+OPiu0HsiTp
THysqQN/NIhlQblJqskRAwLKX8Q3bbmLmHN5MJRjlY3Hsul8qyiylII84Eknzxw0FbUDB7T5xIvZ
ExOIaU0NBAlm+1spGND+7j3aBaXCdtSgZcYTgBjt4Y8zYS2mYvNxJXg5x4x3Dw3HG1C4bFK44Tdl
X4pe70gGI+MVy8DF3DTICEJO9PvJsQ4xOUrslFHOmAwf80OvYavPRPACI++qdnrG9u4r8cKvsQ59
+doxRYBFx4LX1OGozTrjwi63vfdjTRJB/dmXs9J9OF+kZ+9b/U9TAftcfVhHZ8QY6DhjXlgmCNqB
vv8JJnqwc5x1rOnX1bld74JiPA+ABrunx/+WRP9PvxIZ3jZVZxdmlPqGOShsbG79B4ZAY6sqAGzp
Qbdl4HOroPFfUqIPoF7Gm7pksGfD1+k8gjam+Dpt0QI/w7YzQKlva7ke73Jxq5M/Kt0vl7r+EenT
Tf7JpuO5FmncTckK5ZaMugjSAAIaUQFtj/nGnu1t4OuzODqUysj78Uzysm3bCTzjTobMgGRhsql9
Oa2fZ0deOIGEpeWOF7A5wbbJtZrf2CgP+kgmssDgPR8CXTjj5HQiFE2yU5BBZ8b8NjnvnA5Ng6gp
8LdumY1TUktHBti+kZS06gxSyDQ/3dBSjsBt4d6v7b/7QlCXZXuwG3ER+ssJJBIKiF975+1aoR76
1uSWdCmpmy9Sprp05Gmexb7oP1OnB8QGdRz1Eu7GkPQAJZYcgsGuk5EO7ksCwEsLkuO0lWv8mBLt
a8H6i9gZN+dxcAiCxUpWMFaNqmtz6bSpNqu8xkfB7ihqHSbKK4tWaYv21NW58EVvzQ+fhjRSuwJf
KFqEDmOxVR2g0CrHPaYGXfYb7/+90FCRIB2oI/k0IE8lyXlXuaYqofl9Ywq/6eaqNhA8u+9uF2AD
nERcIwcfI5BMIjObIGcglJP1Rb7RojraEZayqXv1kpJzrbH1m/L9qlYO4BpAUXou/owCOb8zDxNz
kCPAYEBUtmMTNStcfG6iZmjjmEgN1f/qy+EuQrcBGcTGg0hti2l93SQH6mTD2om3w3B+S9QAcjc6
lqs3TOToui1vtEqp7jFFTyg+EmBh23ptkp/PfPEAIbhY8KiWnyFsdqDN/cmS6XOlkBoOOsNv8dpq
D5DJhl+hYZtth3sjfpjBSAv4zA5xwJlDXrUqX/fyeTWWtC7gsYfZh1D3Z2oe9Mma31tL6t/Wnse9
tVN3Tnv41e3LKQCOV6OYqINlaRcAd+BCE5jnGrHKl8LYfjKImLAaGtLQefHxq/rPY20h89S09mir
beoacnyj6USn2nRyIGfo5dv3h6OqxvxfQjp66tpyRpvf0bKsLafcn0W2ydj9BViPFdBoQDLdYQns
YvZUMuc2mZ3XoaKETbIljAf3/+wVlA+lb9iELEl7lj5E6D95vWP3iw97yeOXDx5/lFew6MiUn+OX
1j2wkRQ6zPfCP4ACwFFwS7mCNuPwAobvrH7H7c5/bXZLvuq5PBUiKeD8pD+XjnmANsPoJr2fU1jK
OKtD0EmnMfJ6zbey+L4y4LWzEuOPRvCFf57mJvmUiiD0LQoZbUM6qrpULzNU+Cad2vmfmyegCut+
EK/0DDDWUqAH95P52Pj4ceJfUATe4V4fABzv495oKDPNWK05mAMnkgiq/N/1x36CEg90bIraWmTj
kNsBxO2PTqWimN83uTJCz8tZ85SiFBPqMplqFlp4iNCkmVMmu94JB3si8Wa+kD/nGAl7TFZs4tZ1
WZdjj1rQe09WjSRKvwv8IU82M9lF9C/2zOFYu1GmfYNn26RAA5oqRZTST7hpD/jubNFJQ5N2W1tK
Z8tG9bmGDWrgDmsds7oGBGK9vO97uJ1RywTWfqK6POM8x3DEOHRkH4oYEvn0gNJ+Hz+B8lCHXPY3
UuDxQEtiYa47LHWkhMrXYm7foyxYIvlp9QYvWhEoNW3mFBktH3rTxX01w83AFw+FjFEHrm/6sDYp
b04nSjp/jHKRgfwC2lINmJXhyAgz7hf2ErP50w5IpQ5akUbGM2SUlnPtoznG/beGiFxvsX6GHEHk
MCIzKc5XEUQ+OHxaA0bZJcRoab4ymuZ/RWvcdG7fwx14nXnUcs4blE1Ioq3ttXtoDrjIjK+hm61G
JKfHYbLM7ZengRootBn5lcRVnLb/S8XojDTiUsA2fj5HEZ7NIpdLCh15xPTuex7xDck39APshCMf
C65QI10IafJOTMOCV8UKScKYShRG8qiRWcn1KCHN7bMn8GsEuaYVigdLqKZyNW4nyhmxexxR0iy+
2QwGjb7k+CZ1IhUPHDVRYORAko+Emb2/NWirliTo0NOaiQSkVcXotMnjKIOSrsFUPBrcSApXyPPs
3LRqc7WrbDtIYW/v1JqltDR9Ryn7OCCY507wXAd4nCN7cJXjAD+qeZUnlSdLVZkrETl6KFpgtFDo
zP9nMWPTlja57rqjofDBVT/tf80a6Vb+KBlg8aZNqvHq6eCfjhGlFXYmhTKvWdJ94X8Y6AenJ+Cz
Tyu1u6L5E87LdBIgjzzuDPUI2SzO1gHVWs3MjVXhYNKZoAyL8OYpJ7bsZJeYphYMgzVFvVDzwknr
szysIooYORxn2m0oJNvUu3aDzwZPsybJkEqySCGwC/TvBd8+S23YZesCj+gDJ2pGpw5DpBDor0h9
ZZBFGDO7h1Ziu7ddTeg00A7wOiwSlSJExjVLtxz9QeZ/hQiOICnVm6MQ/6KUmBvMvzKHzkWHVZ8a
sAAJeJHNYMKq2JbL/5ZoTCiVemCF/bNnjprmyCy9zXDnYHLF2Rqe6wHgxhrQ24ZfosECXI1pZS2x
7JktoC8m8z42/xbAE/S3wH3DUcu/PlJhzOrFSugiqA+kiOdMeyFeckwQ4z/Dch6vSXZUSGN2Ebf2
78wnw2ypg+PAxVpqOXaQNXk+4lapwpmwx96bt1ZM78BOI6pXj93gAfn5TKKqXJk748ixre1L4+Ac
mJsqWItzQbKIBLkjgpKXCI363lZF9MdJlXUlFqd+I/43eAheaTQgvuDuo+znPVJS6uSlimxNEaJ3
DaFpQVo0aiXHppJKr/Nm2+cbgulmjjoJtAi/xJG3ANXXzvy+0CSk7K+u5TcfLaCxhiZnmMcYgqUM
8Db00p3D92JuhSwLjayq66iLxPo4H2r5I98GTDBUjjzXd1CX75LjVtUTHGt5BlmPnFNLcNEacuxz
yb226wtQqLI20VGTONKaufBPyO6R7ViwM44dE3ZSJLPxN9FG/8KoDluveovDAse+HLSwKGT12Kv7
QxvG24QQyTvV5SDURQlynH7l9vnqxjk/dd1RaUL2oEsapddXT2CiOagnf+czduPvS9n+qmA2R++M
hbrEvzing/258EDFsCEyUYER52y/iSrOIAvnkPqJZK6bu3Zte2eCLgAbYNPOEQgbbroHPZ3iiPE5
CBXlOlh/EjXlQx/aCW8zkJTwuCSJCsgQbBxf+K6RmpgTUxWzYF6BOsQh6EqBnGdUalkSigJNBunb
klYh5aEq0WlerfBnHYsIPWeBQlWBpON63HuxUFTbnIauMRCzAlGn4gMyKBeXpVBpGqulTw/AMGNV
vmGqX+f9lzsEuRu/2UMdoLjClAkcvr3PmJCCUBt9mnV0rpxFiR2Istrwb3kq8S9O+MpXivJ+ln9h
fgmU4HwN8jErpvwrEG+E2hAT9Oqo3DMx+A71HS/zOjapt70BY3e6+wu0XLH15PBGTk82640n7AqO
uP0+og/x51Z+1JTwsWs5AvEqTvMlcxPUKEBi0VfV6iH7kgNQsF9ppYcErcRVDhYK7FSQVRvTWAV6
/8tDlnm0g04xOs3utwNsDDK/ID/cP4KUezWShTqb4hma8PqIciJoj7RmxKn9zqdc8396BTLFBVEJ
lDj1YVZC4DXDmiiP7/jcwBNO2kS2KArdx5M/uv5HgbA7sb4Sn3Lh6Oet2dS3JzTdubNBJbq8JkKM
XM9DLXDVMSNkBukhXf4iqnmb8jJGvLEriRgkX8xAmPO9feT/tSQfM/10mE7ZzgYYtjVwG1TTGYGu
9CrAbwnW1ySaPTQ06bQ2OZVCLg2NkKrouixjAmNr7fu/ODUeC4Jm7n3CdR0ocoXnfAMbFznaiBwN
r7tHurVKqBzIzuxSgQniI1yUt1Ho+LSxvMSHm74wkqcfLXHcOGVmHYUr9fpXEyiwgeU3WgYoqsBu
A+qgPuLgahY58xma5dz1iXPWgyiC+sQlUDImR3bAauF0WUdDWDVxy9KB0fkvjRWjK8V+Okb7496l
5Bhqa7HPlkemg8HwvQ5fe2foJA3rw8sdAsEg4hZYrIAMD3L/JpeiqQtoWP0h3MR20vO5ecsH/Cxl
vClANJCAMQ01ZU24Q3191sTALXjkOxr5KzX1rtGmeDLGS5rjePcclVnRUCmzVH1D7XjJuG0OjSfx
9iTGeQLGNNA79MahgGFidxrlDa58rxGSLZsbWs/2C5Wr8Ck/K96+mr/bFnKs15Jp72FnNjH5haiT
VWatosWa/KtJjCnIUHQGw6/RgQv8evC9qPzm9CD4/M0EQ9jTvVP6ABeSd99Sz3wk6G9ZOaRUDhi8
xT37gKEASoSjXZGyM8+ijpJqleZsm3y4lCTId0QdKUNdfTXlpwAT8dxZFIGcgg7GSv9lCb2iQYtX
/22O6dng7oph82IccQhpj8jeduE5ZKcYDMxji7BP3JnPs/sD3AwnFxM2AkZSoKXOe9obdunSYdiS
vVoPM+F1GOCtFLpeakAjgJ+W4Ri415eh2LedBY1YvqBu83kwBacb+VPgiWQbotN4pe/YCRzAMyHZ
fDNmtB6FQtTQLU3yApbo+3R0Hpqa/MjYlg+aCgLVUp9II8rtehdstwmz4GZPOa29+TuabVx+4KGB
Gcu58ti0MCv/AJ8+AzbhrxnfWGE3FJqTnNhodnIab/sR2dgezEXuUjHEHzNT6MfkMoWRQ8fhY1Tz
6Hbhmqp+jKEzjhikNBCJNaB/I8UguSLA2J0Kw3ZJRY7kEAbkcC3biQuOis3c2GmUhIiX6GBACMtf
IDPFSnFQ2lFIE5Dr5Dq+qGuGPed14eHmdl/nYWxEEgvhvAAXANng5qMRmsHyXyN45+sirat/jXRJ
2/+pnBId/507ZgWiJ0EFv15Qp3YHA6xix8gS9jUV0uZEXbIUxbmYy+6NzobrDAS/HwNfBE3FvudW
cj+eTiHQo1FOKgI3reIxIxJvjjqhwlzRexAcD6X1ewIXnUJIzh13oHemggViwhCaX3Fh8zXCXkNt
2x8xozSyGGT18rXTKNy0zD3/j4Wyaoafak4R+PYnbdwzBli+BGlTXOuW3qJexk4cQvdYAL3yVwvn
pDxcotQq2MrBUeVtHsyaGSWBcFaENfG6VLLH2IKEwGOylwrl7eedcP/0EZaPcKTR1ppFr4pcyNFw
5g9DqH/4tG6SWCkBjKTIArLE78+zkBbhsIy7ZomfpYirSAY7BbPAwtCBkYgMOBHyyUttESiMF51P
9DoH5nFYeb3lAFAZlF2hmJueGD7IUCX/ko3IrYzg5RPtMjEFIpUFuQ/NmVJMbifGySOStvr+u0Pv
CtZe6cJzh+8jWQWXaMBXU5WJLvdP4e03rGVKYbdJFQXcyoDCsEnoYlfk7cH/NTuAR+o70c2MBr3O
5UgKnzSztQxBF1TrYFPSoYJZCpeQFN5mQduE+1IKjnOYgToDRYJ8Gln1PWT7cMREFDwxShN6OTM6
aTW8flbAn04DQ3Zg9SVYuRqQ9SW5b6ySgerFl26apSbD3CiTJfJjFCiN+KU62cce6V30uAgC4BgF
Rp9yir/zgK4Nq5k8nXFsQiqq0mVUPQ/MwCyWdLXcsml90DH8o1DOkKHfEjhZHrWR18W0OVOXapPw
rFNytx76EnobJcexDi1z5BLNLkHtBIgE6igGBGh5fUXaQGtILVOxC6z9PNa62hYFc7ubiT2No37c
eIjpgvhIoK6MCaJUz4SHt2mX6fBFeH23/YW4ZHpS4JtROAV8Z/Wnc7rt8jYvzhp15zFkBC+/+7Q5
Cd4IVpFtjMa19hl0YrKN5gRFLpnPMwJTlItDr2xLt7/m6cAQi68ltHpakY8akVDIPsVOR06qE7Jc
04AA9I4vavn8VnhqQYB4FC/wB4ljNTfybbIwUDmwFk2eyT9u2efLnrfX3OyR1lpumG2TstM0+RYa
YzCYFPlw8Frx+UU/WJhuEGwXe8JAVuwG55t6H82XzXSw74uIj4zs3e3sx1U4gikUxkfCt58i6Roi
HK15e/N3yNoTUVHzn7YZ40BobhJn6WXTP0PqDMxSJGRjRsRyeHWXyWT/lYMd0Mr7yV9RfNjSiXZD
+wZfSqAdTpKVATbqWmXUekQm6EP00gW/GU+Kj6goZv0SJpU9RfsJwd6qKzdjYA6/09Zw7SnEt6MB
HcfbnrEyVAQjxuIZ9dcpaUL6MrUGY2D87K7DIPnvVddCHmFHi1fBHZ2itqzwXEbKt1Jx+FOAzX8k
rNTUA+UjgCqRKKqhrepztozjWUuEZOn3Qs3PHs2nITbemmCMm3Iwh9gBVkC45CO0pZ3XisZdAoOA
Rv3XtnEAay1sMNzXfxCuMNCSGc2lIclHViQNLM260AnPtPHL+D4CAHa+RbNYXITin+0hs4q+WMMd
iCh230NRZeIpwru4e9Itr5ACZlCkFdjDTZq/kGsfLVOuME4rTA+aru0EZgfT0ceYh+IOTcl5JvyG
s+lAZA30wgXijk3HkYyM2nopQtnyMIUm+2qx+xsyCgzZ0D17YZWWUoQcN7sBvaQPu/oXO4CSxBZj
POXzdBiD7L97leyhfYKIRs/ffbEkV1dHvkZNLFWKeHLlv0IGD41cZH8jOaMTDjitpB9BmTudjiG4
Z8lwpbRWdto8gTf9e1ZHFOcWLQOqpN3J8XOpOHeTWPiFhz7QwuwoM4vkIV57LW/jzcGCpVqOHVRw
e8PZuhsxFYlCgPPNS26yOtMAYAOmi4LjhPfuhtDW2ePD0j0ijPM7SlsRr9fIX1dIboBwcq3cX9Qt
l9Lu4sRa7uQJLqiUHd3BX7ASCPWnuk/y9zRxyKxFjcExPZ3/pD2Kgtx4MGgGcEC9dS6C6Ll6Y1Vq
hIPK4Y54TB9vdobHdvXgj7CQ/YcLatW4Ckz1d+/EiGqS5Lv0ZISWq/RR48fXXhibaUCTQtIK7Ey/
S1HdVhh6F2B630IWsT3rZpBMU+rVxxnpS4ONL6ohxRS0br5vaaRy7qCowk3ds4Bhpzu02lPZexJh
RRNMb5BqsE1J07SZygwMM0b0ol+fcgMv8e8A33Hg9yHGIq9eWYKrSZ8L0X6ILMRAMLLzTLmsi55t
6KML5XfhGXjM8qGLsSC5/krZdo80mNERLx2II7av+R9DYRS8m3PdeBD9cxeHw4JaXZ0DQSLePeXH
HnuqJerzqg95cpCHZ8nx7gurLZNTSkugQVXVIyLS5CmwWhM/DNKtyL3mCzwLD6NNUZV9YHcbKC6G
QlxWQy6muUR5F56tY7ZC2qKOG2GZGmKx8uK+vz56cFNiGtRfsWXXLCVLXE3ESDFwkNNhGb9Pf35/
GDBSkGFOa/vNXKPBDEdTnSiEJOp3dxn2JNWDeyalkvXeg2tgKjVcHXkyj/G+Vwxg4MY7w/TxQulo
G26fYZDoReah9sKGrbYezwv8k4BunM7D2qaGvEguMSAAF1Lzs5+zH/puqtk48j2+GQTSZctaE83h
NJa6pr6VgqI/1tUwTk7asgAWoZfkQyMQYkwq+o/XlPSbf7qXBMMaRWEkudCXl/g1Q6SZJMZGHkec
44N25V34n66Yafo1UcN/ZZWiFtnNDf3aJVyWTE9Vljn3dafa5pwl5kGbpFHjzeimjRs8fhz2/Vg5
o1up7M5N9mUnDJ2UqWzcb2lNy3tUr09Y6Y+/E/KN9RVJuBkNg2wZiK4uwqq5TTsfAS69wjtAr56U
//CPWHRxPV6xlpiDMQNZOlzFJIFqg+AMjI+icndwsn5DHCnrgEilHtUt6kEBM7LadTq9oaWR9AKr
7PZdRRYZn/McE9tzGloiWN7+iJZiYspS2nkOCh/hOoyrKcj4hXf0sCKYwSg0ZukyiFE56/LvXSs+
HygPJg1aarQerpS3sPjHsTYxYo9RQKXdSJ4vS0Q7DuBE5XtkiiUzU9mRscdvzkKDQ7R+RfOoQO9a
VUkRcio4w/Bh+K3o6336GVcb7XqYTohiFXl3xqQYSAXxKBSJXnMf6a7vqR8SVjR2AxE21N0T+zml
vGJnWKVXqB5UrmZtDu+Oy1ZI5jjmIL7JyP0Pf4a5/rfHPxEou4ohDoXcW/JgyfphZ5ThpnXk6BlG
sazDzT7nj5a1+mQYIdCkzZFwd24Q0d+1QLTK/rqG/1h49jx8eNTo9hw3dB5RGDO3fBFN7cPdAd7o
gNWkNTVwMAxr32KFONCaAmHsQiBQvw2Z2DEcsZ+VudEFVrnGkATIv7MP/vYy6fYKuqspY/YzR1MJ
8/FiIgzmGzy/Cbxr6MAbI1kaahrhuOE+jgyBlOVVrm89VgLcf+MX48pDfEieDpiEfVVBufyDIM0Y
Zp+aHcGc6jiKnipy4c/JbdNBK92jUL2vyO4R/2lcLHk0MmGAy2vBnK8m55mT/KOX37jOjRwMLi49
sscWUlBDCMxIIN8jL+vKLOgFE7dIV06T6OLkbsSGU+YPzoqg2y0ViDcp9/RzCPwn459iL16SX54w
Yu4yZs90lEzsDhHt6iYi2voxAWG5j70m+WnaOmMC3mKCngoC8E25/nLdhk7hxgoTqz9OCLdKC1ax
bhoPk8jcly4GbuXaRTSSpcsZkwFScxAraABWU6pnvtg1gkj9mXpmumsGSrXJ+Lf3pnmeoUksusnY
FaPw4h5gYoyavYQoH9kXjKrYoXy1eoAY5nVjJa5EH2qYRXO/4tBg+I4wTo2ytCfJCQhu0iE6QWL1
uH9r46pbRg4nkK1CmOq3N2jIosXBR0/ynUIyQZPwzDpSh9qrmfBlStyF0kGtnFla2Me5xITeYIuS
J9HosDIjGAYS03yP4dmybHh1XTShKc7xmCt6Kux6l5D/yU8fK/2Q1i9hIgElu1u27YfeBOW+gsF9
/Xd2BAIDmfKpAD0Brduk3eLA8Gj5Alv+3flpjF+Zi31AAZwQFLAdbKzjS15JT4E8Sx7rbX2zEfiO
AL3Acm74caEyUKhGvyU6LMaKrcGIes2vUXwo68w1XQt7SQCx2022E7f4C5/X+yVebRA0ZiPLFirr
Vx7MmN4iL8GuMMsMENnKLQ+fox1Uq43+y4vOOC5+e9YlIJ84YlcgNdwe49vq5pzCk3xA8fAhVcYV
2hsPdKNh6wzuN5w+IpFOeXNvAyZqthhiJMdVTRRmvEFfb7L+dJqb7OonMxJ3XAXANCzJcMRfB04r
n2tI7c39bNLZRrp6M5ZVvSTmWZ2KX2TBhdieCvBTpAh9G+bNfei3TrEeWIVHa8StjG90fs2X0X+d
sGFUnDxh0+DoeSinHSrdoBi28nsIvyS7aIJIAhDusVtCYsA/iXbM0nlQUXGTvtaqc3nC4qcBAV6H
gDCbuR8T93lDcH7tU7/WZ8u5387NWpNW4jmyhlN6FYj1Vi9IqWsVrskVFet682wCcUmXKrtiE3Cq
8XWeHgFjMuc5mh6CBwR2xjLVvbIiiuAe3eXdMPCqQPbFlGqNHKPMKQsYXjEhEkIAHEJql9BIi7T8
3qcHw7VmZ8kszvK+3JqRfqZwMaKiknENbi3nr9vGewqy1OE7TasMSkdtCmCfhBpDfdjNG2UgayK0
5p4MltvjhC0FhCUrpfdf43sEPmztvaE564ML4nCVvaFGI89Dkl3faqhCgt4VNNfXUA1KCVQsg2o2
TWdFJz7VptONQU1gzz4n783HpfHdil0A6FT0CeSraZDxKoGQ2U2tMMy8BhGNzJ7dNf0Y6zkzKroo
TEicfry4tTdNJ37UySnK+AzItkaj5I8KCsPbpmuRtwXFkBWSUp0yNvSKtg6XiM1HJRJ6+ByLk3TB
OuXIzDbN3CjAKm8Xl6nY3asd6tLNezb2m1LIB1/xe2e08skmLLBqtyt6Xw7j+BYujqacwW5Ihjov
n2cze40tGhMrdv/0Np/xOexBtAMmSEcdCIjzSHPItGYuCzMKso2szlgJBxwTY4fVwSxS9sGysCv+
Ub5NvSrgnK4CH7rITxL62QvS+VQJgdghenxmEkHsviTNGIkJKVZUkjU7wuCBXuFF6JGg0vTeYS7g
ZPThEAdWWJrCkpXSK2TJkcs9m9XbUgPQvmBs+E8wcPaycbZ2p0asy+SFA8MqRMGCy4ya5HN/16Op
TpTzY3e266KfY1psMCU2k/Jfyiueu4pp9/yUytkjJ4QyWavPVeGgzviJK4nZXeUkuMSVlEkZkV5P
suwEY0dRC5Xctw4BvbjGYc+SBxxarC3DOf3JliV3N0LHjGFwMpOf2CGll+fsVjE8No9G4rMfzFBi
jdnICIck3afO/7zoK+kvPgc36scf4EILEh+aFyrpdTdZ//v1oHQ1/AphPTBkTy6tErsus+JOpKD7
I+Ai3GHYn70tt8BrFGVfEebB/BkvDJQrPRd8ZMkbW99ZyaZGZXl1YfFLaqiWfUxgVACS4iJJRNcS
O3vmdFHYvK3uwqW3KWn4XRkjkW8E2tbUEJdR0k9k7dD+OU1RtfRqGy262BSXbPajaGHy6RsJw1H6
zGny8dDvddskcVo4qSn1NrJJ7GlX/m3LOeCTHHbSQ6DfHjkx4mPdZZPx4te4Hh9J4sAS9s/NXzOX
XOiPqcMfSvHP0y69Sh6cve/5zbxWDl02+BSFbWzdHNvFNXYMsuHS1KV1SFuCUFpNiwhgeTcN2E8M
iZ2VGtisCrZWYpUdcm7SmE0+HmrwFnL+wd+cO6v4ZVijfFsAsdQN5kchEOow0cMi2hQPI9CvITTK
vbfdLXKuzpWv4fiH7gqUvlpRiD+gEW6sNsiuLGYgOCK3uBkLuwvqh1o5cbiPSyn/G472kmWWGB6E
xscPn6yJisL8jnOUdX/PITbQx7Suz6FQAvO4SKd7/Z32LLNsPWI9G+9SO3ZDTbjPaOJYcop4wigl
EwjhfLqfOnHKWE7UgCoghH0fDDr958ID5Hy2EUYysbm6sr7sPl3smsACWWHZjp+5OEsU6HJiHgRv
+p+jRYcGmc+9121+ZXIH+euSUlV/UFjvwuUiwCuUyxN3CWVn8o5kX1P7t83a+Iq3z5z3HvSQ9XGl
Sw3F8JUazC6K4fHh3tAQjRmaVrTk7XhoBxTsbrtu1ExWdTixPhk+bVia4GxhJDUb3EY8yJW1Wp8E
0WE/kgb/0SghuH5I4OYVMlHF7yQG8zA7vq6bIyMhCdhHba/gi+XGK3WC7rQy6Qf+OvtWyLde0TjI
tzheyKa6+cp6BQHj+0D2qCBO9S4rCRjmiFntFqu/EDx17xKjKykF/lm+s3iNbgQ07lNh2PshHzjH
erFSw7cC3COvE7JXxcoyLQvWHlJxBdB6P9DlIbiKt3O5awzTm3hU1dOA6dSeFh7yF2sUWsTum4mP
zxd9OFLCn90ZkUlf2C/hdOpZtB3zlApxqoqc/nsyuIE3BbeB/EhqpkDP9x3Lh2qjQyYw2hamGFtd
nX5LJZnLj7H3QBtKMNl0YUA8r7ure/8dLMXj0NgKMojojTkhxGTtTue/wWlQlIFprO0cmmrcOV05
05PhleDi1hMWHLS4La/rjg2UC7B/uSftcR0Zp/evdJ92myczwEtYK4oenEILIFlzNEyUPdAMyWaM
q5U81YK/HHBSyq+v0X9OsE6sW12jIQiqk7c+AY8GPv879z8PlQM0LVIV73n72yYhSvZVrzSiwpGo
LD/wtg0lsemJhlil1s55gAKmy4QZv4w2WUMf/x/FrnjlqxqyRQsvR+XjsDen5vgqftK8l62FJiX9
7sUjlRtBZKLH4yqbAwKT3dO8fHkcSREQDvNLVj9CEsft71xkN9FIb7Ht2sIQ8Agt+1QxzRqbYlU0
KA0EYbT/nhe7NC5B/EpdZsYhiFR9QXIQdYL/iM927FEELa0r7EERiuijJje1krfEBqnnW6VcdIqm
Xx0Voe4PoO0qnjcXWpx5IHBFk3Ore3pL1HDabJ3KssdBkvY35e9zGquFAQAX+4T/4kXNCBreR/Pl
d1RCEX0vYwKobMPtyNZbi41HFtQApl7asRMWnPooTq98I9emrw6jx6Kjgismqv4Ioy7yMzvd1mnW
7bxp4ip78lHnl9qBwpSR671EhoOwJ2bXh+mP8/IJZJLZzRVVhgZMwREX1Mq5SSDqXB5cNKErh5pn
392NQICtiPZML4w1+DyYPk5ImSittAlyCorHO+K1nwBEXmfm9DW82TE3sFVSao2eovrIN9EsBkt3
oslErmfwzI6F17gCh0Zmk+9z5QjEwTikv2/GbREFxdbhjTYi+BpDPYLt70EhWY1yZFYEvFCBjK+A
7Vgyb7SbauENC5/EOoHqkevQlbTV7oNZeMTqaHLsKoT2b8fKuNtJb454F7hzCvYsQBvE23wwPhdp
6Kqs2F9/TkqhZ36fceH7rHulLySto6rNUA0Dde00ApBylSLOGLFWh7wqSJ+6OtYXBKu24sKWxZcb
9IO+oDVkj+wR+zKvSEy6VNs/YsWizaYxiUaCNquX0iKpfrYLw7AVmlxMo5B1n5AtK4ZuSFNLKCcG
x8TuN4z13hXgMCoCiaVMijXr9cx6jU9SN/9yVpTphPw4gGvTdKx6YBnqx373KvXzF3q3ixs7a/dt
0pYn6khWg0Mw+gAlTPVORekILHi9fq5IJh9PODSG8f0nh6aP1KwNHaZMaOEBlEG1+m3eZJ1LT6gX
tAg7mdB1IXPfdfrA62xp6dpgRnaa4pD48cc8z9deD/emyUfuY5fetw7mw6U/6HmHWycjDutBg5QV
Jdxz3Iq5Rmk/DYq1Nmq9U57TICmoeKjPLuogBWBnWpbZuVZRZnA7vY9Hyi38vUkCxn+4NQN6zIE7
UrylNWgWAqPZPy9Gg39rerWPE64FMUcw3NbRT6fR2HinVSvCj65xZJYTzFHz8h6GnYvlk4NSsmb4
Ya+o7lqIhQ52+ZDRewwpUiHhXGZJebkeptT/krNReSdTE7+VJhNdczMmdeh/PdIUxQTVajodHmIp
C0XyYST5VpaxY9EU6W+dwTgrBTvVh3QMgggF3gjI2zFU8x0jam6FnCTDo2LLzLndMrC+3LuBeWpc
Qum0B1CiucQuCcaCnmOe28e6aGOeAzq/v/6Y0udoz0mZqQToT88/y/07zBmSRYYyCxWQSjAn4wci
LLeLSfySkuk1J/cBNGPQJ44RW0WLq6MahzFQAdsuJAmJ26QJhEQ2pbwsPqfL7shkS6mN7bWB9RVK
qiToTS/mhpdavLLe2JJLw8uwhiNtkyeJztBFny+QHIyVUVsZ676gdLpvRPDOBkFjpWKVHmVrSxcH
8luNbZpkKGnzs2KFwj5nFQAdSPi7Pv6TEEBT3FYgS59tC9KmI/8Qdp6nwEHLej5IvrsCHUxR7kzd
IGzD1BF+sdolJwFWsnJd7vrlREC3Weg2C1xnrze8UPKMUw/OTu9xOKkGRsBNETHD4WjCNpwZOAPI
disSUlaWp89ReiCy9ruCfCgVRLD4GcuVbu8bVssbUx1XN5TBqGVnd6FONwvvhh0/jrGbos413UZU
oizxj7KM3CG0Bn7PAE16ZR51VQo8q8lwCdxoe6K/O5xMo1BqPYD/9S2HPTlVfKFhpPOL85m3rJL4
f9wnfgSqCrLM0FXN6RVPiyOVFXj2qtqrdloD98uNK9MRXFi6Gf5s9d0xowkVBjQByMpPcMnnZ2AD
4WAo0ibDepodjsSWFL3tsnP25yUSxUJ6TlTYW51g7yJozSZS8Tqe1CRblTdORcrFb3cH8OxfpV2L
KjyiUwUl2Zh22/D4yoIHJG7V4p9jWkpcSY2tBi+slZa1e39HBO4l8h4fs1h2X9R++hnRGrmrYYBu
O2diID1WSdsmDm+4QYFIDU+BJE/vYkaA6BMYf1WnzkJEShF/Tzqrfwa3KS5xMOw61A5i2aarQgA9
wdsu2DWVZAeGVDbVg4RB0+Da3AdpH/awwbN+f0ta2sXql/u2fkcBUdtB67mIEn1dqxUJkDkmdwlf
ZJlybDkqkX4/ruHTQTT3G6Kn368/IAqLDkylhXdSa9XTMfLjhcrnzwIrkd3CH5DECTmV/3hAD9gW
ISCyxxisqFcgEDrvNOKqklclTvv1D5+6TZ3nZXDqrLCYWhbxT7SQaEM29hrHTUvB+zNMtgXqyNS0
ovsrvdsYmSwQ5bHEjh26QZZcBo4ux0M2ybny+7KY5j19gz8BNz06rQs26oKKlqQVmu9n/qeURIZ7
Ot26MhAwLDZx2iO74NTO9s5YS2EPeAJMi7csxwq22aMzEZ4cgOWpMkfTWUyJkp0yyFCwf+Y9WQgQ
rdTbsaxfyk5K4G26/bsOBODY3SQZNdrJ4jcYGb8bWaIHfhyhgfUTDogzFOPI1Kq1rfFeKHW/Zb5n
GUjmoAXp5EXrDnl/SOsR0U5ljMN1OP0NAs0HuzZMKeOsEMqSqUGdQD8RkFlqy1qn7c0lbj2Mw0UN
naOUIOS78JPsFa1fpG5cQzZ8xXQne2nORV2Qi9oG0ZdWDSFu5TzFSEX0nvwZ7GWg64WIGvpDT1v8
iwLTXnslBDxXbB63VAjNM5EKeTrtWjIhauT+k+znT+eIina7HCs1bqiKYRHqw3864JeSq+DREa33
/ORBhnLptIkJAWXiy6ntmf9E4uCUwdeT5R3KNxhEYAqSk4lHP3vMdCtnCneAA+NBgBmFv8C08N8c
fyMKurhDcqPKuWusv399coJwPvJ5QX178T4jQ1JiGHcqM7Eoo05RxoLe0QI6VZlYJ7IYvz/rdE1p
lrm8G16DQYgHr12QymZlIJsdtNOUN2Qm8ruFoo7AifItdpHPM4Glg4mOWhKdH4LMxt5NdJ8RLDT1
eUsmdkTxGyQJnUXmVzflAzCd87na4Afm9xmrL0ZoPluNU0dMbakDN+dVyVWWY7dhTtDn5uwYeonL
Ki1fTzMsK6nL6CRlC/Amuvi9+YAXitfUqasmgFdywdyVmnK22wvbBKPxIpAbWm/WqRQE71qaTFWW
mOocr0BZEkU9+g2Qwv4eiYgKBHhgwKVCZutOiZA+3iUm9100qh1AkAN31BscnMe7CIXOOHXuKJB3
Ucr0BSivsB7Rhyx1uUdLox5WxmDAfPoThR70bUcn5Oq75+ku3d4msKw9g7JYZm83KKic1iHMuH7B
yIPA9ABK7nqycVGkGCK2SADsnjm745h76F1Xv4EoDAndwWgkt8HN3CA0GwRS3UM9U01lmFOdynsi
RP0Xm0FIi8bktsQYdU0PLOMyg+53VIhIvIqdeuqBZuTf3yA+QcOijzaMvuq9zAUc+zgJZiBZA5rQ
buw9zVI42UDiShKXg+vFFNFZBhD66MqeN1DI7AP5rpuiIgdVzwb0zr+cV+fU346hUZcNzwLyB7S0
KgpGeFV6PJBLmgquEigeiWAagEfvD8LzWfCG01VYigUiJqoLmEzA8QWHGsD3eOHuBsmubH44/A23
yyolW9s3bXDBYDddg6ls/XrYDjgS5XqSdinzk1xXG1BD8kJJ2FmewdeI1N+GZ6j82hFOJz9A1obz
hZSYbMxUNQH/cdYnDoEio/+8AoF8FD41/51BtLjwdLE95OpKJw+MadDC73sXYEjVorrM0IZs8MTo
lfcfHs7n33Bl8TSle1GyUa9C9KS4OPZ3o/EeEBb001ytxLJbdTGMYZLTEi4w4GWZtoPaBYMo9Xn0
+Oyunz7RKtMb1P2SW1ByAAcpUK8yJpN9iBAofBogY53/V0ty8rfNJIbx/iIYkiSmXU2g5gSZHMaU
BJafjPBRKM+yuy1xQorBSe3phitQGVQa/zzVkAN/wnnqVXa4kUOSyKt/rMnosBaNeysBfxws8hV9
8uDoZTD49vOvvG4EaWzuGmLL7y7MU2Clj2YWAUCJMxtTg8M68XiCkNQkyjmYrykL7N/L8u2FckB2
iRzFjl9QXkJaoRg3eH1+23EQeeSDMVhiuDkdfBLH3/LgiGAhWTIAJyV3E7DPM3TpbZ2NrY5JpSzk
7ylM26p/uIqusIz5hrsaTmL804ZEEs7kNlEqofE6WCDJDD6YgffTKBAyn2vmdWRRDrUCa+sS5CpJ
EGBVmaD0oRNMgODK88rJfW9+F0kS0AOw9sCPqa2fqrYo59ilP04xoOjeTK6UXTDXTx8G9u4BfFXz
W3R8OlCSbAgaKrLdIF2Me9HUFruXwJSXLKGcnX7CeMYvXeC/7l3iM+0luZAoc3Lmius7LznLmhfY
MIX6p0IV3wUBMfus40gddXQy0wwzpQZBi23kfoI0Bsam8zyw3fUTspYVdOMOMb0LT3NuSDl7xcry
mI+BgqKuQGsrENG20UV1hVmUkglejoBYF1qCg1deOQOeSCB59HVgkWWiyBlxCjeFkEmSTI5MAIic
2i4/TZY6FbHNgvpi2vyU3vhUeON74d4KMgzrbiqejjFL6IJD48rK6+kswchLMDI8abK3CeUWURF0
1a92bTTGrNc8tHKfzIvrbeSV5GcHKRnyWpUdJqpSfSGy8wsh9HoS+m4zTO/iMJFFLVM0rh67a9f9
XCTuRZjNxK3G4Qggd6az4CKb2E/EHxFptrgVqWJkzmK/PH2X+zBFFpVV6/M7esMrNWxN3c/RtJQo
8rdfUZB3HUHazECz7+sR0QmmjV015KAlMIvDxLAx29IJbcGSnNA+LmPyIpS7qwaypHv8m/ktkdPz
beMTnxMo2mdPgsgbputew8et9Tg4fgJ4ujDbnEHfLOTJeoRIcpOT9ddSkggF+X0oSZHXz3jrpZK8
KAE0SqKWq06aR4FKKs6UO8NwGPmAVkqUr6wzylbNLAxasUke71YdxUS3RXbs5oapG1lxG3+ZYnwb
3fEz2PwMXK63FFxAUlua/TAuW9LgUs0GMwEUg7TrnhDdmP+P69D7Y9UGbrAtIvuxIALZ1NcNVc59
P97Cc5sEa048/EyuS3x0uF8ClkivzAXleeH1kk5w6cH55Oc72D9srxnoD9SCR2z6Ye3wS/Thrze9
JwsGe43Do1/CsISU6QDm7gmsiY65oSbfc7eXKuJUZINo4w6lgpNodRV1IgfNUNYcO6ze3lFedf+1
gWj8lHpYytA6OtW/8G+NWmrO7XmYcblD++Ldx0W+91huM1qf3Q5PxDqXuNMke0K6I0gPwj6nC96A
TBC/QUN0XtkpoChjccSj+MXfLN9q9WwASEAlMY0n4opYYrVAkSuuR349sGV7JJlxXWHXeKIGPk//
3ZQM5Ek6nk6gslTtz0S0aTnSVsEB+ONGlSnU+wmWGZ3QPEPGEeL/heNX7mHSYACaYT9G4Qspxu4B
ukDvW8dMBV7eO14HUZtUFekoQfYfNE7OtM0+oqXhGDtP+sAFjxOyTPtlg47RNHSFafDKLNRYybLt
QC/rcInHjjh04ll66pKslAuSmp0405Iw0KUeuTJjV/IQaYJUEwuHssBLrmXY+DEev/rFdryG2b42
K+Ka47fQOInF0JfSLWOrMFPuPk3oiU4PnrItCo3LCEeivCzozwklpkjRIDI5lkvrq3LlHvTJqH0Z
ctO516NMwFFgKqFs2v7nb1/WCC9HR9mdKQoTYksc/xtjq3H6WDTgEhVCBjKKgePdc2U3Fr3GT897
vV2F4xfgP0Lr2ovkVKfdVHmLzFsSocpTNv5q35dQKk33bMBDxAt3+DiwvJTUtGyiy0fSEcM/reJl
KLvpttjnaamcpE0j6k60OXVuZ2y5twg464Zup6XUqNVdvVom59bQ1CwIpGCEnjM6w0LOrMZ8JJFk
SdKwmbMSF3Rl8Usfy4e8D5hRRZpM32aItTLGWJ+1mzHkCflqayu1yRIG97JidW5cYebwJRPAut2L
bJPIu/HH6vqFPV44MLoPNREz6rys/3o7a9CjuCDbjCarZB1lmowCF0DdCebGPZzdAfDPcbIayAw4
j11XILIYSzuGSh/+y086S3JAduiiOUM0R40DZVasTF+zuWkaiypM494CSZr0jn5LYPQ+fGxNLK+c
kPHdBv2GF/EOeEJGM05OFtMib1mYBlSE0QOUDfKuJ5hMUFuWtVl1ez6nPqYAm8e923PiqE2MrHmE
6mufkSjx/wmVYRHmsKBh3tiHrBY6eGaJI5yOwcirCdF21mN3ctGhm+gxsseuWLJn1gBQOX35rpXi
2OI827xUPsUxMaFHf4BSpcgawUqcWi7nTkMGi4z84GG0jESQQH204JP1Sfc3yjqzES9QyIz91OMO
Sb+Dh9zL4uhOK/CRwWDxnzprUSn+htdBd4VPNW4iAHWNL8CWM4cqVNqUaPdislUArDXj6Wj+veu2
FtF9hPmIRPe3BiePejLk7X2UzOqv47blLEMVcPrPfeQv+WguDBTG+SQQcIiv695aJ8ERymB7bdD7
eBRne8rHQT1CRomY52DzTUTTeWdNrihNKE1vn4m3H5DF89DNEWqyr6L81GTNMUYDvxgq8UW+uDwf
2KL6OAYhRyvV76h6JzqORjDz+fO7z7XpkHzyJl9OWhtfdTZb9jltbanaQ7fg+Vyeb1jeYRh6acIW
Y753ENroCPhdh8QwH0zobGDMLCUrgtrEifPutnAeYJg67gtKny7B7kaHIfZU3Rx/sRYq2EWuRTZd
5L7BQz2YaZH5X9CBYx2WhIOvsX2FCnvgzVXY+Jm2ThEE77kAVafwouaavRcMywT0MulZq38oqbNe
Q3sN1RszdFPSxUR1huhYbXSSR5QWXT0hgTV/mmKngk+wo7WiEmuOWF6nrVv7wY5ZhoJlU1K4EpVP
LMkSmSbBkmM5Vnu1pTzfW76bfK2XcYVRCLJgPjqKIGRtjHXaF8yTrTKfdQV9ZsGunb5++oBLH3NV
MD3+Ws/qCG0WEDgKdTRurZTdqTqwJD2h+BQ1DL5Fbo3xYRYzBcRjzE0LPrNEhPwWEbzIbZ1Uj83z
JgkvxehgxwNQyUAKrKoK/TU7JA3AMrnN4617W8AeBkd7+EReCIhsRVX7m/MP3eZSLt4IZ7pTrKcV
HITHaojrlDzTOIX077+91HjVeBpe/c0ErZadQOeMD3Lte2dhB4izSosON4Di1CpslDEtN7cP6+TG
pWWA3gpX82aYk+7kzG894fvLYTo+08sHJzcnG6P5WjDvivAWamRkMF3GV7LzfDBkXTPsgfieVZ69
CGDk3byOt73xvA4yrzFr7P9WA+9OYagSYA4K18wivSktsI636K75tlJElXVdbC56u8YR64AxyLVk
KYeqV2U74MghEngbR6jKgQ9FG1ewgjRgBHETEui273rI5NhQYD1xjplDFiBcsQwbKqXjIFqiVHb5
pcKIYpoJBHv6Et1HPJ1JXtlMaKEZ0CLm1N3WbHtNvOR4Bii9RBp05u6DByjjk7dI2ygn3VaL6m4Z
9cVk3ZOyJIXLisS1V9EL0IcIC/YuszHSVJluVMcXZS/ZeKoMS/gnHlX4iYF+JC/6jcJ+1YfMG2HM
I6vpqt18F9e/oCwIGWXVVKP6CUK3NO4j6dlla0l/FamORgHdR+tJhw574Iebkgcrx/Se6i1oIHJf
012PRzHGVXf8s+xEkFUqlUW5Kf8pN7V/TQpsAtrMPMXBjKjyTGNf8FIbtZ+8ettvfIzxNYas5Mv9
wW10tz8wjzuLe/9jXdd2Q2QGil0bJWkML9SlVI6POOPzWz0kY3rCclA/HZjNVEhDZpmOLeukGVX0
KuX2pk9h6NBvZuA5pzCkLJ5FopGMTNz1oXTuMr2SjiCqx2WK98mtO3xj1BRtqIZrazA64xHBpOKt
SUoG/wBrPnCWnpFpieANVaaEHIPGtgsoymvYMX+L1natL/srbXGvGCTHS28kD1mBEiFJgrKsYNhT
kMutnfnjSbOBt11hkVNMlgmLYq1gCPKfGVLfJHYE3NX2PpefBgnM32jZ0ubHOHZCVRNzCMZgYEBc
nkY+k+zAKJnHdl2tRZpZkEQgaCFLhZP+dE1zAZNEEtbJ6Jzkzv50KOoWkswejmhWJ3jx6+Xl2OWL
EvcMRDgR7TeaDrIJl7tY6gVF7q5YKiBf9DiqpKmIhM1unydPG5jjU9t4p3rH1uQB6nn2AiRySIik
QqsmcIeMcKpBREH8L/L+SkuYKSH9xWMGpkSfKdlhV9MKVj0MuXBP8327LI3bN81qf3x8AcuJb/Wo
Si0dIH+6unlsI+CAAmZblSOR8AbNVFnVH8GFPAhm+w7sgCOQUgCslODWI0UDI3HykrONan5Fp9Os
qaDkHwttqoi0OthZkSu/+D4x9SVSN5ByYNoi5OwfcecZe4+RQjpQ0pORzR71Obx0YSPuO0etzsc1
suEM6r9ph+YRYUqcA1KWOHU4ezGKLgDFDM1o8wgjehhU4TKGrRbtp0Zz1fd2QI21bWwxV1n4a9Ze
iM98TV8VbGkdi8he+UgZluQbYXuupgyUgy8CmNaF7SYLWbcVkaQr0PnSClt/7nESgaCkU2/nSTLO
5N1/lr2Ceqh1C4ReKru2ahj6jyKv0/FsRNFpF0lP/FBvkkvYxf4+9Cx3inmiI53OUsF10ctQClgE
GECtms/b+Z5QIBaApPG40GAZPJuKjNHa8J/MPKnkMCXYzD0mH0G0sspZ+JCRG5rzrre8vlshWMpP
k25Sm1nc13t60dQejSl1JsNt5gHWjD3lOtBLf+55bKTqWA3sr2sVu1AukipPxHBFYiE/zDcSpSad
6tvk+ts2kSnDP1kLfr8kvO1WgqQYJ2vabi//0WrZWnMUYdlhywAe3i2WVMNFqa0gOiEC/Mg+EX2b
tW4U0ntAzh6xmv0Lfl8k9TJ6xiIEbdjM4Mm3qI7BJZ3qT/2we1OD1njjrfknwOI2P5rQhynYoL3G
YcMK56kQ/eY6k0LikeyapRKsUPvvrhJxJbEUuiaL6FK34y6j+1rPvnP1TcIuDkYWD3+AW7rtVonu
gBkb+aefVqmSVgKA9e65/yn07C9hZFYzWo/DKUt9Gy9b33UL7hcNsdnSD2a7Z/3fBZTNDf/j4H6w
NDvb/4G4gHI30Y/sJifSVuJz3nuJ/M4HkujqB0getcKpLJSt9lOCyJ304Ln61uwjDGpt0egNU9Tq
vzpFRyAdf8ReqV6BIr7tgjUq/t9Vp4QlUHBon+cUWUTgJ/ceBHWgMbwrJ4uUMpo7nXGR3dhbSt1T
cxiRnp4G+iqmMROPhnSA0UXotqLxmGDL5eYQaT5wrachqwbiT3DpR0keyAehPY5CJd9O1b8yseJb
mCfpxR/aJBmjWFJV2nbTbLUeBY0zGFTJREOvZHV0OcycgLo+JpyW52WFonkWBGDBVxcGRYpcPTKB
rSfIwW0I/T+HYNlB4P3FfHmEg5qjfm8jGCx8q+thWC9f9fU6yIm0gR450na7AyKIDnPZOUv4yMgC
rcWLCuhSn3hs1bo+QhDlJjR5hQFdUimklRi8APUnJcqSXGNe5GhzcjkwsQf1CizCWcMqFM5m71PQ
rEhfizJpbtn5Uh2zgDx/a7i2+GXksm5WfeVwaLXRosVsSfkmPutKyIEbg5JWv2apE49MeBhcfQIp
5nVhAshJX/ddluvB+4T3d41KP/x+ZD3hZJCCt8MRwF3eTNaR3T0kjQlpkRnBztwk1EdFwlgGlIjb
uL63aKvTSn6PudIyY2n+SSyRQxZufEv7hAXrLaUHy3513xgS91k6qQVK2TxJS4/ZdaQOi9AuZkRu
m8U0f32jdawzWZEUwGo2mS4qb71lY33NzAWL4Dekk0htL3L5misppPH8Bi9u9eFfZr1oTNazOm3H
7Y0AAjzHo448hYKmZCjOVszii0Mduk+ThZOWTX9dtf11/n7vJLcO6K+gAflRxqHw+GXY2C3kzfhZ
JQkB3D42i7x+krevuzzu4OXJlgB57lro9qPtKWYPfsfjlFcvHzGcsWm1bLSa5ntTXf/GekBHOUOP
5/N7I7KwZkV+wVAMeSMP80MFQZVWLAu9s/MUvjDCXaHoLA5h2Swa5+KDEO5BaQFVkzqPBGblJIVb
elvYbrvcXE0P4kEBMKBxPoJD/YZ/gFSa89xI3cUhikerKL3iY7X6Nno4ZmayncKR7AmZjnALWmLU
EiLZV72oRLW4DA82x0Hxr5KikXXcEaiSUDMbySM2N9+BNXf22J76+h0+qnJ7Xs3PXOX7bAiiLCHB
WLtnqMDeh+VcpibCN1QwruQlmSanvO8IBUD4NKWzA+rKevtSS7hvAlfNNWa5kM4AxJclsQePASG9
RjhVU2t6Rb3i+1yq0I9op2SYZySzVwD9HFSYP0U3UqWS9wLs9F1m+ojy54Ol2/Y14tkp6ItX8pGn
dVKSqq9C3a1cgwFxQd85IXLchNSBeDsvAq/04KKqh/gvd64PC/qbrEG16Nr/JMQDFtdu6SsQoyPU
+cyJn+4Ih5TpWWzjiXV/otjv0Hx+dTUrOwIofqXCML+Ss0agyNViKsRlVUexAb4XKYxPfc4kKYXr
2MwfNKCLsZGk0i65ZLUa7lsGA4zceqW5b1OUC0P0Q9ubvfBdhMFh1uAiu5XfBlh5V2NowLkBBJMJ
pihntRFfrEz/h0ifq3mDN8Zc/HA3MVs9AYFvydYv8XqU92L5cl+5rJQN6jB5fuSOkSYw4y+clnCI
KRW1ygiLb3RQG9tKk2NqGe97/EAASn41U2/TE8q9IHfOmtbFV7ZdvY4VVhQZYBbNEKYfqqPFeCH7
SW4wFl2n+g6lSDOUp9G3//dTwvKn0uMoKVpYwE9sLSb2WVzrwam3Q8Lty8Bi7WSh0jaeFpKBq0vJ
ztqdfiePn74q5wfwCOTx9vpTxIlY1mp0k0aQZwt3nhfJXnwyBDC2YZGAlMajDtB/m5ooKvo3/dX3
MpqjF4Gnfl5DNnH25L5zzMpL7GNnV0vsBGmemkl3QyoRP0qWiB8/Z1VbBe1gTho+omyrVqzP0UA4
BImwarF7n6vT4ARQL5eNzIBN2rji3py+NtyveFxymbuPdLHsdQ0suoM/LqmOq1jcM4zwJEjYwKv1
ALTa4qqDTkAvPiTJeS+YrqaGB2EYQ725MGLNi4NvjiahnmyrzlW3cKL9rLRu9zzpKB3e3cHzac91
+fPCqyTTAXgLM8FdaGEvHgVrRoaY7bqFx8GFVsr05aQ184uWE7hNt+HUoEXqg5cyki3IaPw8KHkh
Bcmids1dIvc5kcJI1znwnBR3g8XPIu7oQquZyW+3stEg2rUYOo1hfkxbtn1+9/Lvi2GCJVpVTndo
ReLlYiaYd3M9/1ore1TktAWmpf8rvszAU1hXHkXn3PjmlUc/NjyotUQA0OlcR3Ntaq4p8JN/Qc/r
318Xwwc4QaqybHN62fCoxqmYrPYAscLRgtq5p8uBw8uO6LMRQTS4FCK7TvXhWebbBXgzc0ceMza2
b9BHVDHl8AE8PNb7BB0cHycZekqJcsLbXuclqbVvhJy+RgpOPAvocAtSbwM3kDUz1mwoMEW+58De
n9PEtzKsZeA+an5ryh6X093inDKLLKrzQBB9QcKaJuaSwNx4AGjPSTLIwBqzmbDVYUHUSor43Yd/
B7Gayk0iMu1rF1pBBZxJQVvtrY8JhUFZCk/01mdpjRfSLYVVxqzlSNH5KkaOWAyih7CeDQBm8T4/
g/96/ApVH3KCk+xDhe6yv51q419fQ9nTBntgl6DYgyYv6wakc8W0s0hfcAeb8piVO1//sEzZIoBV
nLRoWC9DWyFkiBk1Nsxh+ZqEzFmGjuvve9aVzjEko410cl/h+dv0bakiKGsMMQPeijGLEd6KrI5v
LlzlMqZKRKNfJTjjm891KtlLFSUscdPOB3AOnT8F/W1tqD7Pa4ns+URBaOKc66qK4NqrI6t6Zedd
8qwPrMT3qE6gIE0ITkiK1ih/acTUFjOEtJnf9/kI1CKIAilxCWIgVhMV8kTq77MImf/BdVd8gK3A
/h349MgcbkivAdA0zV9s0vNLZnlV737/EkvHE4QaRKgphKVzXk/hdKCJ5ntR7AcW/YdSNbRhIo4h
3saClICcplGS85VNq58UNV57DKpaHd8wEOHcNcBci5bKGpGi2y8wpe6P5DG+FdkfK6WHV1HOP4Kq
ZztHn/1TJizE531xstlCd8BSTRvbbCb9oPOikbOf8oIbybliL2ZEDSD9oZI1SAAmqMhXOMNyCRp0
17CwnshmIo1W0M/bKtZGahIL3UPiUkKCcTnDu8QJUdCodtFWF7CRH5RIMAZlN8e7Njm1XxmtmgDa
te7QfwS6bhbGTFijhf+mR47mn3J6Z1jqeX882xnFo/cNUDDN9v5uYNS17eViO/p7hPYnyvEVTPPy
iTyJXE/tO+fbAsQQosfzgrqzCfI0KROxFI5/qemsAQ7IgBDX80J1mDj16qzi9NyC3QbdcXJ3vbVj
pYLbqql+pJDJ838UWj6dbQzCHndBzH0wC5X9zszkyf/Cv6RKCnCRPdvTTMewF7qRwt6+S9beyxJU
xT3iTK3+YjaseW7bxFsN+Ec58mYBW3iUaF7vJs3Y89pS+/AGNUyZCn6xDOcnQqSqVZDNv9BZcBv8
Gp99JVqqDtTrSYvfbqwe6c2TRajZsRCqdv8zqjD8NMC9mgUt4FxZJ963vsRXOTufgm5ImxSKkOVX
AeV4MV/CXXVSemW4ATs9mb6KQ9GLiYmpoX+3FA5XbTPrQzDslNYrBcrAA92/OIXyMBD2mR57fIdz
DZNdatxd02WJLiL4fc8ZzItrg4N8OSyTtO+noOQfNvyDcYG/lI23oj2LkMWF7JMdkOv0bWQSKrtO
HjDRPaIVFnA3V8zqsndigBb1/D9Ex9E4WfWpWhG4vUVOD1C9qQGhtt37ufAWU+l3tHwz/tH67u6B
2tO+f9bo8BIm2U6iWqSfFAUATq2nZownC1evspJoIgeNsxw55OMqvi/ncVTOkha5sUnijlVjzvjR
rrKI/sbaqNMeYHRYlvNDHANq2bZrMgv4GDkEb7fJxE+AgAPqpwZidjWrDeH17NrQ7g1Lfr6mqzzC
nWzvdgMtArSDQ3UDab7zpa5IE58vQgY/wVeN7OK3b36Eqs+mgP//Ce0PmDj9FkGP5wQ3Eh6Fk4Dz
1qzk39w3ROzHfSMr9n0QNrEgZRpzMu+45IxLYyGgEs3grDmHq+2sLq9ELzM92uHcNklAmhvfOIiO
O0gn8+5Gq8BNY9g5A5gCr80roxrZLuEyLfg2xqUY+DNc+tCGZ4DPaGXlJU4LZkoR0T+oVHxwxDq3
SsVnvCDw51IGLtOHGKzjZzTc3ZmC0oV1xefiYVTLV4cf4OU0iKGx1MlxC9IoNVyT8NG5E8+eXD7U
Dfxq7LlEc243gbauVcsOhE6jlsQjKxbQLq7PCSUk0DGf7/QYHkLaN5uuOlXGqo7A9cLbHtcjZr8K
SSrSPpO5te6b8jqq3IvH7WMdWKHtO2A8bRCRm0VBAoh+BR3z9tuq+PbKk+54ApgItgKGonIQxjRq
saLxXEI2fKGqQ2GbU9XUuPf/EhojEfUHFDgfR0CAnIiFcSrt5GpBnBJ8KOiTO7RbDJ88XG6vm7p+
tzzQ+yWNdjOweWe6JUJ4K46Vs8wlTJsdv/N2wgjQ8PYD1nha+/dNEEnqATZ6xDvaWGAYnKMLkUal
MfR/ORW9Ud4D0/u8o4fjHkE42yBPkVG1GbnXL6jgVyAlRQRn2OxuxIFx7SittzX1GGfzjHkYtFzy
sXe+j0N2P0RkQx3sWjMcOhfL/4ipt3acejKwr1iV2OgEtj+VcSahE3qMgp/Y4fyYunNbExDPYLL/
0nhzUNIxQ7vdYc21lncHN/xgbTkdL4b2LPCGw4U0BF5tQx72zhelAAaIsHe6l5k280cjb1sdte3d
FY4YgwViBYkVgZkoA/vuToN+dCf3C6ok3AHGNKzY9Xk4+H+WqjlHX33YGUbANU9xmxkubtIIcOYL
z3A8O12P6GDJvWXN0HX8u+CTkwz4lR/Lj+KP7t9KABjUpy/qVXET183f3JzUkpIP81BOTJIai1iO
sLwxkMYyY5TVF23byCIGe5gNcZvgMx3qGRf1zXHpzV52YbUUYExzr5FarZM8Taqr4xg34h/xpzrK
Ig9TMBJw7u2u6sI1qgHocvTNPkNhXBcTVeSWKUckgfT1lOrNw2EZb2dgAXty/FJ6StLsoqKDSC4j
DSv/lDJ8qiDDPkw5cf1XA0+eFAwR8zy2k01eFUYfLCmDangp9z+OpsPvVVxVhcftDMYSszYOfq0Z
bT2sc6Hrs1RY0k43OUfOiOZ/76ut5+Ne+TLxSC5eMPBa8umtqZgv6Vua8XwehoFyrr+IRT8bOsw0
EU23IDuOYm52N9swnqozStQMRKDpv2Qx0CuTMgISqt5ldOfU+9Syk6KTzu1vzh8S9uE8oniYuL5c
ckrFwlXnbjX9faFZukA9zexFX+cRLyjzhTBUZFbeoP1rVqabkhqCxRrh1WBdqUQQyCNk1p8URuhn
R+MFf9jRwZod208Nfy6mPF6YMtD1BpN2h/9ReI+SJGvhfsc08osydT2XMxxBh96OhaQf7vN6Q9ZR
wcXQiOeR+eHcQ67PbTED0nmd9aC34L8L0erW64wduGSfWqLk2ZVLaYPTBzLAoD2+KA285+m5cOmp
OktRWmSqPKZ8EIYCvr9mjRMDdkz4zchferZD19ChnJDyD+qlyj7XIRLlJqIdrP+mGrz395jn5edw
lhI/IZOgQzXEJqa40pA+/daMRfhkYUTSVe5Kjk4ckD/9E7W83Z4vEKe2sayN/CCkoe+dSu9BWkVh
PuYzLjnistIbnnbYpu1ee3KEIDcDUaPUZEAZnoLo7kc4ZvEJI3ViWxuugKCDorTPDkbB1b9TOMJv
B8vcOn9LHJXW1uoOjXryqysLsYzExPiS10XCqmFyCdyysRX5Hvi7XQ4ldYqCsa/3HbmdBcbZ6cz4
ZbsJTw93FW0Ny4nhSCCuutwxzT++6uC/+iirIh7dB08vyK9LOygpLpg181b9F8QRfI77PJ/bJg9L
e7q+DeoE3kxMfizt7j2pGQe4Y+sZGY2Zt4LlXpOz4VHmJoSvQj5mCmosLvgh6rdrOXNqlfbQOvdQ
nOv67VOw8kP4hIxVLKjFX10jPAEYwsFhX0FSspjE4X1VcJN90LuQDdmDv9hjNMv7P00hKUtYYp9B
ZWI3fpefsZmFN9clzhKWM+LGJWV18DnUAlklyTVZWd37wgwfwgHQG/CvoYDUL3d6QSLZzzr3YIet
jGbpYyYOpv5gH0QKKCVB52pm0/7JtDVW4uo7fRQN1tIKTbdoh+f5MQRvXGcTMfgZpCr2XBWvPe6A
Kvfc965sR1XcyjDRN9Orww8CGYqhkKVjDx8EgdHkW6CDWCVvqOJ0R2qbLAF0pk/kKsv/U8v/RCjl
wHZiuThPcvTSa6B5ug9xEodcwS78MlXcY8VUAMhSqIBGLGlWGxSfiAMQJTq1mWF4fYGZpEpZTeWL
2EGSCE9G6LBFpgMCk5x4y5YlYYgEZ2pgIjvsdNcD2G1ZtIBxnKsbdmGwwYjUbVymc5dS2MVvd8/z
i6ZJ6paaxvcgzyaE3lw8i7clFbiN2ViTWKa/ULzBEXKKu/fbCcJXnthgo42/l7dv+AoO1k+sxu/I
db4DEpWsH9xXU54KJLE7zE/BWSk4W7XgqLP3hmGrnb21FAdYeAxyf356XZN1hx6qMl/wi9Bi/spt
i7ryogFMZ4J6CGe4y8Si0WwmxsJBA04sElzOEDx3hWIV6BzHPyfC2ow/hg/QSV5xXxWJPQFrejWc
xKQsZ4kdQP5uZdVWzGMPS2mxY4ifv70bnAQS4sAZfzUOjhfG/7hu8bEIJJSkijFuNUsMuys7pPtf
eyRbfJT6ygCtmGni4ABjYO72IKJKKjRJKEnH6JMWKBsPFVIsRNVB8KMCkkaV6c/h5/Rtab16RtQj
ax4E+diXB5t2xx7ofQLnOzkuJjy94I3u9hCCnaUfTZ1bvRe3Bd5Od5p/4DYOpl68IQyjy+6OM2k8
Nho/5me/m/7B6xOldcD+LWc4YIbtuuKsqZN87QhFIdTR3prdUJE9t1KwxhmU+imdGwczMaIUqnos
nTV/EtDIHMZWdEW2fizeGlvqZyMUBBtNZiZi+wYgOQlwxddV933RnvEZ7KPLtmIqCuMhIsVQG5E0
l8DtB4XBtSNCrSnBc7i5zW/Ey0f9Cdc6KjEMDZ7VryUFCRGBTebOfhzxVEzsPyQQ3adT3926wz/V
KA1ZpKhGO+wR8RcakJh/c3nyBn5whGq2wRYrCVbetLHTbImEX8sfDZc/LuHKVtns4a3ShdYymbEF
dqoe3Mo1NbzHqSrB7NsvDdesWnDSOeiBPPTPCKEpnKnckNH6Mx0nktsEc5RVzzTcrZZRs+AZ9d7U
Qi2cP9fhPRZNK1heU8dgAcEA9RO+bIw56D8E8KTiqqwH7Mp0nNLPizu6F+ZEIKL111cMUfyyoRT/
xJb9VVoQ+tRpeUTOTqjm1XrwDo+OyF4lhJwSoWlF+ila/4LvnNOmV4XqKRvMJ9ZA9r0qsTyTxtIx
qLjsv1fyIn2od3FVYRHL1W8J6HJBv2z7LJgBJXzgFDqSSLW5tcD5tl53w/2ZekZSkuZrp5QrJdo3
BKuh//gpUKfhmzQDif5xTCHDxRMLs7Envqot8tOoDK5WNsN85aPyJQGmHDlud7IvUyxH4MjRDhSv
tC4bu73X5yU9xewMeImhsgJ4xeMao0GM1FT2UcNqi1sRcagAPICPZ/9kH+KJLgDaynWpbHzYA5Dl
zL29KrqOx5sszLQtudmB1Ec3wKMfRq0aNhsfCo3RHpbPnNijlfiyhTY/+aLTEYQujmFsAdPx4DGp
h44WckfgnoFRKSVAwmR3ZilLG19r1Mnzp86oSj/GhP7Bh2Su7xPxEGYwMUz9KpVa/DRpQYzvY5FF
wOsSjdfGovNnjVLaHarwzPmHTv7Y51exHLcCFIgfRcaL5NYTLijmT9e1xbr9QuLJL2Xzyo2O0Ztl
DHLKnK5Sfw8qYHDJ1kQF8TgEb1SDbiK/5A8hGcQNivd6YJxdEszlqRTSg8RsSR/QCkQswkDfluVf
MM6vntXL9iDLzCU/C8YgZn9MjHoT1bVabUSZI1WuPYyCmqb/Wu0Yf/3grQIIMSuIUy5NiCfxIAhb
Nafn2iFWkxRkehCzC2ojwu1nPRAQmDUtxJrl7C0U1deezBIZKJPOyK1SI5femDrN8V6YyTOby9Gd
hTeGq+Eevj82Al3tZJb5AvZ+SJNhEpHHgLjRIM+S6DpZl9zoZ/EXVo/1u+LnUlIcOOP+cSC+c65H
+lF2x7XOJaVE6elK/PPbkfC0ZWO0JNt+5H0yxS/m9TOIuAcAasU2bG5qKPlktPCuGMSkxy7NcWjR
AzpKBceiok7sdAmylP7CRPLDXtOjAqJfhmH1auy8+UVvPWVl/QGl4IB/K6DqUCrOrrvZeo9MGciQ
Tyh/ob1ZobEs68YAg/KbYCJ/an+q6Oo/Uerep3uwJdkVjbjIWwpHsAVG4l71fERKGeyuT4s2zZs3
grERtObwOCfLB+hW0j2UKLJkLiPRTQKRiLmdipieFLc1b4FRqfvCCY9jIlUv2RfZXEdMYr13YDb3
ek30BjDK/dgNvlXavsRQzrvD18btcIDZF24+zdmZxFtatam47e2fwE6nG+NFSRgihRWqCFVDO3ql
SLR1oG7oiOJ29UA0V+cx7HDe8K44rn03E3ZyzfNwqvHg2fSNuRWwYuyg4rG4YMOVM0Ws9yWRwjqZ
ps86upBExAKp/FJscDgkFIPyLONU5ea4XbhdGP4sY2n8y9D/SpRHGOP3lzZKPp6dDS7aCaa+msHD
YjnjAoUoey356RgQfbn7YeSlocJ5ckbKlGWzD5lVEWQ/A/ndNAX26vIOWsCLrLAIGYgpSopuk/UD
1ai+QgUlueQVbNerCny6VlS0SCLpw2sqlO7LfHBR5clWilM90NN0NSu1gHqIIyY7Abfmg+K3YhKF
SgZXf5s9/zEoD9Sf8aCRtgjER2JVmDRLP0ziPrUXshEnS6NiDGA/eUhEOBOXJ4DeRD8slmTdoJe0
8/YFJAJfl3+MoT1ufZU50SqxyLQtwcGTqHd8lkcY+VmAt3xGtvNog737rK21tw1IvP7F4uPVvYXd
r1Jxze3YM7Ym0Vad2idn+ycSxeRR2ZSnXtjREti8X3a8YdiQ8EblWCFwp+UpBMhOIbfOVvw95I0P
Bbp7mGqQxDAF9yq2ttgyq+SkaVQKibvVu9qMlhPS9Hdfyt8GcmKzdWBau6HaiaHTxpGYc8yKG9ll
bke7l8XUt1Zk0ELoAgDnF9bBC2GRC4Z4fYOUxmtnHtVf4GMa6F/EG3Z2MFSPsvhwt0/zlDuAhRjq
HtgTFcPwcWi9zGMIYnUmf8aAng78jBt7wUjJXxQYMzZiJ4IW7GjFyUms/xM9lFwZd2BUl9oMZeWS
4pFsAuVr/JsbygkegoonFC+2zwH79jFjOHVtJ0SoV15vV2+uVUgk5m/lwaHa9Z+2DBAdWdxht5gu
C1019ke6RySRDRz6t/M3dLQX4Z6UYbBLWibBb+eIVm+5tMpi/KXxfEYsqxlC2jWW2eA6jrh5DF5b
muYYhsqliCJ/AJVJLVoXvW2wEsPSvgNy35Qo9XdD5CzB7YeqcOE8/GJT7ueVd25fXsrf9GAo+1st
feaKFJDgOjRUeLHy0ETIzX6v1fvb+bTthCm9jlTT9fCECxd1i6YLUu1W+5m9uIR22MHMiW9Ksm3c
drEfhlZAv2wW5OgK1rwycRvTMCJizpoXYRzRAZBB6QC9KHk+usArvONIkUm6Grz5F2fvLdSCkIha
qE8hz6ZRP6Ma3iRYvynHYwZoEUwebueyqvCZcANh4ToUHKXuSD0R9Yb50EpWmC/HhFVimt8oevBh
HTM9/fbTUdFdGB+/8rZtZSbB3VuLAw8MimJziz5t5Tly4OKPhvcutreWzZWLv/e7HybX3pajasuj
vZYhFOsyeeC4TV9b9tpHK9y1t9deAkHtwmfrUeQ/29dMLuz7c2NBCxkPqHesG3iwnf0X8uLtV06D
wOI1SYV5VQZddgjQke0ezZmLZreCosKpmAh3Z5hny6b1fIawZG5FGi/A9cNNdMmC0svlM0pt2kX3
VD2VOThupV9rxKOPuMcb8PqAtkFOTt7iN18/DKl89EhQLW18S04lPA+OXmR15Dn5l/O6EMeteBNo
I3+JL7k5rJNxSL9csJhy6nZUDKtKWTzy9exXe+pXsUxiQ6R9zuj9B2jj7og/g+53CQigONjnqmsM
SspscCRvh+FxVIu6DjKh5NcUSOMJol9QGitCRJdJXJRgF0asTq/CG1MgZwwYpGwyYfK4ZqmK6+gZ
L0TO195lp90JB24eX3JXYsCLBDWD7yOjK0tTMe/SbZEFQ02OCS3zCwa3/g6SLis/4HNO6lJFOYFO
cfZpVqbA24JrBt4hAakWfDjIIka+d/oeGP0CrmvOjIBeUXm/jXWPXZU6FsBbA3ygYOzogfuU2raC
RzbAPLV0B3iZx2Yt9MuNEG1Wmyd+LsXvsYl3B0p+1xAvEkbtqkkhx3FrUImrhNa6MpSlML2LbXN2
iTj/ng/9SayACDy/XAQlolRtsuzZS8g2RHMxOaonwtRolB697O8newqLEfBBVrqMUmVhqUyDR4/o
GBtxKI6T9Re1YPAMv3+FjG8EGIyBUhY4W481JWbBHjb6RTXysuLGKLCMw+XgRmrXD8/6BZWMpiT4
vrAK0azIcDS7H2ey0/NrF4qL80LJ4sPCBeRKrx4VU9bimWuZMugB/Hsgd7x5hbJ0rA1FL3jmezwu
lFgKb9aQpaz9sAT1G2se9mKoNJxT9VwBtGH4W7Je7KPSxWoN1HIQHYCXQMS80qWZa66a4reFd4ZT
8J9095qzs6zYauO6uLDtcusXf6g/Ftj1UgJG04p2LpwYIjtUYXqjJ5n2N0j8rjnsspgCKYJqnugd
ft9NZUShzZXzvG2ka4HUq0zpQBZwAZ3xdGbuxjOVB5PP1bJPNtmI+Db/fWEUuMD6dDUgBe7kRKqA
PP6TvxKHedUnVSZvpsj8Qaa4EjxpdrLCUFg+XhVcDDhIUv94pWdbmqB0p9jlyuZvd/nDRjQU+SQD
WpPbwXjXPp/uLkZ7w9+pPiKOn5VcnqjktyoQUEy2uIa+rqO0dyzZsJAdJ0TUI3enzLK3GGlFjKnz
7RUZLJq8Qe1XODmjTSbrUbzCMK97aZkHuYZq6cR/B+DbQM0aqaOBAk5sGSYc9aGtq30CMpXgdUfL
rROs35uxEIE7iFo50UTPhfOjmkhcXVZP+NSD6thpMTPQZT+PVINqxeSEc5E8yHLHPrqWY9lhdAJ3
GtxMgdF7eqEs5YjsNxgJI2/II3Rn5pJjIZ5ZgH8KuTEBr7uNYvRF6Z8GuCguofCz6NrFh/nZpCF7
ULNeV5AzA15R0QCMRwp9teRKmwIDZktMxDy5ix6Ue03z8aU9nTfY/ZSO2MpAKvqeTX36ia+rjc9u
slI9lz0UHC1OBhoHjwdN5AlR2zrrKDGO+bYLpL5Wm+NQS3Yhs860HupXsKOTLqbl6azb0vOpTjeO
1A85GXJB2GQ9au7/SpvabiSi0Pss9Edpl5nt7qIfS7gr/Xm6NcHq19opjphqWlBWA1BnHppHMdGe
LfT9ylNQMmXM+7lMK4LYI33gIWM6JI55/KtJataQ1tDDxrHk/c057lSN9OMNkMkX5RkmuSftztX0
jWrFrcYiSzkrixggZ1WnvI8n8N9VPoDlqbriInGdsWS5T39N2iYbAqP1r2z8flF/ohM+Tkr6U5AW
HcrutQd/WqgIUAO9faWdrg3m0PRmSYe9TGSA4AtOzQrzAMVav3qYJGybbVpYsSMOqvwNOm1dbU48
FL70G5OG1lJhW3f6DjoB/hb7cnBxFbk6IY5bqzes441Y560MOFZSUCuFMPXZ2/yvmGOauZgXzkEJ
XiWERDoQnJA9TxSc+mSvfI4diqQ1b5Go0p6cjYe3T8QMcDpyHDaBJimJgvyuOoXX/19RYAhHYhTs
LFQSkYQZsw+CGyWY6aDrhO/6hJApblNFrxvjnFMvE2IZ8VqIwkj8dUr3QjlKV/qwYTqn4cHdswLy
b1fqTiFcYWXqHCc1Wj4OIf/QBD1amCqwb7sqAfiWXkAl4AyHS4AubWwKOLBpOEKftRxGENZJ8P25
w5nk11j3smiVmwVZCeiYjTBHxVDdyoQnliu7yadwqpm6TJpNzHA8pbfFJ6trE8d3qIAp1XgpJV0b
ojYeYuwm7gYLj++1MgJcas06ylRK/RPXZh6D/dvjOORBLbMMIMvoZi6brHpqmjeRIioLsV1cO/Hk
TmYtgNaeofy58aWBx3ELt5kQu6f1YZuI+4Sh3d/mghsRlT7kRL+CaYtPILZkr2aC2VcwmQjilvJs
zwTUq2ABAQhQhaYyY6iyPo2OhaS+NsykClDsyaRvHWQaN8/bR9pLaH5h0J1WSWQ4PCzJRYX9aoi3
DZT6gLPxXVHgdG2iMh9lbgC4bS+PRbBM3lwoudPnxlkOqQ7svzaG372eZEC4+T0FOFMm2Ty3VN2t
9j+enIjLalLrpqWODaaQMumh0lmwup2e+UJVriAWfxi7yzxBGAoFCLYjGRo0zm2WLpJ9G/SFb3A9
BZ72+y95YB50MsuXush82eMXRf5gqnOge6I9P1TE71j/iYOJZ+/1PyHrhEZ6fdkFPzwKYBhEv93M
HVlZRN0+v8/ek0SaohMhu+zucf7Wcq6AP4wI1B3OGILCCCljpcZC1VWroo3kdR9p/5e5jjvAEHyy
NRPYzweBeeoA75Ajgrn/gakD0J/SN4uK4zIy/nNQOImT3TNrv6KNOWv/J4rV/N5SPBUxfAGImDfo
H64qbfabli323w/RFg61qfvRXqZYp9C/yzRBa0pUfPwHidpaT2G3hiQE//Jcdiz9COgIEID486cz
YIpl8BackRYTK06ZCOceHUrDywsXT8kTxZj6bI4MYNpmp+KGqWRvzmUMcFdXUJ31x0G4RQy6I5l3
zzfKj7gP92YTj1Y7XjbQpab4DNzwV6+qWDvYGuPs5ji8fAS5rJA9TDijh+CWxb5OTqui9clyZS0N
bh+tSE3UkJt8tmro5x75Zbpg+PFZS69cdfdnHXkLI2S3VRYeKGKd58Yk5P49u925o22xloLCup/O
ccGUjm6YXsw6Xf6QRx+yhQKhMKTDVDe4tE7UaA6Um9v7uoGxOsG2s4qLGDFhK66/b4lnWJ9WAexA
3TnVpc9SkeYSESzyDhtl1N0IgYEv0Ewvrs5gpLCV897gOoQNSWNgjyVsoKWxIHT8t6E5EhlGpvjT
Ig3skVsXg993NUUITxZeIMsf2WGb4TVHpnTuNPYRHWfE3Zw4I1B9XrGU4wHjm5JlZafOacYrksZt
SrVdQIXW8ORLKsuQOic+0gO+806K9IS65gZ5OzhNRMo3drZfxy0BJz0YZ+tMt2ozRpXCGa5ewZ49
3ju07WLDZi0A/ld3HNsxlf5RKQSt0Bm0FF9QK3MrUWOq2JJDzg2fEgN4cmd+bh5k9t7IQ5m27l0w
cZBJ2YHEW9A8hru9kxlWyYLPq9ojTVS7sJGCzhfd0LqoWEHkkxyyX955NmIWi4L4/ftass2fUoKQ
FvycJT+wtBYncpQ8Ww1qAVJZKTZ/UcmCCuTa3+A7ihROOCnAkNra8SG/anTt2ZkS+BZrUUIkqyoV
0dGV6qCVcks3AED5X/hrh0x8LplRn2K5mG6owy6NgI7PF7suCylygs6+/eudThhg5XkPfCuSfw9v
eQCTA83vJN6mqVtC8PDLo8sTpODhIgSVPf8Inrp5mJlcZV6tuHBY6xbkOGDITv8oVB3YoTKRUrdS
rht/pteeraMVtvVCpFBdYHXddiyg/WObrxwEACAROsuAcSyiB0Hs1Lfjc5577bmOT3dOkmbXXc8P
w3mqiloEl2RXR2le5TxovhNaGs8s3hUax5e2cFFncH//3hQ9cVfDUEGl98nwXQ34QlBTDyP+R71j
YaDuE68jpS0lWn1FUJ9I8l2XI0ChflapVynDmOLOW+19K1Xwgj+gG4MbfcmWhzC3LbjR9kYMtgFR
056t+/5xXnW8LAPsvnCc3ilnV1cpp4V9Y6o0eiwjSmS00VOJX6cIWAN2mNQPodo6uklvLsyrNv6y
3hZfLI/0G4n204RlLD6aEp8IOkDzE7s7kvvZF5nfgb6QRlW06yVcPse/+DXca+o/y3zg5DwMKWjX
DTzbZQqsWGOcLnX/CybCsAFAKl+nURFWz8DnrexjlNkxn8e477eqk2PfeuZdkOMxlvdHubkfmMHW
sfnWJAsRPd+RVgva6HLqrEofedKdCB2vdMlDgftkAc53jPMtaUaoHeX9d/iI/Dr7jlcFrE8+RYRN
X0dBUbLMGWaQ7m4qPKcjpWAfUcmBjWd93XEWO9W7AXZipASFS16ySyX84giFD7QL/5lYGS0VAuIB
67dVl2jU0raOFbZqBc8cZcXXstPsDRh1cjvyuGp7Gae4eyW6v47NPr/b6n//51vYDIFCeqFwD/oz
b2ufS6BjLbICzan7EPwL+dciJUWQ0ap52AoshlDVvEygIU6YoCk1dMRUzkHnDrQaDzqt3VrA7Ig4
4GyyAZyxzlVe1WdPfUMgeiluXbYXf0MD+RZSWzJv2ZsbE43vH+WJvLWCwiz/Z/av4LhBkXia6GC9
6CvL4NdPDzXwjP8DbHJazf/mpo/60DzVRF5n+rOzgHvv2Zn/v3c17BtnjgXG676CpCWwKSSeO3g0
VUSpU49Jk8gNdOKQzbJLl4yqb887aE3q0cx1f9KnaHHILGGcz7u95lDL5rQHxB7iA/RtxTOyndlV
Bs77C8i3F1V5ZlOBbXJRD+sikgu1BJmSWHPzfEM5i0XzfRMZuqgj6NgX1eQCQrx9kIJGwJYS3pjX
06vlq48a/VfZsSKEWLyWa9zdKOKf81JLpcquZ42kfTqh/wGmYb5itV8RIDSKlrl0PPxeGy67x7Qe
W2QVaENWyiNGsrJX6nsljw4hqUnvUD+wTNsOGOngtGWwrqstzBnAncfWZYMpI1W6qf8Oev2yYce6
+ixhY0EqIPIX7uM78Qeq0opzqWgGxPGioS11HEpEQhTFVoxrdpAtILEYkPJfilvBiAnGmvftvRdf
cZi/U3Fb6b3QaJlQSVIU6Biz1XR4ql0RlKO6UBj/cyEgELv7dq+zZG7fYlSMP0ihyij0MUICaDlG
OGYRsAkMRHDlFh4WzQqEKL040rdUKqyapl/I+Kp5R2E1yL02C8Vgf+Xgj1Ft4uxwIfxhQzoJzlPw
adhnuklOaw+45E56y7CpLiYmbgnSmBIonXIAXe/F68NPb5uIL8KloCxf80vFWWubuDUKzXg7bY/w
p0BGjlnbqj10L2/Crj+DYiUaD9cO9umxHPnkBjXnnFbDvOCr3LXq6QWT++t255qiWusJ1KiczFj5
lnOpDvUNiz0kBdb2Y0hMWxfuJKffBohs++VtOY+isIGlBpegcheAMKa7VcDPpUrNqB2P7eTo5zKP
qMOXGpQHouOkpXrwJv4XYvn63ASh/0E2nEU96isRgY6clwg6I3at8MKcGlqgVWQkJlIVM0ceIEOK
bkWTpoZ3zaCYd3aAPJoAgV1RhPL2Sc30luQK5JQQHiLXxCM+noqLoEAREcQbgcz7G4fX7YGKyP0Y
xBFEqIF8dKDMBFxev7HazJO4dzFqATPVOYUHO7n0LElLaGJu5Hq9ixHr/StjJDyYtHm2zWxs4eb9
hPoapcDBhXO04/2uS9k/C3zrCE/cHgrmeuLtiMSd2OVr/1pJ80doydLzYFxE9LwHzmJ2Fk+pMnu6
K+lUnwbg4pz2j5dPj4ZdH/YIqJY4mHlKrW0qwAbwztobHC3HKeaVshbts7nNvQb/BeQN/mOzW5x/
feA8rI7SZslJmokhco5Jvy++YLRPIdEg8NGuhVh5kqfkix/hBq9poFAR8cxgxCV0qdhp8T3ftSUx
x1z7XdHMVfBfsfKYwsk/t/omQPievavrDA6J/wXO679xkvauplL2jnul5LUmgzYXt6epETwwJlbL
MkyAD0fqm47rQOEsilG4uYwjEptThgz1nt95B6BqRg4eJU0abDteKZHT27FjkqUCbUtXDFRKQEu/
W4TrL1s0xdFbE8oBgF0l6ZzcJd2lob+rRfVs/yKNJZcpWaGTdQYdPMkaXpGDav+T3GyRtagPqDeG
VePSm06mbqytWznwWKMw8z1Ref6WWy3NXS6tdvFfdLNaPzzZdXsOKiEMZm+AdyT3tJsLI1N6T7Da
BO5ebZVjrfNjGio1fdiNup5TGcB8oR0MJtXpW2YP2VbL9pj1Q3Qi6NLDzVe3ID08Cv1OtkyPe0MY
KhX9o6f5aQ2bInGgcRzDe7lTTpQLffycZxyNYu6v6Bce1VCXYRyDQPU3ZeBc47hROVkbnRKPmt10
J4r0abs5pSMxMPZNk8h9b5T1RqCVDv9GRBTS4E+9l2YLPZfqVMW6bkQwL+WOJh3n98TL+bgHNkP1
l4X2cqUAe4KPj3gczM+qXaSTGIDFDm/s4rzoi6MidvXLWhVpAxfJj9i0dAPYAzasxR79DMkA0frt
ilAX5WxXDs97X/toDZUpCC2SSJDXRVy4QTij5W+I1oRCrdrVpbXYH3jw9f/dGkgdxlUvnVARpF2T
PE6Ab+JUGslHoxwP0Dpyo5SXQfyrrdTZ0C3TaosJkfXAYSrti3AmeENkgb+Y3qpaClv13//Me/qi
XPB+S4c2lDAnauy5+xmBhwtItTEntmq9WSy6vN8IAv8Bx2+TADhvYHSKUIVEOI4aZHJmOLrPPvsf
pNgH3q03lMnkGtyIJB4i/8X0n8XzcDBTbBYqRTNdjSodvOR6BCGYHcu85q2nD12AX6iTlFmVpwQg
UWprFDHt6igGb4V2Eh+Fs2y9HaxU7enJ6prrgQT830DC6g9jwKrgKGgBfPpN6hvaqOIBKadysDRE
V3kvhL6Bn8MDa7FsGGhNOkCZ7Ew83QUeTJVUGfa+22sd2EPIos3s6WuLvD2QUYuuZ+xmqOKifkUD
7L44cRUof79xtRmiA7l6yhOWSjnsKN6JBCbnv+W+CcHG+pOYnsji37174ayLDBoTKwyHRmhAjNCm
hwfE3LCVr+0cE1fdVcQRH2R0IJl5xweeJis0aULazS3RyRgy3eCu1yk4qYl9T5gQF4AmnNJogCGg
h2MEK8Pb2P/TURP6dR0BRtlzaWzD+CpG8fVuUj9ReKWAxqyZXEG2mWK6yA/z7vjY6IFGWb5S2W6S
oI92oBD1BgBD2d9rcldMvxyIrJiiXNVUWEm9KftTI+61H4ixGssKFcuKjZ0ZK2FabR3wv+F403rl
8TIIBCB2Ir9aSPdKvk4ZH+PAftfomcx61lOwhfHeCKbA20ZWJ8WJx9tTIuxKkLKSelD+gKJtTYIC
AF2K5HKs584a/qFljYdJtky98vMkXapctvwYGPiFH8+nB9pOvqK/Sc1KLcHCK+3Hwubajsiv5kZi
ooF53GA9gRVCZI3MGQI80qAzpYDSsJnEt/jDuC7ltqJZykAp7papUUcN1yI6KR8zk0iHw8pfQ5Ll
nUicPMO8EWdbnMRYNwG9DTJ/2ZFDIx71QXeyE5Dp7AvCOHP3AG/VSJmtN2Oq+ZfpGpcMWL/hIhIj
5BFLgG9SfgIzGBYuhT4J7cUqN0RPXZJTH9P6HQMBwmBI5OSZKj3e5RUkxYguxUMmwNtTj8Jwdnuh
HXWn5V6YQyFRmICK58r2uQOPekcXo/CGVH+tPhSffmfneEerYTdFC5rlQxK0hSu7No5HRLqhHkB7
ybJPvAv6aFB2Seq3ugl0+jpHIpMV+HohNk138MRxrQrX7J0L0UH//zxaaF7Qo8pghp8J1SMN/o/R
CavO8svZEzb+MaqnV/W+UrbmIXAawHX2Whj6UbeByH8doa50/oUygEy4XbyKWgiXkZawEuXJkIlS
5m7Sbakr7LTTKsFLyzCjsmiChooepV/V80sevK1BdWhhOQwOn89EcQ3QwqAgG6lvDaTpJb9PE7UT
aRB7OaNJkvdFs9oIFwYWllp0mXpAwnCVkq90FGIyH66zp4JSPAY0wDi/nSCFJtY77RvbEG15/XXF
wyyGU3vSlsgj++M0hir0+wzKIVpSsXC1NUTkyAj7ilGhLtuM/DoaQcG7xdsx/mL/+wld9+U48/kj
VB2ukr6gMThXKyEQvfYg69w+/IA1lLddiQiNDvh11egQ6ji/oULqsW0UBxo0zu44Zhqxdt2e+75y
6blaq2L88v0LWbQqMd4wOhRuVptLjc0HH28JrcOq2kZV45n9cQjGu8HstfofTLj34mgVWQw0uf60
wzQHw+yjFQIFgerKHX/vflFGMLdAZ9VeQYAvxa3g+Izd24Vzw5akJZk9CeFQSz8qSQUmao/na/N1
Dfyav46Com58DKzGh92fyzRV9bNoYxBx0VLjgfgtV05u9LHWif47dfCCOkZTKSXl1sNbKYYdVDX0
ZNEY3ITyiUy2UI9eK8leD/bUeCTKKHTjgRJpSs2X9DXyk8xY2MN5yMjsLTNIqdJ995i2w8Y0TLmH
CNohUt7ClyJnnD3XJmVUceuiiuRxcLzONAomBcag7b3N5iAKPfgJRvjMcUBnlxIg7PYuNuwW9rqE
+7zh0/c7TnfFz7NUDctla5hHLEUH1e7so9MSIEMGF86xezzocaYboFPKLBAUhs9jdncefoKzYbqL
XA+7DTsZ9d63oCg+fMSAI5Ai7nGLgZ46MIpkbwodCjZdr+78NBlbg5xgct3CTWZ7axC/4+vRZ80m
eMXdxE7dG3oXOJWkhqW1M4mHjANVmGWamGcADAptbQCNJZQqYaXzDmGPRWzxE0UdDfoZ7FagsDFw
C6B3kp93/CqS2jBl7GvseijNdkAIFNfytEs5jI0BanE1sRVxtAA8qy0FNZR/QdiCn77B+L1Gm1R6
Nxz3ma3mfNfAdlpnIabMAT7NwIyh23YUz/ATQ5vBvGg/qQFpqiNyE0D0zZ1otMYALfXNzy2LeUSy
hJwvR9jUKwdgjLzFPGI3OJa8xam6B0UWlZhYnp/yYnT51r5tcxYo9Xv1+VziE2dHZKEA76pUNd2M
R29MW3Ircw+mr9OqNcYzpaRL+t5AUdomfTGz6mky2Mq9oiJeN+UFhRcZVS4wglTGAD0GehaBKAQg
RKhDBGhpTWem+vtU2Xbq8/5RciPOygdiuZ+ClWYA+lPwb+cryT2y0pYMQjg2nTOuBIWs4KoSgd/A
KTLcL6fYkOOtqQR8asNvq2ORSNr0/0rDwDVNBcqHBsS8MaJl1fiFKiPXm+xzjDIeu2kzoR6Yu87C
yOdz7kFs/rihPHBsmzYnnx6++6GpeJTEgm4wRgtAfq/7N4WHHRZN996AEbTzPD+DkYlWzNRG5W13
wYAbQtjmcER8YpiCbpG2xBfrDuJ8OKKKLp3ziaMl03ISN0Iqn0emiwX3mDbzME4WjIx/zt1m8Zam
5diAdyw+p/aVUtziOfjGYGhgseFIR5NsubfEmgSZURMWTiCKhg6MbVkNYvwvBac6qQwAMEdeGDIB
Rlr098V4+QHCPD+ASzZ4SkSB/hgxa9+k7vr1UXqQy1x3rael4NOamZyGGCard4+0nsRol19orMaD
hoFbEZNhqGdsy2QKBDw72vqrs1P0NEefisR+7EpW/zaZ+USV6h78cfpFfhwasaD87mbz+sNWlWmg
83qyySi2wNzFLGdanyHNww+Hz2uO39DXpQz1Xme+Zxc5uzoZ+J/ej3ruU80lf3CxCbDF/REcoJ7M
pNxmZYvz/its1TW3kLsSYrLjCbAEICiD2VHypslGfbaUfAT5GwEdbd6rxKqZ2wLIVZ4xppRj09XD
fquo/V3DSfTf1NHalxjLmmCUFo31W5hdoxiov/dhIsWriMLua0Nbc7+0y8muxEQZSNsTmphv2n/O
D0nkTEh5aCkb54jzftw7i2tG2DyDtwz47pRNiK3n0y5kW85i1fBgcZi//7jOwD8ObEj++YagVHNS
r0Rs4xhJNOLvBFUT0+deghAfklEKqkqsrzDTNohjxhm4QJZOuO4y1+AhAEa4MioknsNT9lDMWAk1
LHu/VIKay7mq7HPqLEuC2YixSmyrMUbSioBL4l1vnEOnEPNuI5czL8AK5uRQGQFzIWk4F9bQTgwr
CZfaZYsju8dJjGfrKxoZVxqUSFoOdRle6oZz66oELmh0XbwnFk8mZrtUtaYRY/DNN3Jk80szWlZR
idNvtBJRsli80JR8301XAdhESSLubHeKIfZFMItXXLvU9AdxBksnXF2cf07cW++zuQgA2H8Tbo1k
wn5yJNZVjhatNhW/bMFYFFz2FXuzUewU51rTLOljbxjjHNpss679GL2X0IhtkooqK7L0uqob1b98
iDCCXq8wI6222lOIpwTcMGhZMV5uHMzXCKL0xmmhNbQO54ZIoBSm0f51xPW94pFz3J2fzaYQphTm
22+5x4NKJmtNS4KQhuSTc89k7UMxUH2ch3A8uaGg+W1zcSUuT7HWrEulqNsDUO2wtEGl7/N0YkmG
xekiCeQJxiEzilWl/XSwpXrpOmW7nUI4KHwd2YMYda3nANW5JNFoag2M4rVtwAsKyLq5cldBVur/
PdNizAzmbFttuAkcBuLjFdQQoa6nKJyhTkFMie2NlQKZtxjxhLaQ9/CKucOgtkO6tXyZrDdFIbBI
n/HOqOQ4CJjS7HLmVUKKCxd1thVAhjrDYXJ6abHU/XrHR1mYDENjycK1uUdT3l2kmIWEocl0/WT4
SzNNLZ9ZwuHOiqaZVC1QzHCgfsAhl+FTnBlp1AqQdl4kfzEHp2qouMw4nChYg5fOQ6kGSJKktR36
azhlZncUJJJVqh45M16A8B8xc1f1LL5/N03oG9FFm4jJZonPAE1FEa4hFWUvjCQ/E/dVaSAs3GLx
DYue4PWRZRp9GjnhBd4Rx05gLDQ6AX2/oV7MQkoN1pghyEzJ5eoiltGvOMFMbQS29GFY1yMC1BwM
/KKeJV3UGX2ro8Cy7F2r5PzMgyNiA1LguMv4o4xmGozQQdOM1hmDt9Cok7QL7i9Vha5oWoVQ5FFy
x6qJypsWSDP5fDcxEBL6u/VCHZAxTPuGStJXo64FahpuRoBKqU2dPZxN1XCLtxr9joepGFoe9GQB
EL+99GNalJ818uoSR+l//U1ONh/txUyqjQZbFlrgtH1XrgwexvNkdQPkh6ODpDWNpsMAHGWyVGmX
1kYoMIFk/PKbpeQ81Bx6Q0Z3SvPFwyuNQGm6KNnmj/1SoJ45YYlc/ONTDVyD5nzB6Yq4uKpJ858A
r+a68XwbHoV9ArJ2Sr824qTeOiRcLUWYWgYE64MH1Ve0xmjrQ/i6dsRNJxz6+1tSBJcpZcuq8xl6
LGBiovQN0Pj5KtHKVsdjGq2k6H6EzoRIA5EIk3NyDR9nE9VcQe73zjBwaDlBrWJ4JwCWYG5FxhgR
gh8/fmgV3MkizKkV1U89GStS6fGzx3HUlt0jI1W/HNeZLG1eAZxeXiS3AvFjewSdAGYrhy32ANNa
8akI7hSaESFw7XSqp9yd3GzYhpZLrY4fvUXqWHfQYw3fC5lJw1Jt/mWSE0Pprvdl531ANzobqvOo
wQKOLDPTJb3zPHD5erp4UiuiUW90ysWCc76bIKVlOwpNXTqWOBALjnhhfTrQdhxM1rjXzRU5EipW
NI0R6ukAL3a44TLLBF6m6VZF8n/q+14P35TDRi329FkmVo0/Rnh3zZVBjHHiL7Od5dq79G9M2kmV
/VMwIyfVsSarZwkzM/zrZGFAHzhp/qxC466mddl3FuubqPfS0aLS6hN9o9h3MbciqtI2od2+fb+G
hPapJPS9ilpwCHHa7BG8QOi6d+2KE7YgPw+bKUAYczEHkq/2LEaOUBZQhJrTa070ruFdhoAT+U3A
eT+J+ktswBKLZYz7/GglYIQ2mo+kW6Bauh9ySoYua+aEX8wLzkIwxgVs/BKXZOQhl9Gy3LMfgag7
PkhfKI6+UlMMa6sX2D5fR671PvoofDh2mCf23GPen99wUYp12dF67I5Atx2wxi8g1zeVgEE6X0He
rtUrgoJvPiK4DliteQZB4PP2Rj+Hrt4Z4g3Fy2D3mYiY4mNR/oHM49uD2bTC924AaJ5bDQ3llfIe
+UZ5PRdo5ccA8C+LnuiKfjDfoH0mnDpdWix/cIb08GLLZdSq11tQfWehXCm3oCW1rlkDlnb/MKXh
4SSs628xjTsGOXuyZ+clR8cFZy1tAEJ6fWGhBfHg3E1xfZpAzvlTCKqJeGHK1C+2uxaRzY1EIN0c
G/oJ42R7UPyG/W83849MYjXQ89Ql+IVuWVducSW73+qmyUKDK6EGWBnpdTjg1XAshk79hsDLZhnM
fGl3D+JxfsMLXYEyoNaVGusQIqb3ihsb1G7T0PSdia3LbH+LyBa9/aAf95dLWY4gUYTGa+2EoMXl
uw1BBtEOICgtQYTNW/8nJLf6Md5QzXEFf9Yqa8jx6UxW775dG/9NkHg0tcH72PR+mJB3bqFyqdW3
MW6uKw22ekRfox9BIh2+l4nb3+1YFH5N5ZXwo7jbykJV4a58FdWOpUhyuNVLkI5fXGlKXtOpcqBB
5kq5w/PJGRXM4vCqyN7JK9J5l4aQm6oQEgHIJLAVfW3bWhFy0tF+qqUXXdq3j7J6yHRicuwDMzDJ
vtARxvt2wjSsHIfEnFgSCRH0a9hvXCII5XKfXVOHCMJKmA273v575D/AHXzc34YymMeDe2mCJscv
00XU9a8FjMxWac1SGmNCTcez9QFs76rsz16vwD0OP04hOUqv9uHGqGPgkROy103GADKWs2qL4fWC
GNMnyEp6uqqe0a30CNjstDPmspbpv35T3pzUYAWfryScEhngKF8DnacBDB+2B6pzKnKYWaxlVRkb
y+ztEANRc4W3Atk3CUJU3MPefhBEf2H4jMwGkzH7AiBj5aDsXOE4pHXeHNO+5nkl6HjxT2WW9fPX
6FqdePnmIe5f/IsRFleao8kEcL8y5vfemnBLdhJeqF0SnQ8+53+0JpWpEBF0ne7Yg+89Z9eUSWA9
gUn7SP3cSpu+6Y7AhB/uTrBYjM3Pg8jheK+YUvzHHtkedVcc7h/0V5yi815lseOJuMRt7bA9+IQh
PsFj4sBkEHPJLM7aZjfzXqXfeVrDCxsSmX09bxaviL2bm7A2kR/TVzbRJZYaWPeP++kFbBH7jmFW
2wVmCDkLHAbsRtRyxYZQGdKF4Hi91IimX1v1eXcYcX5uTaN/jo4VGbIhUPfyY1f9ERPnt6esrOmB
7pqs3A9KehTy113sNeP5oGMFCXOGfdmW3Z2HXugiwbGjwyUkun/DDxBoFTwnCZtb30mMVsj9u8bn
97OGZBAdl7W42CxrEIu0pzirI4D9wBWGwQte83dKGgoA8t/vHeJon0hMo3dlPBGUaejCNiljXKP3
mh/8cMNkAW5q9DrKwufs7mvAgpHf0hm6k1iHD9Qo7jfeGFTQjiTN4aw6kTjrJ6Z9kZUhPPcocynd
/k1GYq/xljV+WEdL4FiHSRioXl5VScz+1wHrDKSHW0i4YGQlZXrkxlUvducLGtxnIk41CB4A9zHI
YOoJ2itiNl03Wt+ikgBOEAR+xIuaZI6iIisdnSB4ggWJzgQK45EXt3CDYZZhnr9Vkl56SngiHoPk
H1lH/zbni1xoQyHuZOpIIz27MvY1Hsnf3tq4S5e149AAxWJPGOmUXKS4EpbJdR69zDDomQR6ME+M
qYCKsZF32WtwkWmZ+nLL18ZddKk7+fm5+lfnEWdIM1W5yyauekqMPhUn9GIBr7sFZLmZ2JiHe9LX
3GbiELThtx7Gssw91AzXig+OK+sJ0b8PjTk+fbEejy9PyIMD2+k4959UjRelCiFOic3AebqX3veg
fMHpXKDHEK5WUqSTBmRawDIi6Rr+RDVSDYRoCHhuX616SQdR0EpKzyj7+RaAZgWTOSZgkJct/CUX
9hmm92QMTgdfQvmPw0m7MFEJT7Z8VDwPqPEvBBtjuSNmEshmLH7j3C/nqStIYro9EszI/3+sEG3m
FOPB3QWEY85knqJJXpSI4XDj48Zv/Z5JK/IiK+iHPTmXYvhSWvU6anBAzHVyGswZ3RGckB/pD/3H
5ULhgzd/7aoDAfltHItRn0MNSLXke4f5yu6CBxpxyYeG9DexCYmV5a1exDh0Ewpt1yRtxLSVCkQM
UVY5dm3lrq8KJVrDxNA67SajwIZrfUQer8BNPv8wcQDb8DhfSj6SAKITFhf+qe8Xdiamra1tNnAf
WhRGKDvg6h5pfzM0634FRvaUBXzXs0G55IQe7P8w4oMvtGUEjbZXfwarZmWqHmxm3iczi68Q7bml
9yRdSqDgGWmeod3LZFwEBUDGH0w3kDvi/NaLWmz1DBP5BjL22wThImzFKYVi7mMxWZXjp2VD+H4j
DhLE+x/O/2kXbF/9BWo3qpfkEX6mvNt/Zh3rJ/vd9qbVnCD+hg9IylnE3mbmXCzkwOHlEgRmIGfb
CD6QyHecUzYF7CGWqM3vzeRWhBn9D31oZppIpbKV6zyaVFwS7/Y6XQkOkDYQCWgBpZ+d/ilRiTJE
WfFWSjpi1RFUD24dCl3Q1nDQ6U3rj7iCp5vSr2doImZcNCplmMz2O5IfIgqWIxAZk8ND7AI7JXiA
8M+MZUdNy5L0cXLdK0pYKVywQp72Qk053vXRO6G1vXa4PkLUUgm2KDag/7sOc1inOpoe/RVFPdrV
JV2Z1te0EVJzIck071M5jmIWUy6pAyZDqkY0ji3jI0XrEHVnh+oY8saSgQWk5L3QJSfPiVEMyVs6
2Y6iVKC/k+6iyLh9Ofm5rlc9grJkdSq6BRtVtHGMx6yn+tvKrYH6l7IAWwa9vmzL6j13sQRhdjrX
YIGlRKEujgsa6jKj1OKHxadIu9fys5ovVdRC816y9J+UwBLzVMDSME8XlZn0FGNJzhqHVt0r4oVC
ekMeKh1EEyAivRHXRa7dNs+xMw9O4nnSDAamYWlYAUbRWr0GB1IRgsKdBS7PHNgeRU5C86ptgn0z
BCeeV3G9D32Zhx/1GuPI6nJu35/KQ+U2ZsHd6R03LyHX8cw6UbgCTyPn+oqwgKC0QDlMXyX040kH
ibYrlrVu1hrIF/1veTMd7WngAcCaKH5CaoBeFW4kAd8voUzTpFyAAk74y0ZR4KQuoRCGgIM7bF7/
j1G/TnDH4CcN/KIv/KT7A7qHtWN3A9mBs5z/jZvOn2lArZSc23QVdl+iXsl1T7ABLxyHUPnTythl
hALtsr1aWIXoy9gLH/ZWTrQYVWkUPqKkxF/k9IvZk1oZz3XrqFHM9Q2KC+MmXebMbym1jrHw3tkQ
OAp/IclYzE9aewxvwpmYNMdoAWUgwzj6sNU/7Lo8bc9+fNZovpE03j4rXjFHpg3x98/nRJ/bnkhw
LTEkrRy4SAL4aVLhcubsofecdW5n483a/iWo94HKkoNC2cB2pkI3vZMI9NrZjRHTiuy8vpqhdztD
T/vBGS2gyFIOsVFTBGEVlz05Oi+auQSoTw3FyaJ4jAavOUAcROUJJS6244lwL5h2gz5k+Anb9tt1
OE4ZJuTTTzgCzuu4qjL9YFY5CxNWnSjxi0oek42I8OSR/GDGoiRzpSfEhgvftc2gvVvgw2RbqytT
VcqWQgDsdEWnneOKHwUV/XlaIg5qqOKizWVmpJYMCTmUi8wu4dSW7FrDC15F++ASINTDc34CpcMa
8PHqjpHtVtHRvcmdsu8SqwMP6yA6arbrLHUVajR0DzG0GsooPIz5qbqd2O2x6Ben2vrdbqwY2ceF
R07WQb+6w2osVdZUsOFBZA3EjYP3cBlSfkghbm2w8j87fvflfJYRWj2J5q5q6vOWoSiNCotkhrX/
2qGkYaVVe5x3mBCVF9HKBSUTwi5vJ+IBHUOBFyeqL2xzzTDVqu7paVzyf+VbZ2DCqBhfEtELhqP7
zOq07x4Q6x43FtDeV/dkcxEWp+If8M/gcvGbtU8BIstZPH/yMaYuWnXlc+Qs6qJjCIwcwOyxRK3C
Thv3nPIZEXCaT87oR3nQmoChw8xTfL7qjBqF7CXz0E4Rk4+QKt7/Q29x1fTVQltXJag3RoNXXzZR
xbXcDLT77RYZtP2SsAnX9sSCesF+rNCr7+npo6rbZ95NJFDohAYLg64po74i97nDl4wz7aT/VgLW
CPs9k8ea+0KtkBTZljaw/Dz1TFeJEZsL3mPO5KppsEwQCSEVnNtT8lyNMpTAqyhjtmy7KkkiYt8E
tQKztpSjwfunbP3+1ojKmdfevpyPx3x4BEEtHIsooVTWf3uL8nwsTmKzmGpiWkkWcstIkoFHMWhE
ybQP9+yH8goc/qb2CsgsTnAPkhBc4GB2nkBmIIAAB5THWeArJsKlH+QcYlA4jtZz19/a3J/ChFO1
OT8fSME4STXsxNguhEDQvg6fDumVRFYx+W+XQFqMR2f2zwB7/6PnQPvfPb8h+/nkifiJbI4ZKOYA
gY6SmwB5Ldg1chjMtYQNd5mUQiPY/CjqNrgeliROHjIPmBL95yWcCivsd1zdOlX0j1op6ENmBFxF
gh2G5zdGSDDS1uclUkbTXg/v7iPAS6NhXrb+d5UuTfT1kx3xb9wm1Y+WaJtCzkcVUrN/+eJGie6B
MIpdCECkMxfNZExj7yGJfJgCUwtbc5AjlnT80vmQP9sFdICIEV44lwpfmEVKJx41tjl+iGlhcNn0
LsI80xrgSqkkwweM8pGmR+vF2nmRSBGzXT+OHbcCPJm6wqwaCipYbU6Wbb2M41q2zZldfxT6gj4f
jDeQUh5hE09wMfogQdtWjrditcTDeM+qenmww4yWn/2R3mC/hyxjgE/29iUO2Nem5EsBupRoRrMO
oED8eUhowuu0hLtIms6Lm2iHBGArBv4h1d8XnWVM6i0vlRMQAAYVgC/6n27V5JVkm5/JHRBjKgD6
BfQMBuWn9b9gJ3g7xvUxhaidkUDJosOdzEX1y9mOhzQ3FfFM8Pn4aLInjwYIdyiFcAKaVXLkMzfN
iFZKfhckV78K5QcyIZXD/aX4X712dTbMnl0PZlI62a9OvZmidwnpsl/69iEZipykCkAjFypjejQ0
TM7IZRMnSCQhtfyThT2PLutw1GWjcqMrArh1InmhBqcmH0RhpGUtsCOyTO1dI3ZIx8Waw6t2XgBW
MqUSdwCf9CEBS5FP1TMZN191BDAjqLv0gO87hNYMHnEzBL6Bsd8QKIr9UwrQ8dtM2I8QKCmusGO/
FlA/412RGYJKANzWEZNni5XFUK2ux2fpiSE4XGHlRipZb+cFAX6AWJn1Xn5ccnjnWb2rDQl3TKc1
QX4H5KVu2hXM+80Wkzufwq7rHgsBuR5DTz62/7nwU8pcocKS6hrWrYQiP/gKNxlRBLToBOp7N06j
5CYIcEqgsdSucjFehKc01yFHp8J4FFn7BZnfNSPFgjsv8LGTdHvDC+iVnwkxCQ8SJS2hHrU+MYHj
jboZ+kkjeDVO5qMS9JuZIhZ6BJYML8rg+4GCiLA0qruTcYV+nq9EdEs37nEhvU/t+r9j3WteS6gu
M+PY8bw2wrqKKD2UvKLIkvmCn0seRIrujw3gCvLCipagr7LBQUqiNi3T3fgwmWK6NzzMVld6WlWZ
d3ai+SlGHI4ZE+OGalW+9YFtxkHZeODPbiozHGbQu5dXj4oIDuCMrWMlduzEgweIbuUjOZiJttEI
GcaT+GJvKIBJc1T12JHMkofNPK8wMW2fSP21NBySDTCxx8Lh8Ne6Vsm/YNocG2Nd9jbZYqifM5Hb
2sWV7OTbtY4rVINeigPzeUgkFh4tEIAQCEa7JBriIiQIbnDiOMkGvL5Ie+O3x6mjVv4lMx63lYRw
qu0VKJNNSWgoqFb/cwLFHFALCNgdLj1dCfW1eM0hAATAq1ZSUL96+hdFg9BisinqRNCb5ElYTHRv
dI97XyMofNe0QhlhKxAyTaXN5CDoLiIjUviy4Qdl+er+1rcVMXYgg7gVYvhfzAXTXnlE/92JZWRx
eoF2ku7hxvQZIEhshOosa1vpND1tCtbdOnfk5mjzWtaS6cChRixb0ETEEEmFCNBpS036bxoeUIn3
oAl0J5/62W+QN1Swj4ZH+H4Eb7gMo6o6C0c2VMsOgb6uMQYdtXvDzqhkIhsVNle7yO+liJcTc2ir
Dc8CV1MTEU0qQiuSlQpk0MxYWTWPpBnAZ3NR7bBBBzf3Hxf6uSjcZY+S+Q6IjdTswERx74aiC7/Q
XU2RCnwxDv5KB9gU7v5JkYLg0uzmtuo4j1UCwe44JWByVn5SILlbalKVa0DgFxnbHtu4BUEL2Ylt
NSjx3IDbDarOCX6w+qCyaLYT/aFQKNoof5VGuka7OJ5QrrbuiY7tofwqDrAI8Il2dOdPwhNg0Ira
jTT8/XU5xFQTAjBO6iDsAoqAKJ0NN60jfGLHTh2ToXRCejMnyOfGRvxhEIsBlF6VaosQ3SpctUz9
PyAOs9CS2vhiuR6rbZtc/RAK0T/+w6yUkXeOZ13SZfox4RPXAwPYbnnYAJUFS1n+cJbzYRCGCQld
m548XZQUFPpu07kViFHmby/n6Jd2PtBmfLdz3EMm+tKE6HBRzN9RFYYKaDWL59JuTBVUaUfn6mt3
h4XRsgM0ki28U2R+cYuNCT2F6df/ja1yHOz/srZ6kA3BKqOcgT9rTqP6cXhGm3hmztpwGoDM2crk
hCl1K01PEqVw+lsHKB+nXX73BsgKp0t76rUQn5IfRbyCXZxJZ6VSSgz5ddHbEngW7P85C7zakqPf
FtYJ5ZH/0N5W8HKqQBuBqIwODD1glLfgcnmpg78oIMS0U7Fj/eS52tGWVvlkBbwVvL+YIPd8D2/x
xmZQeyIh7hhZAF1reeqHY4KvsCMPWqy+oHmTsFNnNkKz/+W4y+nw2vwqnMNeqPhur70ZHV+67AeZ
SLA0TF3DjVpKTrWB8f4biw277Gt7cDcE00jCs4wWGdOhEwUKTwioC18pl5BdSo9FULRuxs8Qck7Q
QfReUBvWYkfOS9IYTcKZoc/jVrJErRExSWAt5VIMkGA+HIx/os5yQpyurKSXnOD2o54fHNLzlJrW
hFk3cZHXl2/is/Pw8yvTfEH9xSkWy4VGvRWS6ac9F8+ewPMObrPXo6TCUDTga2uNljtl24ah1yZS
whSGOV5Pu1GlXA9iIAPBT7m/zmRSd5riqwSrmExeTfmwhx5ZjkFG0yOGS35wSyrY4i0pHLNmUKJD
kqmB3tQ+PkBcngeWTB52EIm0jlPIzOC7wlE9C6TAi2KsKT3obzvgwAOXx5TrXiAqT/IVdeW0J6PR
Wz5iVfC/89ZqsRvawky+6kaRacnWWICDr9xCUhb9LZMJPpPIHSP64Xcy2HC1micHzIlLHANiF/1f
CzFzLtSosWXueOV44o9WTv3Gc/JYZCpchseE339LSwA5ivmwFZbwdXs0jLapOw1xCv+6JBt5LcdO
rpkn+NJ8b1MBoh111o2imHmbgkayzOYECOdG0bNpHbXY9aMZNUkvkZqcIFEvyJ0ScvABgiCI9xES
ykNylDfEkzNHVz2LpEliVO/cN7NY1TUeTY0gHEQc4SXc2ihAkVLnMm0zIXXgwgSrriqv/RrbESme
UkPN/PQndDKWiNulWx7OySksKvtHSC7q5c4tgNYJvbECnCEVWxg7YgjCoj3MMmVbUl87oIvGk5zL
3hZ+SfHCBMfsiAgb57JLzT2qAXbiQATe5B9o/0O6/CqrE2XAEA2biArxpuAMn93+Nc4i6i194JRr
iZlEybfT7hhCyGNh+Ugq2Sz7NeVWIVvRPjjDI4N6CojB81imGvYllLXX9XLvPjTcidbYFDHFh4wB
B1OlFvX5SkcUOoIAQ0+gCfBhDVdwW9d1u0k3dR5pBYXeXsWtxs6NobOIEOtutbxIFJqAmJJkaQ3k
Z6KArWj6cee/SIHwI3KsccC78YLOXDGjD5Hlzt4NIbhZCH5veWD/nkrA2njxVkvCbT3juFW15CDj
ls8TgdfyQUkj6MvUYLZ5/9UATgLXBbLea7TlZzOBUVYHEenSdSbGkrw99nyqPCR43j+ROXbQqkUF
MHJINiMYzI+5QNwuPSqiTEwsZTso1nXIDS5boLTAJWgo2SzktmajTeXhxuyc/hAIcF6bhfZRXVYg
bUgl6wYqaUBg+aKtow3j27QWaUEahbLdPap9265LB6X86emxE28p9JBCrnj4bkZZrG2X4BThLxvW
ajPTUsevow7cLpdn9lglRQb9bY71f3/HNrLFHZENyF3Hy7SMeeEH93r/Ma8hhwsz7bKB3xQvP8Qf
QuWJR+1xJqqiPDO9Y//xEUVxpxmn/QhMrJsWCxegW7t0nrAPf9SE9Mxmivi8qPR3n4peYoK+ik1c
k4DTKIMZ9Or1WRjsiPso7uuXJVRbZZFOAaeANTuvt8gAdjGnK95C1oBd/LrhXW9Cj1eXwb+J0oR0
u75QAUfIl+NIuPBHdbW+f9XFi2TxsqGH0O1uV3dj8gnU42Bf+dF9G3e66IRB851P2/s1pIoCWqwG
YeeRGxX1oC/5SMXexj0kQywKF14YzfmEbdnANJVVgiwnLZbkznNTGXTc7K1/UM88SMYeX4cfycgd
FtiUOiVm8n3VD+4YR9zwYwKB44nC7WRLiPn6Zm6wVs5D9l5Fy19sFCnvzIa/25+pmPURtpR0DR3G
2CEC+dYchVzA5AcW1b13r2DXLjBYodRTcTxEqbuaw/f1CcfqikTBfAdtV/tkDLt66k0o48/Xm3IG
dSutA0rSgJj3qcFtTrt2q6KHaP/u4h9kqgQ0BYP0IQOXGwfWzSOsIAh0sBs3sxGm8DgR1XTslkAm
dhiE0ZDPcKvcko/wjc2+4aKTVmKGEdhlwEfBoAhFYDk9STbTuDYENhpQYn9Bu/7eZ+5UnJh6J8xe
z8CqfppjeSkYTYI8vJaCewu/yJ3BGOnXdNQclrTs8iCpv7ogkfAhCKO4kmUA2gBy5+YyEgIgiuT5
6RPw9P95YrkKKWnsvwy7dOr1ipuzyxCQpxE5uWkVPMUQayFEysZHkTZLRY8mONd3AxcOQzr2aN73
jXcr2TRR4dI0mjOBiF56kjPVw12+EsPOqDeabjGzy8JoqrhY5Qjy10DbdP4z2I+JQAZnDXfl8+it
ewgPeeGvIj0VyaFsOJRfaiKjFMHrmndFbKur4ndNDS6JTdByEe0SEKITCsw77NE0QIB41Me4oTdJ
lpYxwqfBDI6eRujcw8pPapw6bYhgm7+WRMhAOvl18unHVvhgeKDTeMB5GCh7TA3tGS29oZ0jxYCT
skCVC/HI/h5iSziirCnx0W19666Yfh0vNvmS7Qk1cENk2gzNnXDrq4Qo2ejoKxOvLJDgNDfdx5qF
UUBwde2dHdJu4mal8xlRWCDRPVSReBBUN+y1GswEPK7Y8VPz5wkOeqtHV0Puhavsy281iPBStMjH
ThI6h+V6goXxm1Qfh8p3U4W5UDLONn2hWUbGgOUOyroVcmAvQ0c1v2DtyBfjNyXCyxfI3fgY292A
GgpLC/l+l/Rf8/rbqV48tFKrXDWqW/axI42kDr5RQT6y2LDN7d13HdzVUCDPBfBPKZlDe/ZLK7Qs
xoL6rck5mNwlT5BC9AHB+VOCohzSVbBzLzsU+iK4p/qhfvq6QzHhgzFCEeMANiKn0KDjvPeQFaQ4
ihcbMWdYeMqgQt6DG2ePGRfVB4bB5g9DoQ6wCev2RhAUzO18DrZsK8SGmIBulC+wAKEm0yrm/xRj
E1wP20vDW6Sv3MqGUZSH0OCj4y/bDC/KSXqoujJPZsHJVr6SacYmeDBZbN6+OpQi0n73Bet6Ohnw
UpVM57WH8yG9ni5pITr6UHnDpsqlp2EkXCIpcYx7vHD3zh8Lu1idfHSbxv0C22jD30CHgqxozg6M
6urWMhmkQWFcL8Clv8HsuCTQ5LK80ckg4l3/VaPFRuvAuHhzmdVIPvPc3b7zBEh1j7p22C4ctfce
Ug1SASIgrB1XuzVTCaarnqa8UTLIkkzRqykE7JWbXyCtR8QDVUCVNQYRoTKwhhMU2t0HmblbkrnQ
ooupfHAwV2hYu5pq8uN2Ty6UYSgUS8QGUB8UTfuUKo/3yNb/7MBsuuf8jhNsh+MNCqOp0wSzBggl
6Q+CctNnM5TyAyEwaaGr6hozppbI6xoZkJZLVp08Oz7SOjC0iNZ29Yg+s9KH4dvkZoP4ZZmq67ko
gGUkX33CoXHfaL21r9nYzGWIdFfNFAXgrhC0MIhsY1uV7vt5rsnOwwxpqcEc9Pl4qk7A//XKIgHB
WFlHo0XPk8bENkQdPmmg0W1B5/2NBFV5WQgbkcUVwGtKaDssTwmoAFTvYwCJ5k+l3IIitancxwpF
Srci8gtr4QXChBoHvgQikPkzmNdS1I3UCXdtvnNpHtTLdC6GjfT9Wmnp6hn26B9xR5B9cZiIN5ig
kNdzXGECbaK5wprfxo5WjZU/3e2HbUhdd5PegwH6PGeu8eTcVVQwL26VDYkUFM0HaU99lmaCJyac
Z56XpEus71uqoJrP2Ei5FoOq66ffIphynnE2avHKpx0mtQL8B+mHX63nXgx5pIc9PKuXNLWMnwvM
jx3NLBZvGy0aAbyqkbKwIs19MJSxyCpjkfjHJ2UB+MBKkIdNIOOT2ubLJ/EW53A7+vFXpP7aAuUe
oQ/Rx2Q2OdAPxsVWPNLI3acZ+HFtguvHOt3MDias7UnQ4CVX7Xj/NG1bPoDNG91jBHY9yoIb16eo
4b9RiuQJupZgrh3eUJBQIlhSwY498vt/1r/gkfaYMLhZLPb8T5Tmqd32GkIBGDKy+h5PwRE+cgar
tqdW46iMhVdNK0FDDsKWPKaLHTYKzr9gaIXFr72ZqLZaGWCfQj7uZfh65cZGciWWhKhMb08LDTpF
MHUU5a7jdReCD0g9kpQeHAbAleifS3bZsYYyOSiO+Sbc7vLgeQFtGNzKjouXHW8dFnPdh8Ni3a5W
wf3t1LVrvYFqqXFdrUT+mqpchFiqHXSh6nZPnnbXgpKIZdHIWjnjVmLDVN+g++xYW/u5cfFm++p3
ZLxKPoPzvcqVSTv4jH9OqF2oGpv7jGaZYPorZnScjfY+BOkXZdJJrL8TjO1P59GqPBnzLY7WOUeq
ghidR7z82vZ1OerV6BBc8j0ZVggChCJc0fFM0U8fn6maaBHeXZDJ8w0xHxUm50tuDPYlZi6EG2Bm
N1649K0tZCsRpSFpbz8LD93r+PYJKV2qMjYvfYxWBWAyDzmxbgYjcKTamC16SfczYZQ0+555IdJq
e8c6lXpChtyZbRXQk9EONC2OYyemTK+N5rBkCrBTmXwRtqqtVwaTt5XiVbgQTIn0FQ1PMMrP2m0B
WApmnkrV0UtqWpL45JkDdOMXL70jeODyHPXgX9Lf+yXFesyZMpJBJGw19HoCvm9ccQSGITpOCZY6
j4QjuRzC3bGyrkVGkrVTsUVfPlv427ih8Xz96thWup2qq/RSs+/G/toXM4sgEE6ftw/+r0bixKeO
0UgjCSnZw+rJCR9/MdklWcGVi1+g/YqBjN5jwe/JulMLB95Iq6JW3xwx/OMMMvqf1YB3W92Y14x1
eyTkr6+/x6e1wbfwfeUGjVT+w40fQsLpIjA0qHnXL0NpzG4KWu6nXmSkAYJ6UROfL8NTW2YuzPEM
NE3QqCvqnhUnDaM3t8U/k7motseIKW4IRZD0kO21WiJ+OK/Hbh0dDq4ZwkVjUHgf6tiiC/sTXKzu
+c739kHxOcLOQJ/dZqvI+eGFBTh7IlWkA5P7/nZpawHBkoNZ6IcHX+u2mpyVZE27T2A6R6kvY8PA
PdqbuYHFZktQjXoHYfR1BEvG4iWFdfE2g3U3DErZ8qLiX543MvSdpXXyQV8CitFtXVrL7VQc4VWR
4Ood80Ll4s5ALTtBskUYS+K+v/AP/lCBHT/THZyILOXRA12Ae/cyIR6jgNaXPMa6hSPyy1FG0KGU
XoI0n3oQyqkYi8je2eK/CLNfiSl+BdUN6721EL/a6HmREVulGvt/IzJmNRm9wWi3l61TZQDAzNkx
+AiK6IHeaU7EVR2124rWdQLa2W/05KRt6/5sint6iGt70DNz0L+kWQkcoQFlt3hdqkqWG8arpb3H
Qw6QmT14AMYMfujH0l78CbAQeL9mJEQtNW+uPp1mqJZ2XCxO83RWdVEiPsBMh5OagTU6ogQvYadV
/KfnFGnWpT4gzk2S7+HPqmLF8ZVkCb50W5zu4Z+5NRnYpRV0VFKZ09m+AwPk32ZncUKASfyCsRd8
ykYune8otEM+p4Pyv+X0+/ZZ+ZFqqyz/sFGMPefFF+1B52g6l02L9pXLHzguseBGaeiEld7DLfSi
jQjHtURRzxGM06+5b5jVAIfJ+KfpaQNPxFgCtwzrT0fllzRoH40FYIkzu+6U0Dh4vP16rZ2A80i/
PWhHUvFTCaGX+sYNhV8yjbYTvzNhzuoCTUNm8rbbxPuiYavdxCxH/P5socq8j/SS8o5m0UPpWKcw
+CoPOZzueJG6Cpj7HDwf3TLWyQ9PytzOB3Stdox/lgmtRNL9P9kXNNQMPUgn0/tLU9dumGGNzqAX
qNoBpx3P81XuL737EwPzD0vvk1KTjvOfdS18teUs6T0+A3JujvnCiVCUHdKBpRxWzQwSGqOGrm07
4B/1rkhrzcpD5IqGILJ1eaakuSOUXlVDzu3RB4u3nr8UhF399RRJAtOglOoOA0P37qFbh2/p1ws0
ADyqR4byzyIzn0ICSHDVIei5O9vnUZde7sa3RIMM8Qtng9oX2U5JtG3Z8NeY7aqPi8hDEy+Eo5Rq
FmcBCQWnmVFZnq1eZtpmK4R9SgF93vbPmu/N5E/iaZsiHPbi3O39IL79Hs6r4loF2yXK7ZQsz5Ml
K0w453X+jYHHqe5fderiLlRlCK60KxsV8otCn3LcwI9gTPxfQArbeqapjD1nAipFXV6cdkC1IqgM
wE0B7m/TeWG0gyjKFu2Uqb2AR0neWNiLtFSuY5lQJeMSVgvRckYHdPzl8bL1wAe4qgzi1qa1zUNw
FT3+J6SrAdWLPa7HjITChMFVxIlunM2XaJnanper7aiulWrKoxo76bG1OO3xQWa+Ebs6xghgaLid
+JBR1B8oiq321FyLNGspUivfEcy9iksZ8+3LY4MyhuRxB0sSqHw1jK6PIPxUWC/dwNBTmgYhptDj
F92yCjGnabqBjhdol4Jr7pvSxtkv+0r+TM3UnLwnmG3gfOPXeK4giD91Al6GsiRmt68w7WbkGG1b
vnoKpotV2WpzM5u1bHwV10JxFslrPEDknRZKR325+I7b6Q/eiXvzjb8KpdDn6I2+633VyixqH29Q
pa3vWdYys5eGMCxf6VSlgLfIKicoy0sNGUiA9WyDmgb7MV0INUi9czQMhotETyFHn1DJCQM493tG
ygeHdZWpB4/Q+4vR1eEKRl60puL57HnSCfbuB9Czq09zAqhHK5/3pUjm7mdxL1mJwgqrJIbJ5Cjt
aLilbGcl0jXOxU86dg49lE6eD55z+gXgjvATQ0WlU5lKqjjlszeDN41lscEemmaqZOYoJH0xPtJL
Zg3F8Sm3UnD+oLfIKS87asiX093WGbfR7+HEM9KIv6FcSXMMMKGjpcXjDAbYel1+1pEROTcHKJ+a
dP/cxegiC33ttAoEPytCEPwbQga74+dT2z3zfY36+IYnSTdA4wtmiq6nMiXo20kGgNJi5UbHfzHY
8mrwiX6+WJDs879HjOvECUrih1CeSZSNfanHL30Ig6I7WFN0icHKPLzF9zX2BYmnLNZo1+rtkNQg
0xQ/KdoYxZqu3yAXsT17l9WVoFiQw+AGnU6sQsLQKWHeJP9j5GNhDlHlWY7voLYmQR/uCSF1ZuOH
p2BzzI6EXTUda8ZNP4A4DrW1nzXfQNGIVDr+xFuJyQmA6aLGb9Mc2W7l6r8yL70DJsbKmybvuT5l
Rk6AhciYzmozyQn15jEOnGJO6RRZFSU68BmV9dV98VcSDL+3UG4l/WQI9PUbQNHKz0mXgLcubYRg
kIkEP9nAgKABIrlCLumRJve1qsVhyufguD+OlvFEK/ICNQPvgxCwmbJPqgVFAc3UYOUTrfYFM2Gf
/QVZlkKXTn1vHBs71+3z4rRELxdRbKNUvgaknooFPhj9BiSGQb5+slL6cMRmJFWYrwiNUDZsnVFL
bmQx0IHFcTVma1+57Y9g28ZhU/g2Ku90kw40CoJWZCYj4wD9p0PsVahMrmSTtpVd/1JbjMrhHyTo
iNk25VSh7+ZkH/h4kD5lyYYtsRmSpmJEi4bkJP+yvlW9YIEeO3kVCeb6E016Q6qKy5qp/HBxP8JU
F9AHiFCUfA6xW0zRA6CfieBOAIEuF241gAfIA5XX/BrmCGtAJ6W0LkZzOCOoMylgfikDRLiHsN+B
14QCJ17hiRd89YWp+LMHc4+Jwg7FDe88SBWtQgCJEI8KpmaQIMqaq0ugUqaDjsVRH0GdyGf7R2Zr
XtvVbIgTVOUZnSx0s85aJ/LrA/e5JIl3IRdntP50lehbLGnxnQ406OWC8WavvJojOkmeR3xY98Sd
HNkrJOXICOAHuu/xi9DGuQIWmXDtcrwlgjSXUKTACTAYwFSY4H2QBzCCZuorxaGQpdoPpSEji8Uv
ufsJnNHy3mkraI6k0EuA4Ev7lhBeDlsLaxb0EdNAUb4oQgD47/BmO8jKFjme1bE71PkSFhRrwmW5
SLi7Ta39wZrXFbTT3jqC/RhXuEY0Xt9HqCQ5hcH9gjOq8HbY9bLtBnG9m1Z5OzUUYSNnmI9qJvT9
X/UCD3z0+KmoH1TUHmX40YJbWc5vTLHWKPOXevohzOiPL6zPAPo9KpvnTSC9GZATO2YmOkenb/Mu
f3QisnFrgWOVGJ9KiDMn53F6gtn5Uk1VQAsAK4Nlz4V4AUw6koLfMIBf3y+pJXAy1cq0JjjsiRt7
1VFUYGmqkNjVxaJpw8P6zGrwGr68dUaC27MbU0hLk684Uo6LHg/HXpMq63K6BvReRPfDvceUcXDs
HJyb2irlk/OUEPXz8xmlOIyDm3uJ8axJ0cmjO6fMVtT6zVX2gk/XwUqpAiLR+UB4sPAcNdpLkJQ1
QtqxEDMgnUjwPG4lwLTWddDXL5UL1XNMGzj9ZW7cvRoVrpuqWcezRo4WvHA51Yp4C2p25o9Xlf8K
DUI19onAjNL+g/cHuIzDq3up7mHQAfsIIkrDjH7dWFkdmJ3q3Wx3EdKeU3D1voGqKIip+nj6dUQi
fikOFaWZlZAaj8nclG8XkGF0/pyxNxuiZFXaOLcdU5IHMqWK0Xh3VLwsjNq+e9SpIztXCn4r4UL4
x1wCOVnayC4JDuVvQVBnGzMlAmvhi0c8dhd4Ka6rjq48ahWtYZB5FdxjumrkiZIUT9ftZdEi+bLI
zTz3YuQ932NhfR+wbpT7cbZWIhHbk03HWXLRSzHYLCIb2NrozFTn2P4MgEQZz4ShZu/P/xcVhv8U
2BY8Te5G3KC/wGbKSMm7qaE6HuZX+B4nplp1/cpdVpOATzctjxe3LfP/tNciLI+s6UZVdIuj4/49
V760hF2BOBsoxytz3O6xA5Mp4hIqJjeB5VUrlfsk1zZF4nAc6jrpfI4zrBlaj/tzHR+bL+SllzJb
/l5sF5nexb1Z1Q3+i+/8/g28hbSG/Tk7ai38G0FGgb3V3E6VOgsw0fhbEGrZN5Tu4vpnXutbqyt1
E/nJOsaf1W50Z3Ib5aFKKUcjDmzu2faasTk+PEsLX7hXtCgyfnYx1pMUilZbLPiSqxzHSDS80Kss
iEt0HBldt5K8yrjZTw0psq8xcYDsKXRQb8jkWzKddwZyvQ4yWbiI6SySoRhCKtgYHZ7JzcAjJ4Vt
JIbRZrKWk4YjPEbwfUH8kkAdt3+tS9hiGFz1fQ6dg+76SY4VFprTdUh8O+XFLSlWlcBsEElzIG7m
NgmeMRMk6+wXDOiV+Lq62ROz1FnjUMXXAoU+h1EFtcU7yNJjSFKheONObTV/Q9/INPffHQZAffnI
UxrDMuIMiWc4gcdleZNlfFphYtn5faOn583MPzraKqiTrRnrHnBmaeSfOfcu5bG54uyYDxeYqgW7
IBa/4mAoYtYUcOMmSGlyVfOmh7hMokh5rEHeln7/FYP1UhHefImK1JNXdg0M5eAkE094ViBWIz7K
6fzWv6ElcDuzRHlJzoseu4CJEfJSQnZsJ7YoAajYJbKAgiyBii0R58JyGhuJAweNe3UW8jOM3Lu/
VPbI+f/ahfFNoEvDNOh8xeofmUww5pt1wAsbQ7FdPoj5azY56YW/L1woDQeJhAcFNiUC64n1oq4E
acJVoq7njAZFXzSP/r/gUzdolPmhLPpmwpw1mM0T+jn/Oblq23Yt4VzXycNBGFkB3BqEMv07B+Jd
s+o3ZSQi7ck+yBMjJtcIqZeF4vODMDp5RqZ0h3ddCqzVxJ5HSAmYvO1mEOTEdQs0jaYhsjIrITlY
WaQbfokNICWLVOMlHcLw2EA5PlVxZSuGY+XHggXn7qzSPrW342FN7uLx/jjeRtIzYJ77x02ZizWD
LX858YJBqKH5YtVIFkXOAICre4xnLX3CbfNc57+/9BsiKwh4RTtS0ydX1URcx8zDf++4TF2YEJnC
Urbkg1ssIrfNuJy97UjyiSO2dAJ9Zxvz0jPOlT6eHS0VJwgznYezkPXWK9D0j54yyTA0upgP97l/
kv73h/uOo69SL3oZYWiyogxjVbciuDbMR67tPG4oS+YhCNV927+E73iiJpawSPZdrfC/OmFxGb95
8rYiQ8+QNA/yLFh+9FouWpbiD/1/JdWL2PAt+k/H2C4j/Y2SyFNBhWYR5r3urKTbGuQ1JnHkO2sI
l3zJ1Ef41C7bV+3uWH58Zzbl6cLJKBmszXVVX0caT9pWg5eBd/jWHSZppRAPN8zRvTyRGqvaLKq5
6DKXHGoHQa5T2KlHj+jO0yO/Y1futkthQKchwtDn4qjfefrqAQ5kraQ3ErV4fpV48XaQr1m5bMGZ
pL9o0eWY3I/yWycIcdflgHYmLpljetuUBdZivdOr+sktnRj9MKwI5eTYEH2h9C5zWa1ESbuv+jGu
E6eDWYdNBxMWfh4fbkabvMSCweHbkhbyVqHBHZ1TaeYPBcI4paUedvCXTR391/5wM1mgOS+EBqd6
BB/J8IrJmnLMQuufOmBvX7BeOEDQRHW8+OwleHxEErEdSSmxSYhP0iX+2aYOo2bqD2bIW0oPIxY5
ReuU3mlh9VV5Wnw4CVIPMJFAfu4SE1Dx+jMR0NUyCd1Ch7qkjHTaUlgIlh1/tTqMr+54ZMr0AU3+
cTf+LYBdkqacYLsNUqidBrYD2SH/0cJWfH309J9NGlVKECPjk9slw2zc1uCWB4P2zCIQVQ1+EzjV
xXkul8iG2xBwE8AVqJx+RDhbBgpPCXGp7guIwuRRyCuE2AEo6X07wxhURkO2RAXsjCAAdf5HW98i
b0RZkGJ3JBSIW01+HTuS1/eWLc026BNK1+zbehyQHjuNMmjWOxGD56FhcRO6rG9Yeo/4+KVhY5k2
JchiwtCOsLI0XKp5ySNwL8X51yR42Uw8F7rU/q0PsMHkvYuyyB9xtj16IaDFfF0AnRoAyVnXVkHx
F06e7Xyt+MXza1ARFDx8stBFk13K45LyG8g6Iv3QNCXhG7afBlZveymO58s/KCexV0wRTMHc/iM9
FwpRKv6BpOoeynvZY7AASJjJD36az602dcYONOo/uFNoJ4WnDroAhK8S4dJpraw4WmDX6iuLqnNb
UY3pGW0q/VXgUsI2zVw5VKdJDSobjDLsX61z7aXOkbbYq9tM4fNM9plKw6+q04J2QghYkTD9QO9h
gLiYzcEUVKySpX9Jj9I5UZ4AN3oiA5bwuKPjZ7/+us2D2wvaJC6w+eWvukySaWd2x94p0FcFxXyg
tR2ESY2IZ0RtsYgtiD7b/eWMjFqeEjyoy1GpIgdTukAWItkYQZBj1DustS1xQfdqhie6w1IdZi7k
m5hzAdqx0T+aIRldWcfNLT+0HZ1Ln7fcGmnAJ6BI7HOPZlzFGFvEpsV70fauKFFHJcm7P2KLmMcw
qQhwp7NpQYz2TYWRBETz+FNRIYdanFds40PCG1xczW891RP2qvYWAdpM4hnUbYtUVNb9kNSEzeKL
m2vlOaU9SvNfd1iNbiVC0nl9BrkpICUepi4hGW9TNbgyKZq/KgoilGrZbTQhrwbOnsMUg5t3FqrB
MZaQSWTOZ2F7Ia/ZAweBQOGS7id7L4BSKCNKl02nSSEPI2XSC3z4VBx5Tbs9IDeYtFLkYANiK6RY
+pdFHO3k60+DhRD7mr3CB0BCoUdmoY6wpMYrRITN7ILiJFAVUZ4QEQNcbk5QKQ7R/liBLn+J9GAh
bjjeUKnHj5vgskeuUWLJhCgeqg9qnr04CoN7JJwiWQAssaEjNm3DXHFWQcULmX5FcPRbhX3uUoyj
t93iKCz8S0g9JJSQP08IbREg5x3kRJIjg4txfxV2ZkgKmACah2sNj0SZKyNeIfvDnU7jgtr0P7UA
NvAynjiFHSXAHgZlMQTY4yjxDVirxF6RubxYeHHt/gCqrYjdy+SW58KdmPsEOpZ3lXM3J3i4ZWLu
30Qowvza57zoq0CzMAZbY/MLYfFcFTtuOiWRJwqmQ7C2L8z0HddmMjyl5vxlVHy4pwG7tJX6YrFv
+kvQXolhLbd1hicRRwK8TSTkewaLIRC62MQF0j+AoNO05IkfQf282QHQ1PavU3cSh1Twdg7TZC4w
SVUBhggcP7GRqqS3gtDvlI+Bs7tb+9VtSojm7mAX3gwn8ZxtDFCa0HJ2nI1WetvLHOPiQvW1oEwO
4lTVI/4+nIeiSDczRBraYTB4OBC6PxY3KeAy3/LkLhOcUvC/uE7nbbCiqaFXzc2fEh/+4nwhFbgj
Q0a37v1AsfNxelh4M9+MJVHmUsTdUKvMIohb2WIMvb10LEW44sVEEojA/t/ui5EPRkJIg7E7FsK+
VeSI7dhv/js5Z4f7yfEQ+39faGAFZbZ/nNSzLS5koQrhlHk0v10DV+YLxf6fZ/1X1JAWZICZHzAW
An2mbLFltoYpt4c5BIHm9beqOiaiR3oLWP7yAdehpu24gOWmlN3MwE1QE+iAzNYUFOt++jbkeD0B
TcELvcOzrwZmtMZt4SN+WAv7YOIacKjmBWROOKrPYf3nOXYTCd7VkQhLHVoibixqKxPTP3YekATL
AfAqi46ROukZg5BNgLi3gBAZE0671gJWw7vcHD6Y5Ym0Lxxo0E4WGt1pJ+QWxLz+Fh8aWrHFCYuW
e4EbBVEz660RBr430zMQBMkwUWsjIVnEeXKSc5yufoiMi7Tv+dlMLHIxD3xggbdQeyFFV+xkkMW1
658nfXsGqN6etz+Y+HBj9AAnbNAiG2XAOlAQQ4MmEXT1ynCW+6ROWbtdMjph+RyXaaG0LSo+LuQy
sxe/nCp5pkn+EOVncH+muVbPqQ4pc6aCS5L8PLVFWrVXnV/8UJ0G3I46LqLtBRwiJgCeWxBwFc2t
vXRXgdwv34qVMTom7yKFIcJ9SvW1wKsFESjIKbT7il6WMiZk5bxsRCQSxJQh7GgX5+flaA/djk6O
7gcVZ7ixxh4nqHyeyzEb9VSorfeCMgQyFO7HFFopW677jnH2CjQQNrPp3szXqRUBv63+aj5nNX57
MznOLU56bxMk+VxaXPKiOvUEUnjecHbbTTqUs0jnHoDtXjCZfKF8z+a1KgRem7RyMTgAZUGo/Xsj
8tNFpqXfLxaYZmYHWSSMfheUf5A8WrJIT3G6WZjp8PPgu4BjcQ0pBHeCBqt2PzvHGB/1IzSiOyVm
TeAKihcgyOZ6sQ2WJqZyNsfQ+f1mzkUT+3DpPhTzH47EBjxI6PDETgG9G4Eu4eyX8o6Os8/LJtzX
L3Ud/9cqYcW7AJqGjhTmQI5DVprjSIVcqbixfYTXVWMekTXdAvUK93Ky+XlolVMdLxAUXnpt0B4W
YNK/Qerk6hIfIOtknlC2HsJFNq7eSeoIwndfGBOfLFruQaOlRXLjDqgYOefsVI3wJ/zNdw27AnPy
LWBOQXpOygmdX9Z4oSu+HGHLs/jX9tkiJJUjO3bO9U0zyF3BVmivhk2hpkc2rN6z4ViEfii7SpdS
9ZMzeRMb9MXCwuIHFo2CylDvQGgWt68fwoftoEzzOFaSL/Lip7ssRcZcKNTSQ2jQ9X6kfOU8SB9y
krqq0JV6C132WkWn8Hy33ClIRDpVhK3PTr8OfwksU4eEfTsJkFvKq475cLPj/MruKXe70qESpHI3
hgvi1/0QqDeTFdAwVNEbCiIfHvcpCDrk62nXy6PSrxtgZwQ4fhZ0HLgf3ZJC8gma8AtSei3FA1Ka
t4HpskFsYcPxIrtrs47wU11j7KxqzjB4Ks0o8fmYZ6c7sJ0fPu0YtHykWBq70F8EUJmptolhOCaE
cVhHq21uRXWQCthPJHsZkHa3TW4/4+cqcPtAum1dgpYTSULTBij0bg2T0tA0u0xcNzI3fpr+l30k
j+PSmaRQbAuNNpZY131woQm1N25GOc3ZPLL0g7ESAdI1+cDWwj9Td9qgOKio8oYGN5M7c/xbXHcp
X1fFv5NF0uiA5q6wfrV1htlwLJQfpD7WE2HNP6do9Q2KWJxFD/mLGJfutM3nT5vH1wgVZ3OWsIl4
Ex2Ki+hD8TJu9uy0Oy7YQ5iGtcad926F0JP7VEbdGNOGKKPcn0BH4+G9IV2IDlo4lE8j0qHzE3Nn
PcVXntNTkbVrrueTAlcmxWTmoRys7rjCvm91vNKYFJXRCRxCqeMEvcpWqdyGHYhxIayTYwgdpsP+
8tc5ZCesFTCLH/tl2KSmJiB75/rzWJmmDS8fXFf591ViGlzfuNFltZUqooUTCUnR7mrnc+sfr3/9
V1MxxAcU5VJoLIIIDu8zsXFVhA/Uz2EMYG4ggDhdQKZnR8IWeo90EwsyXRmWMLXKla23WCo8cTVs
IML7mnYeLPR7v550agjAoJe2U68AcE/gz9Vt19LsfKFwlERRKOaGed+K/wLuVbDVlLGgNHx/Y3BS
5xMrUnH8UoKmjXLjy4ZQCM0etqyWgIcPrUVAfkPNRDvDQFyxlcF4iwrauPJaoYEIMduzaoaJsykX
xwy2R8Z63jW4WM6JWvZZpZNiE+RQpV1IXjNGSfwO8VoNxNuG3w5A85fE3GsIRxMVgSJZ3W2x6ye7
J3ZZeqbLVyXFGZ5VoHK3SAozD4s7zqGz6xpwXkbRKRQ0eKLOspPk0zU2tfmFlxDfnhAEHt1p9kfD
GrfQAXevEEuV5pGEQ19svkw13TTJczowV7HWOXqRsf9XSmL3QYVi3zvYN3H1sFLmGvOVFWsA305X
LNSaDWsMIsDPsAYnwyxyF7VybOAzU8hv5f/MxhF4Rl/mg7kvLYJ6tF2t3S6MNQR7pEpzE1+/lGWW
P4eCVSfdtaPj3a3c/JCUA6cjZc4Kif6hdQtXX9Q9z7/8hR8SN5iAyATi8V3+UZoGW6f+vgv9d5U0
/08XR/LCy5091AjCzNLawRhlj1VO6Gk1KX1vVyFya90byaIhYwdEUftvAhLBRrEaxf9Jr5ZplQaH
ZIJz/K/TRH9l7g1y7AyFuaFzFjSB74jmnzZONoHRJ8EkDPdiIKwf1rF9a6DsfgdY+nzWZiQ1vSzI
MHdTZ4l5Eh8e4AVrPG1z5QDAtrQOL0foZiZiV1vxwUYhBZy99l9x+SMzmZa9780ZSfDP3eUcHIUN
fIn+lNh+RfPolAy0T4IsHwOALoskVdCEY1FLW5yxuFJmUq1HdTQ+y3joCplCVz0SCY8gNTFZ1aUe
G/iaM56cgPqOyD9+bCV9Q8UdZwI3pn2Y1HNLIdCj0TEsLI2rByCE8BcObVbVKWBPAnBQdlNHkgHr
PcftYKkX5U1fLuoRb9OoOFpkk+iNk8rVtXYDLHJrET9xBjVODQeVQExGzCf7R5B94M1Sjn4n/fMM
1AEOk0aypRziI1zq0LEPY8HnRvBzybItv4mgoI7MhIDC8Z915ev1OJ1UxXfSAAsRnqOEGwkZ16rH
zKS8qgqTnKgsuPh8d7TMbl/1W/sbzVk8cjNMpCfR7YvnOU6cOoFKp961mUqj1PhzdKhOhyKzmt0z
5ZCbVTeF/e/keWQpRsAgd6HvGg5LI3wPBBLI407syYdfvFgEoxRZ/Af+WzDwA87lPGkkI7ONcJw5
AITMgtmYJPdTr/m++8wfH7u1eAVrEHBsVFAS9DmZFQk+/knSF1rvLApPFQxgqiN4Ggdztxk4F86p
Y0I+N6euyl9yXFw/NOfQFBE2ooyrjIiFnOuHpBR4hH0BdJrffa8a+MY0iFS33XaSroIn1TTviI9N
F0uOM2bvRnwPBvSZSG85j9nBwXiDiui71GFDgALH6YHaRiIIiReMaOZ/rX8+WelPtbPPmDaxJ/Ky
jG6faahptN0H06oAMc5CwAGfiM+mVp1LMJhVnxO34R8szJ/K2rlrYcq0N7vhQpzNG5jb7zbCN7JI
81ZGX/fVC9FPyM5pWCYRdkXPgejbjsQRQN9mnkQxHDO8hjBsCzbqPKIODKTv9l/hqS2nRR8sf3fk
KrSEBhhDhF3ciNKDVw0fF5UKwsluvm5ysKfHzECAeMR3r0u71YnQiW5hrVaHyNRpUbOWkia3r+c5
KuWEarLwvzTtp6/BGslPkUicjbw2Enp76YTRl/vPtaJftqRkRG1owSvvyYb6areRKbpPc2V1VlXM
X8uMLBf5mylBuQJCAM7cNZPjwIRyRDm9b6ew/NGJTA16ofMWKy9eXPhc78ZnfYNqWoIJPpd1Ok6T
lgcxtgOoSoprlm7lSn2XGE/LSguVYDPMXUZpr10GrVIidFF8M629qr1gfznEPSwP5Ws2BA3uWwjp
ii/59fu0Aw6g0rPpenj3RC4LJZa+WJ2ekoO5Zu5Lta+cKUZlUanJ6960vr2G8i5e+96TuPV2pdYO
rYZEhYBGKX+N0HosttOebSmdg2TxsYfLcSYIhbVztC55tKvpfm9qgMHEEA338qfswnq3Z+rusmpE
JloDQdUENdSIi0g4i4Z6Hw1Lgd/1BUKYC+wD8PlKZboTBZGlhacEAo68qucVQL2gSUkFAw5SJ5XF
bnjhHdFrJSDrHXCL0zMDPZvBsjhX1uwriYJ9AbY7HlfwuEZ4OjV+Ptj5bh0VNNfi7iBgg6tvGFel
NI/Fq9XHFFSApWIumuopUkaM58br8M5QcNolazUGvSWnOLweZOAciYKsvbu2svYOd979X5LuNgMa
d2gmuepoXRqZi1rxWvE2MImnxNdmYXPCFtDoIFn6XJrKVBVv6zjXNcEYsvYG+sbK/al04YqNMvZU
xwpu5OrRu0UnWpctR+8bwcChhJTo/ms8AYEz9y4LkUqIFLkYp4s3x3qOj491xiuW/zHothU0QnNY
jp0TVzouF9Ve6714FIyp73ekPdugyybc67f+9Y2svHfSAjMSpuXy9TjAjOsptlEkhwjedAEU3VhK
mCItK8HDXVjRKHNezSra+acsJfEnvSq3hHniU+XlIoDM1Z+PaTx4lpO3YC5994UJId69YCzxHcHl
wZQmSFJMJJrWBJQ99NJq1wuC99xDq5a6xF9fTG4EXFi2rvvWzFk746/Wra4+GTa0uslnbRJmPO/V
DvnhXc6Dwopl9h8I5jgwfgQPN4/NSu6OENBx6pVNfPkBPVT+UH1Zl3mypCoS/NPgpQySbjiPZsxt
r2MMzrJtnxxss/26IQhqLyZ8LER91092FQMAsGXa2Ky09SyekVshY2xDu+2QNZYZt5w/m7Du+6y1
228Ojrvj19C9wyTqfaqNibvnRXin2lQQuRjANewP7o+GvmOgvO+4mHOgrbwCq761qy97cu11CAJW
VlHI5pwFPICWhnapXhWOSjXAEydC5BszX6let2mzrpv8uO/Skqln/cWLEWETO/UOXIOWd7azavUu
ZUu3Yb/n+bym03mbF0EOHxATrOr2Kgo7Nh7MGi/ge3DKY8ME3vk3hRNdKP0/iUejKh7okYLl3EZg
b7dhQxzjjb/CLrlhyyXjBkb79A3IhodEWqpKdRpMuo7fVxo9z2kjHocPiyWeKAd90qRPFGBTvtga
uUsmWEAcOLa7AGnsrfGTH/7tIYYogFruglPpgFMkOd1hzUVy+1h8SGs13avSnwDCw0cgZ+nfNeIP
OVAB8i/QK9YJwDDNghWJwnGlqn6xhSEGhyQDxyvNy8ByUrgAgERuaIKg8K9g8maUa9Pc7H2/i436
qDwQCpydPwcZMLqS0kr7AkaV42OT12UyZKY2L15D0+OSY53/AebydCExIalYhjhIJZqM4hmXxMw2
0b2GUREUkwsw+uvzT+k5PESfRP3S4yq68pUxtNVAj/2MdjrZivLlpEbT7IyoxubdcNJafGOh+9zX
OPVfxMYY1Jo0C1iKrVcmCdDhnODJDJNcjH6lK/+e+MFilaAuG2OSrn3yQfvDXSdtv6OpzfN/bvxa
XaaBinR5kqNkRvUj+xLWrM51EvtOFsJJrTv7t2EDJuanJmZOagJxDx4Q7/VvAJKhqBXt63omDu7D
s9RIwOoczutSHATHXiRVJ5DxjwDZGnmech0xmdSwrWBXyvEtQcBgu5YvyGjsC6/zYovp2ARyhzVB
teTk5oliXVwG0TDnUMzw8UYm7MbmUGWw8MNx8/b+LeyjCMSKjNO/H9EJsZC/cBVdBL61+txWu5vY
Q5JVdAA32dq6oUbfZRRGZI1+YT7MMS+3kIcgDOiolstlycqCixHcwSVNDrpfzutaMvMb3MMUxU2d
5vg7Vm4Ih5Jm5VGNnllVsy4f6nFzdXOPYbUDKtjlGQRliBYT1uyzfyB5xQrwK7UMaOOwAUrXZjFy
PGPKdCgM5C/rXMQIx5fXVB/jtXSFXrHYhoeWGqD6/ZUC9MtQDrZxmmdsMEaTsraeN4QsxyjON87K
EepX1kLvWpkFi/cMeq5Hubj6RgEsQXn+pWH6OzxKUFnwm+yv4d4X/zIdvLIbJ3RQnfHZwVORj6kN
sUYQnIXsrPZFbCtE4kf+2np61rFAURo2oUIPDj/Ndqu49/t5IqLykOh1efGFoXvZxDAJc7sC3AuZ
Ql+fLJYmWIVt7rZ5YhW4IJ+LMjjcd7RWJvUTJW8XkAh5NIkSoFI6eZ0d19NHGLZQn3jdLUbOmn2j
T+uGNDJeKqznGwXyV2WFNtiiAznrDcUPyXzfTj8Odeu8l7S+4ptZ4TEFPya0UnarX/gVhXLeNHAy
aE8tRl2T2sSaXz4S1FxtO/9Nrwr8BaDsfd+0Ox4QSaIiuHsQf7xSFiM0OTtGMOkL6H7rMhKI1vR2
eC2KIvR+eyalvtOTrCc5qgPDkszMCOyL7LhGsVr6sTGFiVV0KMWQRwtBjxuBooCPZ20KLfbCReWi
5GhOZ0IO9NQBpBOVS3IXXiWc4Ooh2Pi5QjrImsm5L1kyYb0LJFjb+bojRnYA5o1PrxpGVZjLQ4LH
JnjBaDT4wCcRvtpZEiyCwCUNCvj0k1FwSBGY3gBit0eR7DaVbZlhO0Qw9ETLVTlRSVDehWdRAXeq
fwAUFekqIEnkBCfJfd5HjwFEUH0BbpuDk1POu7RNRbnnABE+nyIw13bRSAyYV0XBS7PzjQJhC64h
RbPGryX6QhFVpplVwqf2o0yKIWSCYgQi2kMGx0rXaLqPZ5ljtwyjXRJsDGu6kOC0ORLITG0uww5p
LdYrnJ1YMud0g+1bIWGSUOMUGXLDancmrGJQ8nS6cSZ4EnUeHqXb+WxSjX7E5VOxtYkmyEsycCoM
W2MZ6bVofVF6vTtp3jsRElh3QFK83x5dcGTI1EccQ+NMtTF74FQ+iVncrJYo1GtB2spmKlEYSUFR
kiNgpgSBnPn0Mpdx+XF481pmpWPc2t1/MH6tIRHEzBNkMvMXc7xdoCdjJ1R3KZ8PXq+JEcZqrLVd
j0m1K1uDI3lb5/KX3sH197qN7KM8CupYHe9B5R8TS3aLZkfkuWV5kDmHB9SQurLpTE+WQAutVqQG
EYGG5JPuS9/7kQTYe5kFK6IkrE5xMIm/KEOj/kY4TABu3jhYEAiT/+MOsNroTAo/puAFQlkXC/WB
Q4wAKVGKVcb/P8IyrUpWsx135bgkmxD2NWqx51BLfAAAeMnMxKOaRi6+7ubAq8CXaZB/UiTtTBi3
iG79CqteE0GgpuBZRQ3sE5fzmo1g92TcKhwsHa3Agr0Q8gYp7aHIZfFDC5Xk5LCWReUL9H0eZ+y1
J8T4xuOhc8HHnwWO1Ptj+gcrdi3PYv8LSjYKHeNck4KstWCkTnrts3iYvRq/K7qsk04Vt38BNgn5
wZX7V6961PacbA00eaQAS1KQp/8CVzWxtl9DH6MrM0sBORreAk5HDw1lTTfLJ5v+wrRUDzg733HD
pLFDKGjh2Nq2IKnigqzfa9y+MI6RknRcm8tSIIcwaPdTpbXLlKIG1Wib1w9EZhAah6JA4Z+V1vOY
WVs7P/U8sG2pHpmwEx4iIh7NzBB5G+HcdG0Z82vuSdkgUBZZtKWysG3P/hKZ5pixJq3TBqa19KYn
4J4Oz3vH8K54BIftmfFmUUjtc/1DF4ep8ezVzZFwRshcyZYFmwjhubhL5l2fsEDlQXM29NKjWecm
XaeUTLPOwaY6zceEAgckpvsICEHgmGXBZTyhbvPjCfuSn3VjwRvgJsx+BJD7m+JqVJI66VCEgD/O
+jZhoizvj/Or+x99GmXEWxg3/ZwdNWj6U8eiaYWoczcXDKdx8g8MpV+HzvesYWN4eiRbKM7RjJ6T
4YpbRQuL13apl0YgnHSJvYlY4C7nWoSZaRTKmlrjnMesyhVx/fMlnrs5SOaqHoFZXKmRMBkFl7/7
NsvnM6OviacKMw0bBc8FWax7BwpNoXk/elx332FUiAjzGsbGfLgT8s2ACA64rnk39aF/RQsFpRC4
H/3qeUosHzXxlC89QFbQXvux2rYqU/qceE2KP+92tBgC/2cSHZq4r7Wi8HVQjOIGoqTiclrmmYwd
5RTcorEHSCJ3f/yWGeeYxXlMZwtfVanSaMUOwVkO9iZ2LKzg20mEXJARh5C3SfM0C/xEw6qNqo0E
HAAejMGGja/xVcBzX93PKzvEp6pYJJ7cdEK9ttVuC4IINmMrV3bK297f3uQglVaB1Lw/raOMrC7X
Nlgco+/IJDaCUs8RrigZE16QE2ot/aUuyFBI3rV/C35wvf/bqGuUE6ULka+IHTOhQQQ7gdiEIIAz
Tc+n8VLs7GmVVUjrMzKQ0ncWKtV5T36jhFHuoGY5C8buZ/3epJ2bgg8Y8akbr6KgcBRdr1kBR9FQ
pe9H3LhngLdt+hlrvisRDtDyhajDGIN9l3hAhCVsH4TBdquQL99aT4/0rEcQk6kj4k+LC+XKTqCH
CYdM7ixNaFWxv4uS77lhEkqtLABLJti6cP7af3KWiQBUzvIUmhnaIs0Vv2I8zzzU01Bg6bGVYWG2
dBpewCGgOPvu+Rb9bVpvd7oSfd/DDhML3/LFDQJm9l+ukoSppMnd1x8VAaRmGf3tAMK8J9L1Vt6X
gg0iekQQS6PTzxKqgbsPfVmcCV6QFW5AtLDzUQo4xIYYhxRUOvORXHHsdz2/SPFGlB5YsfOb6W95
5PNTvXn7YUij0+bpkryL/srbXeT8ig8IS7UYA4i/y2kCUyMu8yWdvcEyFYvkjzM8laZPw41vJBZX
OefxNHDRgYj8gsiN0LkcDhS6daA89+14mdKm5+8QI0n+xk7WbM9a0vOI6WorgpNOxoP7YTmrndIR
BBGqNwYf6VZYTnHgexWdxM3SJ0jhW38gQECX6OgBsYLEAPzOerwhEcx2QkuOuMvgbWVYLRp6qwa7
Ys5jBtCypGONF+PI945hbPFAD2FbDc1uxYqN5XbLz8T0CMERAyXiE9UU2khclTI+jL8GcbnyYa6G
eS+PxiuF3FLTiMGhQNovM7rC+BG+eRXa3J+M0tu7AH7B3SNW++VdzyBt50DxvAkaTjuMLJ6ArZZS
6ROlaaQezE6lUXiRY14H548HaemQfY+S4ZGbln5sv/Atzs+uOeHFMyZhOod5SaTc3ITSFsTWgixI
6sq6V63zQ0ux/pYWKuABcvfCCRpmc5FVhUyT0H7HhpRAI0cRYBzntSRnucXCWNTw0X/uEh+j5nQa
yK1ezH7Y8jiZ79/F3WBRBzuNQYyernpVF66kHyBHUXwdVlZ4RwRo6IkuJqHY6q9rSg3grFTN10Hp
QZ3K8KgUP+GaTUie8nV3NEq2CFWdpY7vhSTElOqhyK+YxkxJKGknVurJGZkO6l5QOUTFmzJkoD/y
22+fZlac0sFYbvh/Qs9Ca4htU+a1TgMtqB26YpVo2A9RaTI6V/tbz1Go/ZX1fDkrm9xmSkvftMPJ
NzGQjG2ycHf3XMs8XH50jK5t+69dJs73ZP5QJXhPjG9G2b4vQoOsJxnWiHHK66lcD8PJ0endVf2G
vZHBJpgvdoGif5QVIs2JzjS5yG5WkqGlG8UoZh7rw2khq/zDkbF4N129qbVEUUfPFup4NTJuquuY
ENkpHPVV+0nAQMQy61CvIYsI8KHKHQlLMAIVaF3SuJBOigcUQs5nBZL4d5HCE0dxvMf0SKtslkbB
5O0S9gE17SUXZSyBexYHx/U0/dS2agUN+Ar+Y/F7qW6yDR5UM1eENrYHdwdWQycOjPzm2f7gyzAC
2LWaRCcA3KVHaUWGCInoxVDfoQ1NFGo0QN1jTGNMxnk9fKdfDpWNIDDbNHkWhobQRmcJ/tO6sB8O
HItzqcCh2uFjAKVjmo/EJRCOay/dwWxzWQaOV2nLmuNvvjZJoxrRW/j654rlD7XG9Dle1isPTCD5
0TRYnB6LcKZA2ZRB80UXuDLp+9xBNiD71dCggoJ1ics9CDY+2rNTNdMkaDYiDAmeBJYDhs8hBBP3
bPPke2ayVwmIrQ8sSgyxkoIwNniGuQN6Th0dyfw9NFL9pnbCnyEAykLyLjtTub+mlN8EKNxitjcV
LCh43JN3B669EWIIUBkQGy5AATZ+7uSmkmDqjv0Ye5+AHou64qFnTzmXXOm07QaHHy7+uv9CABBr
D6++xXLO75TUi16YaPKLy8XPTE0Gd7oudCW4X4MrShWdRTebFtPs0l9Pv+5HA3aU49uqVwVYERp7
yHdNbRUSizChWg3wSDOJjNfvZJSOqwyqsP8utDm5Pez1oFiXpXGnu1kP7ul1dviKVDcWootJUsYo
FsCqhgOsEJFhVFvPRjeEiCtACLOrtWov3zGgpKk2B+byxJfbeLik5g/F1D/KRHy0PvYuan16PaCD
OHGcBlPRN9MDOfoZpEwN3tdfadofjGdHgVRlBoi4QyBhAG/5eTk9axP6MOfvKMrQGZ9jjM4My3+4
ZdRNa5/b84LwZ/07qSfx9fnfmJ3FhiLt5tlRiuTZZlpZhg6R9qYB02iWylK1ZhtOKwzmJR4jViiY
89AncaPZOEiOl+Viy3UzuuMdEu5qFaN5Cmcu5urc8nMIHf2uab4gZsIU2B0Po6Fg+C9b619Lf7CW
dR2yrs7I2ymecymkklODtFvQbWhiUpRb/VYewRmiNzrJxYHP0nBwyJ+63t15e/TL10tJu8lYnFWT
AOz4avugo+CseaprxZpZIv/kJAOhucW0Go6WuGeZOX8rGLa+E9R/Kf32HceQkqbBZ4WeUmBrbpMc
Z7n8pEKpgTsBlH4q12+KwCwb/3EsW9lkuk0ilmZXG1IheYPALDSROGG6JEK+uOjY/BxJAoHy0F5h
jAI2uxCBYBGB/qCBNNE9v1XfN5uIEAkHEd78MFgsg7eTfyPOZNmLR0dQC1dIjSY7ari5yh2CbHmF
Z+ELnbVJ0rlx6pDCql6MEcRfQErAaTKPcsrmGeLRvTLXKj/7tTJta/7rR8fpfOGkZnhoBsKBjlGP
ftQe1FXuRfcCVRj/GDE0aK19msiKaEonTdkqobe+L182GddjXOglKP/cRQQkj8M8muMxmj5Tt7td
vY0rmvaRSSNQRGCfBl9mVeEXhuWFSY/sCzxqknBKeNoHMYkKmDVjT1XFinK1MbIPq2ILPi3tmKOM
0Ois0qEaATyv8QKu/m+tYtbKWMMQ622IzWhFAM7ugPu0Y3nnZr8EhrL3CfUws6LV2MbD4nD8hNUX
bZTTBO+jZ3dQnltorVuG988lmsmy/NgXhkEgkkt+mspy1IP9krgBWblSr2IQj9VERmKjwsC4/GDU
INR5wfAqniEHYn1uUOxPWhx+Qu4/IwT7rwEhzepHaAkKHIezRDpNPxHEPYKsYyWyfBDTLN5zm3kR
Yek+KEYUqGysCn10Gy0Ovc1WZrwyFBzl9r7iOa2l3y6wOLJYZJKkjdkqCGc2hxljjDBUp40Aqjdc
FO07jaAerhpu689Ges8S3nhCDAswLlW+yh+s/4KiCdvURn8euiH6q6fCEsFAOwjnaZ+MfMyQaeF7
OAYrIm40G/VlQoQDVbRXfqo5cKkyqYKNgvm7505ZoKLO7pAC4roQLbkQI1mkFwxidMuZ13PnFNep
QlTkqniMVdKdEPcWQE72aLAKJjIhmH3z8GPcUoU87cWN03iXIJkCHjsz+0Zlo0hp64VckhJSU5Yr
j0GE1a6rLy+99jj4q9YM31UyyNLBxwLja9xbSUjbwah/3feK9HySsrlaA0hexwHylUj36TBTVtTI
BXxh76+hzS14H33so+qfHfTlfQgUaWOJG7J2qhUwe5OdczH4kitJmrdSgal4ex6+ajYthFgdbmDo
r56NGyhy6gtfALIzufLWitAvIaerQYx58JzvnPx1VvkWVKYOIgKOrly3p14kEcGjTYJdIUk9q8vJ
wc7v7uOFxdc5Eo5qVD7wd20idOTSUyZFJs82KheAto78KLums/UxsTLcjeNFzt1okvwqJpe64V+C
J7t5/ZfCRlgB2d6zPFhEIbrpXpH02Hl9/ZJOtTNXesgbdm/J9h9Xo5dn/q2cIWqEffUpMqOMAYnU
Wtn0dpN4V9DiJRPUrnt0gBbF7ZjoUyZ002E1f43U5JNrQwwz7uQx96Wjwf+U5ZliziSR3IQHWp+B
jvSM/8IqEPm631xL5xGav8acnzX/NyDa/4S98mN11PuXSzAH5mtRTUPDFOfW4irjt7kZqB52t26w
pXcMk4eeQ5mflrGMc5pznCA5plQoxFmvzBv0J9A25xERbAzmKFCC8Cob21AObYivu5pktxHoPgOc
zIElkepp1YoyBmjJC+IY8jkSr6eSppa5NVNWHS6NIkAyCn0RuNIcYEovjZP+AvQ3yKZ7LwWHWcn0
8WwauprqD+WKKiQk4ytIqHFczAclvFO/HYXfvJ2Q3rZEe8l7g5k1H8LgK9tsPa7Dyj3PrTGU9shu
zGSxngjL4PNaT9Z2IIuKeGP4jj+ZiWa+1kckPJFkFq2f2Qnkb5yWNVIM6wkkESnkI8hX/Q/KLsvr
Gma4sHZTxFmaxS+LRA1bVBOH3iwZwUnpbSxqz9R5agsXe5AQ9lM7YjeKNly/0Ridr8LGpwBSoDLp
KbRXez1w0qo8lIDccb1EW94PLif2ObQT1iKd61WQHIFiuPwJuAQTGUbvMgfmQvTMDoKWjLWEFnGu
KNDuZjYSi5NQiJoXzXT1w8AiC4jew1QPHqB56wn6q1/BdeSlD8MwSAL04thtNYhXSAjjBrBLUVsn
3usxiAqRxdEu/Bsj1/aVZtKGiYqQDoz8+uJmKk8K55mVsX+nGr4kb7rZ6myp3cM1mjn3GR9fmBAg
haXKbIDVxdfYmKzLnsujNl1SZ2ko0v7jDHEbPg4G91CYj+T/1fdJqtGtcpygC8Hp+4z3tIg/1sqz
1YFvo2iKtNNlN75CcNV110rSBzKT7IjS7nJj8yqy/ne7TRuYu7N3vj815KsGsOYRQVC52D/B1GeO
aEPQcRAmBylTwa2lDtCLwPgtF692/P75AJNVAW4Aty35hj8qbYsFnnTQf1d1S88VLhdm5yHWfP5T
sgb2CIXPcn1+dy4XyPDyXmSCUi2BGm/Ap0u8lygO8JNnR1TMxXLwh87h3+aChxDiFudLqEP6LOSI
3hu+vFazIVKPtBX6AMr9alHgvDp0/xCIRcLZxQWF7vhE0U9sOxhAkR542Js1r2KOwbuQ2YERQtJD
yavC5xHHZYmPXtlOWjYkw2P4EdX/CbVwsEPFSKUPyC+OCV+MKDMn0Q7sCJHAu1LRndpzC7IE76+K
hx9t3DlxqHk0XzxCzYdPNb+a2SHW9f91SwMtCZgAqlCXTOPcUXVMY3HbB9g+l8cpuby/OcAFibT+
AMCXrw2XkrZkEgvSoAvgh3VeeWNWtzifnU2TWn5JAKoQIIcEkVe7xzTb2blwSyr8EcFJih7lYRam
YwRzJMJ3u01ZAfjv1TlkMJI8lCAZE7EmPxkapTt8+QjOvcqQGr8bcZhGxpmQ4XvC6ImABY/WxcQS
dMy7psXh857P1SDArQz16UgsNUJwNp4KBR6R3LC1xQigSC4L6nZ0z65C7QMOiKjGCuYIZsU82wBs
u3/eNvoA+U9FHzTkfKf8eqoteYxLF++RtyBFmR5tSMNR9fmbr1eJD7LUJ7lCBfHfiENrlnXIYumX
EyVnGul/9eytu3o5OTNHNYDwYw0NXRIFZriOigQI7M0FJqw02B4fPkeHDptN+9sAaOvMr4ABRYo9
ERw81TS5urBWQGpgeC7HZfVjRxIzmZNC9HMz4302khkGIK2nDlRDcXVc4hdR+5z1OdnY0gqzPTaI
eJTeOGrFZ5xXHh0yBc0foCRgNXnJF9eDm7aWinKDCwk6qR4j9bAbh4tnPEQ2b3xe4rozagM+jVVQ
o42hgHAuM9aiwYPs8WfO3GKmt7oyal7iui9KKjZHJ8KWw2unYcCQChdD80kMQpViEbaFpZklNbRV
QmW28UDyIJ0t7/YWoD3mqaUrhjCnR846j/Y2UXtayzGiPqptq5iSK8Qq4qIh7hubjT4mpEr3NG4v
iSHwRxpTSryfXURnQcl3m2syFPRBLRZAycVVdXNaFOxnjKjukYJbquAG5l+eTYDcP3UBzvBrTLOx
zJQkk6xL244r+EvgxygKgqnc730oLevT/DtJGj3rfRwucaJPm2JRz8iT0nWeIqhHCBotC+LIVu+M
zKLXuwRpWj49AE5j/2O2axzVHpEpTLamcvm6dK3euhdhoc0TPHpTlFRMFGw5vJfqeFjvNtVVzFaU
Bvi7I8tTKVLdEWy9BjCZdrIks8MpfX0IsVseYQuBM1W5yLpJkNuQ+x3LjKG4I/a3dHeIdo2AmMSm
+yqX75lkBkGeDerySULgoW4eGn/Adock9yqKD+ef/8VLrhaUFIvjWl8Z3OdhnwOzlfINOiN/oo8+
ciltqY27lL1lFuHRbVszAIMjKnkJmKrCEezLcx1rETQBZPp6TWquGfqb/yRR3xKY5K0Un8bt4ttn
SF2WGKrye/ysvYaY9CqulrLK3xNc91KCIi8AlfMVMAEg51JUr1a5mfh1sguSQRch4Kg5T1D7wUu0
HeNMRgt/HdJmFhS9sfqQ+6OrV0SaGrLUoIKUPUSSFeJ550vdShRyWeL3WvDxkRoTLMknHwwhLsE2
rQitR+LL/HGFVMOTvNhV/MOypOSWPZOIRT9+oH7fMXLQgIa3byiF9nlWyjrF1//ZSoriBWya+EWk
GX4fgNZkMCSCFV9ZoPk2vjrI6vn+J5b+pYFJA6sCaGIrxnEtisS8QOiZHzq+Slb7SVkHovDW2K10
7CeTbKmXTv5RzXqEVutUfVZ8aXm2nJcA/R/HmWgLK7MLtUvCQ7KSsPRBqjbrH27jXml9sNX/PqZw
sp7ppiUY3VHJZXxG5XiOIxn5zugUI21TJwBFQkHU+AGuj+THGg+kAKfGprAK8yAK9FLNurGySjOP
69cTa2oRTjPuGBMSG9xxmODXLahvHgXlhzKzGgcEOt8VNl4GSNG3o+sksYU/E7UhL/mB5gTwkCJT
LCOCpVd9nz17He7m29EMZe/OPkZB2FORYQaexah6QqQf8JYLiXv86fpoQDLHY5oCe/52xhzVLsJE
u4SYPHfpv1mP1vdtomSlza1V74NfRzfLDAdTK/gf5GFOvNcvEKLzgpk9XxPfyf0nfhRwV21B16+p
CKdTxj6t/MWDYfL4UOyIWMX1sP2zW7915F5qPdFsWyGwHqIiFTAkpInl5ZtJP8zuIczXbqeLTlHO
wAy0WzKjiQyVTgIfXXX0r3/lun+vPUa42hIxKCahm149RQ/P4+Dc3/WztCwXpOKGwliArdcKwOIV
sXpepaRAAXGvfBl7o5gKUiTN/RqbH3QiUkc452u7yo9rbgNbTOO+hAJH6YQk9b5AYlf2sFAO/71+
1iSOo70ijmj1miX4JcA+IJFKSI17q1bNZdxdnaYEs8EDwh1RfMpAMrNM7UHow5gLfyzAentUysv8
bRw4n4/GwuBkiuaK6XbaGxrCIfb7ALfWoIRkwH00yGIswIz/6d+G4CuDRlQT4he8e7TlRwL36O2A
mlTE/AgUkFiz3qQPFA90mo5v+mJd/1hypf+MMrJ6ktXL6RzZXBlE2gCnWeP3W0eE/LR6AaeQ0RRe
pnUBNs90wF9PuXPYZM1zG8jU/p50+HjUAIPFCEaHDzIyNLl48peMTmlSbD2ef2geJV3CvqpVnAIr
RzEBm1fQrSRbrgvF77wQ5ILtm9wjgBo0ywA4WnV8oc65n0PDarpq/ssuWRKZF0pKb0j5mh9QarCS
A+0b84Qz+EfCniHjUxFG56lgfm4GoiA77TSRvHQzgj0jREkwIVElJgdfyWEG4Bb9RdTCZIek/9Wy
TrjKiuVif1HzBwpUNjqrW6IQABGni0jU64X9ejmXhl4JpcYRa/WwEeHPQJ5QiP0e7psW8lfkqUE7
Eh/eApUi6CKGfn5h/QWRii9vuh6/0wL3RW2xle70kblL/uBEDNCE6OrqcX6Iid7hPiiiBRG51hIF
1WZLE/q1WKfyGJA8Lxrb7zC7sUQnkJRhrd2SeU7JT1xGoQl4arr2siJrK9COLyW7O8TXHFysd3Qx
/cFCKJcuKdMtsdct9VeAiuSDFNRqmn3kMgxRdAHyeTuVtdod5BncaEdmdbyugRdJFtCGZPDdKsoe
DG7bkTJ3rkga/V8Y6PXm+DAcVsAAi+vJxwx1ytHoBfffbsVz4SBnyTPVbqKD5xzbwDJ8snO+vtzs
2C79wTnG4cqUnJqjOUEWiEcOu0vR+oA2Gtsx0kef7naPhnZzOAWxONKAEl76qg8kCdg11VZW5zkN
WvZn6qTMtQ5x/J0deemjR3ZANxn/V5LwORJo6q6Kfdc7YOmJqGiULx0+K44FsQ9DkvjfLYJE9uY6
qWpeidkes3wPHR4cDifOEuPytIf8Bs/5Y7Z290W1hzqWEAhzllJlFBHSgpc15lLsoMM8R6vj6ReT
5qVwMSbYlnEA7M+edKk+DKLF5uQM5KRAyxTFVLC/12xidzFLBKxlhyNnzQZOuDQCjqT7L9QNXsqi
eBd60/bik/W1KPCfw8iNii8qaYwZqSOPa1fvAoUg1uaCi2WkpDH6O28iQgXLNC/rm9FCDM9rWJO8
v2OoiVHfyxJv/A0GRxG8IDlOXFY8aPJoMXSz/5A4L+0idqHmBG8ExNAnLe3zM1stbqXRNM3+iNST
UtRdHGvgAnLhEJOAjlGhdhRkAzlQXM7k8SMbPpIZKe4ehK6eCgPmthxJN5PNBNaubjb0xNJ/2Vka
Ay7C61hM+aMaGNHjx20pZsSlCozak9dXeav1Ty58WNFLzdsgB/vvj5ulGNfbcdbCCgepQS7dJGT9
9U2TdcBXmn+lMdIxGBDlGxFpBKRab5WIiuHqFIPbA4AlpoZcwT+zRaN0Pozw3KLGLFyrvFmqbINo
LmY9p0ymB3/t7+uMYnHr7PCPy7HHhFm/cPSiXU+AikSU4YiZoSPtP2WL5eTvhZNUGmWnd8EF7C4+
E7QxsrHZ39Paj+T8u1z+ytiwpCNf33nLI8ebuw6IuRXeuEVVdL+cofM9pt/Lp4Y7uOQ5Qg9yY8Pu
lzTGkRbJUbBdB6SXFVrSmuAASSr9+dc1aP8WWTH4IQT7nQBXZuGU0Dcd5ciQKydRjdlopZFWxsBS
hL8AZOvMBZlfe5uv13AGG8XskzpmYkIa/R6hFbdE1dwvcgNj5YAWrWGkIAQSixFwOqt/BQ1yNTFw
ELvggUUEoFyTUOkJWGVFY+GdzEG2sJysU+4i2g8Vcc4GyvRc5HrcRBaOxRwWnlVfle2k94X+RGsO
ZBWlDUPfVolFcDxRjCC0np5gEonv6qDxEQaBmsgCAEs8sotQ9RoU3VwpTAJ+gHuR1P1mPZ1pPcCI
GbgU4+w4Jh8rhy/LmHzK9SmDvn0JuTYstgTXv5lAgV4Puyws+1k7e94SUc/u2j5W88ictJZnQcOi
3veK5hSW5le+829mpvx0S7229ry/HmilQ1UMojWLjaQR/DDiHMshA8kzksJQImbeEhljNmI4eSv1
D8vLzDWMevcIiCRmbPrVVY9YfUg9pVr7s4gkHBLJQk6HZM1T3Y3TYsxgqgUldOlWYmMZ3SP8i8Pn
STC5sWJPbhXl99g+pOujiPH//lXeNsrz9qKwCiPXn9IAC4m8co/wlhxdYVj8vBVDNYoq0kh6NHqv
mMDVDrPT/3972e5AZhFWVNvX+27uWvADVvaUY73Gmd11sFnu2W2q2po0Wa/4ANYUMn+vgNVysN0c
duJNlmvIJA3CUjkfSsdgUPdUte5209p2HsRsZXKmYKfYaXghG/fQnOw/IFOz+x0D+uWNTgYhNAvF
dS+BOtKilTmtjP4DqD2bwqGPmXVLzO6zJLCya0WI0IGTLwYKWyxvA66uGi1395qWFyV9VSnsneCm
dUJk77Zi5XkTTCJvoXrMxtGhoYY/O4zTSbMokgmM0SYhAFf+OMD2jHUn+M7zU+YfFtgjIq+T6Koc
kGxkdVBiWAOfs5f8qG6jdE+7bnLJph+pTQlpDuVO9YeiM4qNSMNsPMHwsLnKonAwmpK1bPukLo7z
dUAjlDy50CfLj97GSUtmc1wvV+KmfkZonLEYtZCtPI/nyfeaxHmDu4+al49rERG2kX9aAyyeIM00
tXHlJwEVrL2mCn0nTSOn9QghFczDtUNarYNN2lTUtfe4LLa2oOU3laj8f39IGAj7uXykAHMN6vLo
xdymmSK00tuTt5HWE7KZWrqWCcTZ8uo2kp914Z06wA/3+lGvfGgjLTxTsUAWG8QEpdzqBQQqxcdJ
VVvI5TxNofOH6AN+J+kj1bsjWq6QKVUDUlAZvzeOKZKOd5E12mPaAGw9229LujAYJgc7LuFODdIz
3k2WIoRWSwKMnQVFvhm4DZJoH4QPO0LUixreba6WuvUZ/JKOUvIaS9Hw7krq1yM7F8kuC9p3UAai
eyCoim+LDmTySFD/tlWsnviO1rHKwQQb/e5ySJfOL+CGUDhlOG6O9KLc9yFZp9A9JaSn000LbVPQ
yDzbBz5I701DYv/ZEW6VehYvpxZ+LxkeCoQMwhdPuvOXf3e62j0xjdtk9xb4gYXU6XpjQXRTXLD4
FmmN8RNIR6szCkorO5SyJZawA5z5wGcG5YGXH2Lmesk1I+fQaTVoRKUxB2RNx9BHqT72XE6wmf/n
MN5lKEt45X8NXVzsm37gGkDUBjFBFGz+gRwADRyHh4ilb78QDzj6ENAzLjrge+VWy/2l8PqEIYOd
Sps0LDM4YhlA7R3pnP864NEy0utPK5hr8Jojyl0do2O9q/z2GJDUyyzwUpRZDVnumVhDp4Y0jtMv
nuAeAKRIqm93A6ROxJsq7y4i0ut/F5LESFFi9MQSaQ58BJ4sY77frE7H8c9TK1/Xq+fNugMIRfe5
Zw6I+l1BTjZgpttQDb+cQw74jK5uQzKwlPqvT3U4aYEEt10IJO4KP4B1gOzoeEAY9t1MbyO3/LHn
aIyvGpX7FCFnPJujYBd6M9ZWus8XQikEsxaPtHuFCjdXbndlsOgQ64LrMYUKKWetsZZ8oO3yf27T
TGAxZ5Z1mGCi+1X3StvwafsoTmfUDPxiYArl/Qng0dbunM0K7o+ansiXF0NO5CsAgKdoaIZe0wxU
IaiFWC9x9jWzfplvW8jCZQUokJ8V1laIx8ihGl1virLbMEFRUjMp5yHQEJ3RE4eCq2ta5FcffZ3h
P8vSV50KIpS0g8reWpc0jnOenRws6cMlnlC1I4DkWEeT5r6RR/lzcno/aLOwJkp9PRhXRke6VJh2
1190p8qbiG4Ip8cFJWrrY2yg6llDqIFM2xZemNYJR6Bf/An+rYBq4CCWA8hr2MRuBOksqRHqtdTj
FXBxnlEdCNTn1Dx7xd9h09rn9LoAO3nX1puElY0NDcfi98bVUmOVyP6UpXhzIPyDjm3zC+7l7eIi
oIK/qEIGXrEL6NuOHVhA8bD5Pv3CpcPvx0aA/V+jhuZYx3ZPiC8r8SUjANvq1a6A6O55e294nPwg
e6QZY7vhItvuPn9cun9pSVLAnVUK5xqDqbmJhfVW3uERrVEVOH06NRPVYR2oC5KSCHwRnYtyyOil
/7v9Vnx/BIyLC8ZM5qN7qji/ToAofL/JuRNYjZC/C35uIKhAF7zSdNqOYO/GJH7bcZsAB0jjeGBJ
YrJOFWgDp+3ApLPEHbZFj8kO6Dfh0F3Ac4VQS8vpP9bFRDxBzr3rWVXC22MiIFYbCqNVANi1YVrG
o0ztUtsSm43CbeSHDPsPW1AzcFnkuT05TrYIZki6tdjSF/sLh4OR9vvYdDI4OxZc3JJcvi0+/mrS
xwOhuWP876wvYEcHA5vG83ikqQZQgjhGT/lzNWu2kjXLeZRbOdi0V9SYsI4zj8KRBkXGcIwW2SKp
9Dvy39y7YhLiRETaG2m2t9EfSGMOzc25HgWDUc7/3SezgcTvwHrxGJgeREI6rR/9uOQImQ0u+7a7
sjRZRR889+/8gPCIrDIWZ4AzzrK+KIu5Ba4MznwDemUK/YyBnV43Mn9AzvIjTW8QT2XehLqS9TI9
0h95kWNh/eEljyQL4FAxjUP8d/BBCw5/c6b3l6KDOnO/qwKVTuPy6YJqFM79/ycDGR63OMdPuoHs
hwYoBhzueaemqz/NnSL039cpbssioAFthit0FU1g1HiooQCjmy3bdWWzaIn1udwD27tgXKkemQuB
55IoXFxDtnfTk9A6MUMVQsk8FJZ7rD1t2UIzwOwLkj4PdBzfDtZjeZKbYxURNwLh5eaynsGWJKre
JcozJ/CB3AYbd8jo6I1y6KN/aXQLRMeaPLMMDe0VWu9IdXJlhd4cc38YfRqxTkFyHQSanYBariDq
vOJROg+SavUJAbxsYnyZAkFL3H0/6MOGFPLin4URtwAntvQaXFDXDSURFtA1X9NjeoSkdrOIwy8n
vQh+I1QqPIp6ziYppK8fu6YeJKAAKeF4CxHHe0gvAL/rUNhkS7KsqJ/GA/gJQa99xBQuUv9mZJXO
HPpJX5nXTuIYFudysk1lM1P/BcdnlsrJ93j79OzW+1K116NdtTs6nwYFxZjjicbDVHRiLsoWxno/
TO1Do96GglMGVLRTnBtrASH+q2Btf6uS0AbGESrULYy7EChorxt20AJHSikE3SPobznXjKJt7GbK
meIwNp1/4Mb9+82w4gFMpg024QVACxBouxZY1wJmIC/LJbqo0GQNVNRUJoJBPOG1u88Q5ScJ0diJ
GsiuHHnifFbtrZH52bFBsou7kxn2GwO2ESkl7Z7A0VIQk/dEEOhY2dfVoaApMGHLuIKiHivJuCPj
JowcB12aLYo0abOu3RdAsKHgn1AT+HyzQ0X6a702IS5NFpfX52Fd9XKtKsgIiFIdb9pB3+bdeoW9
VvrmOhMnQdKg7t3OCRhVrXs/pHt+mKkVRmYM92S/9vaM5M2SKMiIOBJGsdHB+DDXw/iQFM6747In
zIBQZ088drH6PLEXQOcV9aX83RXXMtntiVDZBiecioCN1BOGdoZBIEaraSJMRerQr5SGcbtJDuiy
mm3fxefI/ShBsHZfmdVSurNscdj1yKK9u7GLRAxl8jQNAMO6uGAGH2oOnkX131TAdUZ91yuAXV1p
srj2+EmcHyDVkIxfSoFkFdgHMzEnsldb3q4Iai2DbKr6L+LSTvTcgpJTSI9onDgJonAB3z5y7BGt
O4ulcDLsZHu77G+cyJ+U3eAI5DOATp53rFBZk84dd6QwmR9BMPRElWfueCZyyzd0tAb2zhGnHQn4
99IR18On18kCnqoFLbrdihxYVi5Zntbmz/ucMLD28qe6e86ukvud6mWG/lq8CVa50FRvLUl2m1fi
wBk1CftLdMzcFdu7uid9vau3IYHvlT4XCNfYW00Mmf4eRsEOgM4Sm+511Xdqb0IZwOOmTodLssIv
pgxLBAsDMAlVvjRoBAjpL53aUK60XPpJO6ZpCEsHtpM4LOILpUzNLH4P8YwdByJmy2lmCKSbxNN1
A9uvQ2/yZ02hkRnADRyCw7t4vPycIkGzDTwodHqtpnygbiuWfDneJ9kXZy0bOISPs+/prPS52978
XJrAS0QNqawYc+jSGlabaIitjo3q13++jcfJKqL1JA2Wu3m1DKTfhJaed57mpRVHsVAiLe4NxUxO
VwwMdjqhIr1qXRen3hoE6ukgDe3LtJDeN4JjGF1ZOuB3CAiYyhhzJwdRB/IQcXgkzDluz7dm/cYe
Qhb9cLE6obps3VkYzQGk6QAk2PXBqzdvWAi6AigmPBzRjRmJtdDjAET92H6Z/MTZVruaYWYda+XI
YRpey96G24RjIAoCtwskjl/Z7TQ88GjnGSYAOUMwkbdz2+CGMF+14NtcWBGDLjkUSRcOu5/PIx3i
GQuE3ZZ82J5sy9n1bJO+or8Jug07QnQMq5dKf16wmUNwv2XzBz5aXPmIImZ8EWrSOVnbRCphEec1
ZSIpKQ39Wm/vlSTfLjjitZ9C0SxzqiOJyZd4UBRC9mNT8UWPGOpIJ+GD7w9UgdaxTl2zWR3sXMea
XhZ4xzqd7h/PGhlfG0oFE7/Hlo+uRid1ln2MjEZLkQ4kx73kptsaqYX28Y4ajvk70MAWVDIGTq0H
nLNVNAe48ykdSCtNDHLq5MX7DZaHmmslL5sNAz1iKr/CK2YXTQB9/e5uBrsbNWOZcZAOS8Ecbo82
uj/SiKMmAO1Xm7lbD+bBBOGApPem8Hrp5EQsvoiyvZg7ZOrvLkerrBxWcPio93Sf3hjwAVDQHjVl
dh1CvvrfYjl0KlwhpxZ6/Jkr4RBSm2vJ0qtYKLcfUTo3N/Rk5qD/ZJJbnvwi2T/xhABmzCG3D6x9
hkTAtKxdRo3gxVngtFCZo89NZ5DtqSESWX3SX1xGwLoRcxPDNov8ExcXsLyKZnA56Jy3MF9vionA
1aRjyG6TonC+bNBPLisI8Y1cVLqlW3pw4J32hWyhyz/LjD7FYejpDLJZo0pyOhhz+exyfoUt0xAS
4s3jaTlglBM+rQ8in29asCxPw9H51gAkjVAPJVlKs6qJJW+ZaIqqqCjgm0tHNONYOJUSjMyDd97t
kDqM80Ohrz8NXBTw1eac/hUclYATiBgZAErqT8P4mAa1an3lQMeFgbLJVMjsqfN7FExpVpysHY6i
FkdYj+0mJxxz9gIKACwYaOWkOJ2Am0oOv/9Ynj8FVdm6v2vGMYIA5R64OhoWVpmZUKAVQ5MSVhax
KNhgAY2t1K7UIlGYcYyoaPhJkPCtxV+04ucoQnQPHaBgi3aUXpcn3gnOyjbJcJwT1ZmTFWM9R2Fh
LLf+1TL93iREEA9rpAUALahe6q099ARXNR2ENOlljXVA5WNvl6KqDoLBx9eZ4t/ER2qIbaZ9bYqm
9Qq4YPtRvWyd8BmTYNv2NFrdc9GNfC5eZOxgORY0BXAJuAbTs8BkN3QrbLB7+b6FnMKbkLyfsLFS
rUk7GTCakM+N8km3tgS/YbuyafoMkXgM5qk4wURccM36dNO/Z4VGjSnsmnu1jZ/mLQ3LMaKXgr6V
i1gVOhELidg7bQumeauI0mflSDNX8QfkUvKRjeMAwwlLY4F343r4k8NwvX/TbKiN9AQVjQuX5coF
hKnJ3SUkuTpw+jaBenNa1wl6HXC+uambXJe5y3rlrQQCR3gK5KNpW+r9JoSFZPUTQ08nHSPAj7s1
0f1chFFnWHYGnGnAV8DCQ4fAcdmLwIzBrXFgc00Ulg+Y6/PU3x2XvN5US1ZQ7pZQhW+BtpYkKd2n
ma1WH7kyK7GTA75aRKwzBgifrM7FlPYz2Rddat0/gRVvZvzUTLYsqRxXZj5aouzjJlxVHvY3JWan
I8DbW2cEUAJhe1EWq38n3sIZWXBaxF0nnaSZCwZHh7ZiJQ+hccpjvSFIn8qOgiGzrN4aYcyrYLkZ
iQtjFo3DAaAIHEl7iZBSuYQgyg2aY61usg2u2QUQGwdeyQFrb+3W6YM44y7tCzFXBgyrdLfme5ja
jybCd0oLn5xuI1PeBZz1PH6B8CApHBP57Pk2dMqQIDfQqzysv063n802Jv+QUsKPtso2qh1oJERE
rPixNOl26vJpe+eFTe4g57DRu0J7JP+KH+iz0qjvdAwLS4qfHoaxzXKeSrWoJ9w9bZXW3X0YP5DF
kS3Ff6roqnX/QGqfrjbJiLcBP1Is2+H2SrERg7YfRhjVoObI4LchyqPSyj0nb7ufs+6f39g+RFna
g8OK0PidfFkPP/MQqpdD+K74Bx8y7U3EO/9NnjfOn1/6fy4u8sv0+PdJQy5jHrtnvnIS6D1nRj2U
wedrrmhyvoiVJj8dRoYf7g122oHdRe7t5Lec17oRx8na7nHJjnapd6wNwK6uFImZa92zJYnqmQWM
ZNlaHfuRA+6Rd67QQbq2Hc58O1rATqDzs2JiiMvwvOgFhO7puShGF1n4ziSgwF6oORDMbGLoNMdv
/c9E1s/NeQImC7tq4TuyAoef1AudGsj5lBp7f95IQeZMn0DHdUIlqOVxRK0L7Ms/TXo968xaAXqw
7Y3VdAl2k4BRFpFK7uRYrPiQE1j28HWys2xwQMRRAeZEr3dAzHuWDt3sq31kdBtE0feJnnCqiLFG
E+HdZ7KEFF5HKfO0STZw9iBh/tQlFN+biXWf009Bj2PSvfDRuHwfLZQUw8ewRw7bpGH1mXsD3DeM
fyiZXAnXrbhkI9PgyIv016a/ZgZewhzUSDm5xdJ5xtjPWH3LIipflAZBrGySezwX3YctVRa+tXt1
3fAErpLOkSIT0nam92UEoj6SFnCCX5PeIDPcxTZfNzV+nSG6AycLCOq8DrGCY7RTAC/p0ohXbkGw
qeqKAIVXrDyp3YCIqq7782KfCwV/vYudbj61hVs2c/5LW0fuDYPjtsn7b/e7G3fv7eRyG5cnjJO5
WLmW0/jBLHEQkJ1PhYnTZJC4MWK6m4IQRVI6AESRoWiYzKYyPExQ9iGykEZrYm123aNenXgCFTHZ
UxccYNG5UwMB9jQjqt52xxtADq10W+fcru6y2znMTs2XmZg24CvNE444bzLBYGlob/3Jz48ey3ks
qERFloycIJCzGLGLl0NECW8LzSP55Q2zyldsbSTd2GHGxWiIMK52MXvDCpXj0u0ggzSe9revwXgo
FHa7zDGHgxT8ds3IrxhJP5PZoPGGa+D6sAENvOH0VR79ZzrWnbkkbzArWLh3kySpFJZ5qfGzniPo
4uV31crj76bEEbvJTJJkdKzsMTXH6Sx/vdmU7xum9ahdIcJ69ckOurZnwjnikLfCzueaGkf8QFwK
SCT1ebKaAMbTgdO2zC3IWQzVqyZGlxJ6YTG5QFmrFYX7jUcScO2gXrQX9tXLbGmCv59NV2TrcEbd
UcMQmZd3DK2Tu51mehLzfXte3XUWZywM8YKHqTn44gInauhseeuYqJB5HNDEtnODalkklCExPktJ
6HUyuvSZMBXC3MKFmL0q9fAh2CE9OX8OP/kHMPWsHIaCu25B8IUVljHMJfk2eCTXsAqlh9XhujT+
Dcl6WoDOIzgPzckOvWDw4+aj4RWQnf9Jo4/cExUWcg5LghoZu9NAmDfcan4QBNA5yda2b21KHtSS
wRcIxA37lnIPGsjNfa0vSFUvE505MB9MraYT3quzfo9xqvwL6+Jg4+rHfWK+cSn+ZfOgwBkad1DC
cAZDJirVyHamfIomJoxSvSW4dsv0twEP4lItvWqEPbCZJAcKXAjfT/Y1Zvd0JIeTMWkyIgWr/MUw
Ov7S0pc1WkKi5+Y6nUm4Ai8vPqy6e8pBoju7LHmnEDXxnvRfNO2+grs2MTmPujbVPwZ6/GLWAfKd
w5fj1zTt8VQ+CBO/GXxVRipfPyqPB1xtwHkZ5ukzrfd7tuKRJH/sQt60ZF4zw8RMLRGUo9QhjzUK
UJ1neI5Oozpw+Jw9GKcq7JjwCq4t6m+tUBSicfJvZ5+EUnCaSl/C4lWwVWjPiW+gm7UJseYcx0Vh
bMbqUwdMCha3Q8a2TMLZjsjn/r5f05Z0R0oIek8aC97xZ5m/EBc5OHOZEj/NK5nrkx37x/5DecfT
KN780lqTGMspEGsDZLvz7v73Zdcv95Mcb6w5J5aYWsrG1z/M+FYlcxYiVG/nfEioGoi9DOxfrUbY
Gk0k64m9jc7o9wkVoS9Ep+DeaH23Lo9klVijKGx1/wjWEMj9Owe8JwISJUeVcQKwKMUK/1tthZ7G
GcrLbA9h4gHaLwOn4zWOQww8eRn+mPiyonugG+7QNP7AzBykV2saqmGQJMkMnJFgetcMwUfShvxQ
CG9hb5LOfNoJ4JktwpdoIHuH0j3PnUJUpJ0qXRVPwyQSzxnjnhYfOwDH7Q+ACVRVpSfjFCdxZ0CU
wfjDldqXM5nOn+cfr1nDVdq8JC6TMCGCK12B3pOGTQ7FiWz6Mp0qbOawUiuRbhMU+EPO9eUAygZV
nXGfimOuO1E+dEovO4Psyf4mghrE+e0u6PRN3Hq4100EcSMMFLi0QWJmkshvNzkgQnRubAFLxH12
MB8nirl1th6KJNcIeZhmKLmOF5s+EBfeWG46yuU3nTYZRYy5QMffFikZYJxOQFaxGUQiYWuYPtK/
54WSTeVwlWXvPrqmpqhIYxm318NYQABbgWdKotoLWMpyJ8gvCDRrpPz5N/TnTgfy0kg1sZNc0XXB
3XkDjC1YLoVr/I9AzU2U//+Gh+DtvqEfDLnsFgNny//5XpH7jsZFL+ThIXLFlqXf3tGjEQUfpu/w
BhduV/zqo7tlv2ydNeQkA+TeSMgNVGN/Rjvice55FDUIYUX8wFWcFPdWkdGiNgbV+7jBVCrUfBkS
9Hlk/rXAyGza9gxX3i+gE2HUoL8mmYCoMAgRuC2uBK7jpKG3X7c2pQsS0zXe2nqTGcTUt0yVYeEF
otkfRhhgDL0zPosM8JiQLL/pra6fWTRIGaKlwhArqeSANsxZM+KjxR/AVuTIkjOZKqGgbOQjYWAB
s/rDcBtfIZFHxhyqksNnrF8/zow41e3kHCSgzf7EQIHtxwjWW5uw/bpvsupxX0meJvY3Nb7CqCg6
4q9y/potZONXAqn3uN0Q4h6BuVVkv9CbW4h55wJ79rCzLhsuW7bD/PqhFJDGlLvsYPMvX5EBdnxr
h+QmLLOLt5qMaTEJuDvXDW/RcfP3MvDD58VmGYEBJRwY0EheZ/trRkO7Zuvl9WNtLZrxyczG03+n
AEEUQ9VzCp0EdepHKrSGCflLEOH9r4GZ6o8XNP5gdcc+0wa5egizKOn9Yss0F68qTtxTWMYuMBz/
u7Vm3NqDr45Y116K7yCcQMGNWlFjKQW9twSJE9orWiitjfrynH5TKlXZLg7yTDCjsSNnp5Mz7o3U
/AlHe3zcyx7R6hu6dIg/LV9NnvkGcZrk0CEm/RlxPkIxJMcLIxHVgPiqThV1bUDRZukfZpSC6/9F
O+a3rinKgwolOD3agIqH7BwEKxR/H48YNHKG5A5PIe/g1NVOPfVrxQ37ZseRdnYACPaEdWs1po+m
37DF+LYjReGJmkoH8d3pZ8fWTtr3Bs7YUfJTadbF85f5qldHF6j0Co4MradeXZuE8kppiYf2JtOS
Fs3YAu1aLcbwEZsfdMu/Zl22gXPKgh3mZgCnPibDVHzvwxfx4ZIvQlJR5flxVq+o6abYIiifvN/k
0ja1SnAIT59fPptK08UwatuSZIQuOFv6PfiejwRhIJ1fgxb/FwM2rBC8nZesentu7QKD6sIoOY+Z
tpRrk0y3EyxDRIXKKmxcIoPdERQQaK+Xkir7ikyvGuBqXxmocYSzoL9GPiV1
`protect end_protected
