`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
bx24XPMbQl0ZuYgzgnvmK2UJsn5v5rHRrHaBzymEsRVRAjuRN3xRCY+goyOwSGiaL5BZpex2sDSK
2sd0nljSnw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
CSRfZVLMWm0HJLEB7NOFzWrGIhgXL0zMCnVPoqKjG5Ur0+RK898D8TnT1vzg0/m9z9AJo34CsLar
7ajBwWmQaStI2T7HakgiApYlcuC6de1XuIEH3rZRMj/RWcjpTLbgkrbMj7lCzKzQdvZHARVRsJHt
n6KxqqDLGxMs1/m4zV8=

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
YDR4T6HZUUPDmkJ3uEF/8DG9RH1KIm/Soi0XWVOdqKCDBSgk2PKH3QgKdeu/Ygc+E4sEfsdQ97ZX
ZNKLn57bC8vQMoMyVXHXP/gB1IkATHDtiORbiLIN6gz0rbLre/0AWJ4pnD6+ix+zJ2ZtVx7uSjJD
UeDwmSaYOZQhEg4QN3w=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
b5TzJrebbTGq/pRucwAvmRYTRYSTXLJ31UHhj7qPdtWGaTRXaKbjtJHLK6r2fdEku+xRcQgb4iwR
VR2WDz2dfhkKseFS1Yxa2DFJTK597UszihjnkRHDocjQO3cUY+io6Cbq8kFDe4t/wEf721IVy63Z
z1z8RoAbpBZZGG1+seGG0kHDtkTe8wOMD9mRo2qsutfBPBsV5sK8/fmf9Y9E2sAlYwKjVvsGOjpr
dIS4pkfWNQ1UbQXn1WlPTe4wXcRDxSDWm2NMDLpVsB7PHxXe/ma6En4gcBeXFN40LqU3TWcyfbF4
Fgd267nviONJrvDRA6uaiECsHX40iXKsaxsGyQ==

`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
LoXyfjLEjXF6IqzWN8H3K7nR07wwyqyXVISYV16h6KsboFmbDcRTEPo0gH2rwN+AX6fpfnjiQCDi
qZVj+jq+3Jpyaex4T6xZDGqASKvTFZ53Vog5975jRBzfQilhyEnt1jyw4Z0UhtEM8LILdgabJqA8
cXdC2MS8KixvDgzWP6ABnTAwC9pDqbLUIqs+coqVvcy1nM4qt9WlS3/X4SHWNrmKgZ5d/HUtKouY
9yGUMGTi2nl4U+Zd7UaI2yJjVCW8JLst+BTCam4lPyVXo4ebpoEbDK6tTwa5DlOxI45b/ZooNuYE
Rpmlrdz/peCtaLTTS4+P11HF/WIAxGHuvcXpOg==

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
splRKPjEH+uTzvqD2tjFWmYXGYcB4TmcJH8LhGT8ueKKhMoa+orNkr7mpiSfxGo4nOfb4ddB5A74
rXupMEGR44uXFXmGFms0uV3Mo+LAVOswYWiSib2qqWdsJAVPQV+uS8kwf1pFIhgSfyhJYccE2+LN
qen4ppn5nmwPuAnPwhqNoxWgV6I1SCeKHMvOOim/bGhWBFyFuI4F9GeL1p+BC2DYSvijB6DHJgjd
lmuMd4WuXe78W//Vv2jhHriZx5nGgRFuRWE3VBR/38AWtMEOOrO4ijdAV2GyHZrphPmDHXfSwU6z
9JSFgLsD3Pd9zxwPDkqCeFOIFV991nTMDEBaMg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 16112)
`protect data_block
McOR5osfN7FhwOeAmCNp580N4F+RByuH7EvhgYojFcBg/8vpIuQzG680sV7weUct28y0SPNs4e+w
qQ9lTSMAdVIcIfpb7kmuFm1wYejIM+Am73O6WYKfbLSXCEK0ff7fudxRcaw1CHqSKP5weFNy/W3J
xRHGYa3n+7/drRVlEUfoidLOwXLag7w3mk26EFheXCHy5zKZBEFdTDAySFVBOQMKnJuVkr7TSWy6
+HO0S3nwkJb2t/2Obg+Gx0YFDulb9lgpvN5ucQIgofgaL9RLMFmlT6WC0QoQ0AaSw7/55vDDzjDV
jaxpTEajXxNZYkEWyl0jlU30mSGCjVvm5auF3L/r1FyUaXcwoU2mKV8EslyjmFHakpZLbqsULgTF
Z3RCXvU0B3gSkWB45UlnFFqWlHdxAud9ph+KM9n9o0n0b4iQv8ZCmtvmffNXncTx1J2HG020+mz4
Cke10DSrkd8eQKWWnTa0Yidx/iULtNjVOq2PUACrwBL801bboIvFcqupEhh/fZaI2xiAGGJ4N/aa
mU8gjWZ+p+mXH/5C3QrOdww1gXr6EDCOBrIjrNuqNvETCyVsU88lnIyyKpKoSBywYVqvlkT5g2f8
k72MoagO+tyPqA5fY8TJdVFc9ihx97d5gB1ZJxMFPLhbCb2uksKeyASA3+krMvdiRaoDYgs5V1vG
uLzMuSgAY7IbL4Unz8FbU7yyoOM4I7S+bZXAdGq1COUITbk/WxmrTQEsomN9JtZbQ7650Jpq42Z1
PnIaZSulvU3KpmvKHMv8Rk7ds6VKtHbnwsN7E+bMmBTMhEW9owkRSXUC4H1puygq/SQFoAKVdQqz
z58uDiorVDfwRTL+SmykOihbxcYzKv05VIAmgdlxlwPbHZqZQAvPataV8bOWaLAZb3XZ7D7r4ehK
A4MP3YHhbrPb59If4o2XFOzsq+pwXkBQ0qo4X3Mg49CG/U0tp6Y2ykBZ7fpY0iOGTqcS3AVU2+Bj
V2Yt0f4x90r++6CuqRuVFqTfGZtw32KVn+EJ/0Wnuzfeko0TrCb52SsI2Qotvu1+WfvqkC+vFa1r
B05waKkVC+JDjJK+1opjXByZAk2otJIlOvLPAmNsOS58UQWdW58tBnCH4ROtQC3GoK0lMghVsNQV
kicneUY2/YZ3kMEJxH1Qjui1GciG4aRExQXzsGax+AO94AXGSTUzEKJUZdW/KvVjqaHFhVcanjPg
/umkSSh9iN1YyljLhQZaXN5wwTwb3gX0xGl+rWIA+AGtrgvDcoNNgnjdRBIr5/imM4mBnEHcazfL
EkHeL1WgffEklnQYqiFyI8Qz3czhYwkFCUVAZDjj1TL5m8pBBkQEIlVWfg1pVubC34JG9FVTAhz5
SLtyVzKu0RjLXTg8eSW0t73SjaUtm3uZv4YlrpLaaa9Qa5Sh/Fv/6EBtRTjY0Z7znDHr7u9dyNfP
rjrjdqR+S5B3eDWda784jqVebprfV/u81Od+HS2gWaiQZxc5y30Tg1EGAumXzI/jwRHGck/4uUBn
WyKLBuHA4FQi6vpQkYDzLzHdskCuXoZ9Ovn8ANicU2TwDfqSFAue0Pb2adM7Jz2lCQ5kWkeSQXsJ
Qw5cBwWPsdPtnxsn8g7EeLslxl/TS5iZwt3NEq3MBheVs8/s5H8TwA204ok3uz2wNtajWvZBoYpv
BtVvFop7tAnwumSIhkZxx26oC+RhM/tX1osNh/8rMR3NEeNE40iBIFWy1TY3/btmyBdpFGtGA3P9
0VaNky6mopcpu8fUT1vqkiKeTSfwRRjjvspmn9pmBbeKLbRsDJNDP+nywudJvyj1Qg72IjHWRiKM
AGsSFzW3upoCS5pIWmF4VZEkRf+TNeUTF4Tk9VMOoYeHZciTzFCr2TiWBLBryxPofaSZPLhlT3Oz
b0bAAHWDv8XBvLj7wqlN9fAhk67AaKeeziobtPkcRFiUighBBdUBkhicwj6yUWjTmyv23SAa3/C/
iOyrPAYtyUNv7VpVzN7YlZDmK/vCEr8dp2pXm1XRTZNGiVURwPHlC5ESiN24Bw6s36ZHR+TAH8PC
AMRqKURiJXAcUIYJTmTAbekZjHbT0eEDiRQ8j8QIoTP5joiNgmfP1HaINTWJmi3INHBy6lkrq8k8
Zq+3rIfRRCEqR83tS+v0/XA6nCPoSKd3tmWknW068ye0Knpa+Bk1Eu44DpWqNXlAMpdq3EeZLomY
1ksrvZM3mCU9IMCwFafunPykHepD3bu6C8gtp/hv10VD6NozhoyVADUyikWml4+TUvJdruQOpfgx
YaOPSVZVzqyQHuhJFrhtVKso0JtCHqc2lJM/67p9G3407Xcpi1hobsToL3YlmbwGmL29++Q9bff+
O+ftK4ym5W4N6iIUeNObuD2ysUJWdM60S0GUeq0rn4NGo8gcxIJvwpNW6TL4v3lW0HpkVSQ/hhFe
iQz3MmUu64ESBFwD85JuYkKyy3ZASkZ1RIF+XMIo8ZqPQ5bYnPrTlm8JmemBo6qMDaHGtyEJkCJz
e1rlzO1y91YtGvOaC+oHaVCzP20rKUM/1tYWMn0gMCPlZCx8LPGsK5Bj3UE/4wONrWiRUBX7E63v
vnRD7IjnT57Iog8RP438SGeQCzTfIyaJxGhk3UKSZ+dnqafULID26RoyXCzJNWHYwND6XJSPfq4p
qhlgkR6I+gEWIFkgIfFJJjxUn81gs4PDRkh/xLNMSLeWSSfPrj3d0ZtgK/Y+qXEOZpSGFMec/86W
oNh0rTX1HI7IgLOzcD2A76QIglPjO0fJPIIiYhy+41Se+x8A5QOdDQp84fDtnAt8vulhBQRkQgxo
XX/XVpgl9g6Q9Uh/CfoFD+UQLdVpbv8+5aez2YWYWK2IO/hVenNWF55+eDfy+7WXmNy+/wT13QZr
XbB8crEylPIMfap4Aml3245O8gFj24uCDUYdzyt1Zsc87tLR+LSiPdi3dMJKfhBWhasEcwJGkJ6J
dWoN/t6oabIhNQSPyRXspq4RpggkqvmZE92NeFXE1bFZqjaGXZIUdBoPkPg/t55OK5T+cmkoBx9p
jWSP+rW7j2Lfz7znAHtE5tOzL+tPU8+vMOWxqqFOC8RCtqUhLg/uGPnik1KAB0KQu7ulMku5mUJQ
/54VZRLTkYYpfXd8tGDdNfx6JLX224bWRq9n9ST7fSDLTUG1cXhF5bzKHDytU9ciZLrpMxMue/ik
XNKNP6hk3E0M8WntECm1Zqk/rOBhrlrwujcDTG71Ror4J4Jp97scLFFaLkOyoc0YKdCh6dD2q2uR
4POnSrMa7v2ZAQah6HKwA8LAK/1UOSpzlq/DHf40n0hkZ2bqVq4gE/fy77LBy5ngwu47zFlWHk7u
iCcM9c9P9Qek+SR5UZdGAX1eZZFHp1CxzybYuNCWmWoifm39DaaHnzk5BDsNG9izs0Z6AK3Jickp
4kf6zOMmgBauFn4WNdK/ASM47ZgvHaA8ymj2iKnJrKF3Z+fiKUzTzEgffTNmfXveK3COL+4i74gi
cbKDDhYIrKPIbIQlT/k18l+ZdoA5mIJHYUlSU3zEtkjtuizMrl/dyMMx6jeQBGMGp8QMRi4QfPEM
xh27RV9UVs6Blqg9Ugwhlq34LlqjzWS7pRK7Ct+fhjDUmGF+Kqw9irQQaFU/po/lUfMlg5vQizVo
oFzZ0FwDddFwNyTvD8Fm21bGXl6iFtHqf6ePngKiTRdve2N9BvzcAUCbfO0iOp98yWURkC7+NUl0
a5J9JVZLuqwCx8oIWsd542e1CJ3IZsjjeCfBaZa8gs7ZiWkfp6jbnfokwKB/yvbCjnnZ2b3gGwnL
XaOfi/tWBNcZdwIe5YI1fUu1gvTxMHSRoyx5mNmkoII0BJB4YjbbzBZSldhC+GgtOCbINsUUdrGu
g40QQPecAMyQ/qRn8i9pH5KQDslrdDNcZgcKG0wGr5+rHr81BJbmEzy5wSB1GIuiLRIC24U1ZoFx
ftuqE8jA7MjEYNRHVQsdcy1GtPIR7ZoFNFwmdRKgNpQAjAJZ3Zyqd0IOq/Q+6Yx4jAWT/XF/Ndn9
qNQiM6oC+r/ExiMZetl9HDNP2mf1BzXfO7Z6Mu80uYa/7qOe5z993ev37ttNW7GWDX2+ay2Lq7m5
EYRt6/WYi9olO9xrIYxz+O4tkffmdFWjNlDlUqDZ6xZyrcrpSXt33MY3vgwqewBroJ+1iC90KhWa
bfq4wLN6E1vMdDBSXg57NZL0fx2uKrSI6poA+fBksY/5lgWvd33BuygSUzLknRd87ORS+8rKeOJT
ygevFucLl+P0J2NtKgjBziTTQcDRzvAZDqtK712wLLH/syxEeUwR0qi0wxvcYi2vtBF8Pmqo8Hjf
v/u3FAJ7cuaXhQWBcQ1nSMYnf+x83pE7lvf/q5MoeLhmAeLKlX/bKHom/dolVPnTWT2tFyPBduH1
X7rW45MQONazXtXt+nr7/+b5mYbCS66YZ16fzGOc/5wgfoEuNkpTZLZtDgF8RI+IaVkG0vSfwwEO
Uwz//aK1UX/oURBltzsvV7UZUTe5EWa7MRoRBx/EJO95NkhLw5wJe1GiaiRcjHSJUoOepfZifl5Y
+1aLwTJQlrP89EvSDPqA4jS22cH6FJSTNVhIsxHNSh44c+8vo9NYFXN+W12zwkubnUDoqBsIMnWA
toNERGmdoZFF5nBpTHK8z43X73XQk87ssPzd/C8zptQEjEyQro/ddpLi3lAN76IkjG5MOjnnBcPJ
pcJSocCJCAIt21kflMUGRrg5O2K9ghJAc/v75aeD0xdG4aMBiGQmz8XBRsJ0wcRv2Rj8NPJ3KodW
C59voe3aARsjuhaQdgQ60rmsSgPUCgGyyv2JJmiNKT4XdOMCIVuzv53+w01Vp43vlcXVtezxYo/Y
CQW5VL7yjgpjiOEY4U/oVn/ZS+qcwC0vU41Lp813PvN26n15hMzZpVOB0Yy7OtbUyP+zaGGeLINR
esouHMkTLBcYk/L6pjsMXrWp/OXcQD9GRsF7UHkk1geg2ESEZHw6HhZRUU+iQPj1bFwbNdDOB8e2
Ir6hxqOABoZVJPLNqRfdRczBenXnPDh9eiogdOmtNvdgjN1cYjQ/WtuW1X3B0eGaHVGexLAXUskT
LpEITXDwKJV295WWM23Nf0FxxqoFszC20z5t+9puc0FdftScMUd0tySXJe2lHptVyFuUubmYNsWY
Zf4Qa+j2f0p9g3FHUQb9DH0cflLlq0ETDLynRMmQdit8Gfn8DVzzOKci0+JiqgAviCsulXeM56nG
/nNh7WLu9UcBx21txluRrFe5iyCEsW+g6CA2tAAjCr1H2Z99YSH2oESo5jEJhjJy4MFvtV4Vq5iz
+uwl+yqk2DIXSzzDSN/7Vau40wUOWJXsHt1HLzbD3+7BFhHt3VRiNzviPsTqOT+0M5e3mYvZ4VLF
pveDh9pjPl+seyJvZo+++vsdMiX/JSEeana2ahvl3JgI0RtBVTGXFMZgUtvcgBicBtXXb/K2nvNX
R4A8EqmuVRQ2Pnwgl8rdkGue5RrHQTitHX7iUB1jIqiH1JujCJUKh3ktWEQaG9bAGHBXjhq5R46H
f/uK7ItY1yoSH2eX0f57WSw3y4U2yoAn+Ml8KxOVF+2SbOD6umVJCLC/2mfSsjBNTtNWaqlUo88J
OH05Dv9MOArF+4WnFjwrcdnfFu4AAWd3gkwt2CzwX/8OaiutUExKwrD5Y0gq+o8Q/p/Zaa/53dkw
qRfyHJqY6S+ysORkBi0+BP7LHOVrLEnL3GjOxJ6nyITWdxi7VsCHJPOOXNP7/rzrxt8mSI6KkkLe
2+r/G6hcPW0xQfr3Ygf3z0CrqIW5HKRGnh6hdJL6tNqAoh47830hJ3tq4yFfuQLVfEqRtlfeB/Ac
89D5fYk3bmpVPQrjVfMFE6db0AbxYWQruoSZLPYQe+zycoiL2m4rRHMvMgNtr5dxx9WN7TVGq6Ij
8jWu3AivrDengCFLxd80k1qZbxlVaUM/yzY3sE/RjrJOEJBzK0eZNdKKFggVHuWvXq//tYZ7iF92
Lb7CW6ElGXxAX3n0GEo5dvYwyXETqMSkS4gCvGRzrcF87WSOJ+BJlbW9VVJCyItPI5ePl5fJ53vd
PJarpwRwVPLTSQU7qT8jPwYlujNDZ0MXi8syKyZGRSVILJwRDthINP98ck+aNJk5scDmlJ2d2D5+
BQodpO6Hm//IW5titXq0vAbLPdPUSXhMLEQZTCsVtJog2xd3UYcSqZEJUqP0rCPO5rrpIy3tvkN8
p3mDfO2rEnyzicfIj7E3BT2G4TZPtYTIIptGTJ9bk/prx2kKkEeMfUvqBIZR9pcwDeZKbPAKj+Di
kH0G0PJXQ26foVwXsDtqD2lFvdcGbhhmSzvfsSI1vVF9dO7CvgfsZBjRqTUDNvBQoTWuhQjfgrQK
QxiELPtGts/RY45rOMN2gBM4TjJY4mcj/HHfMAk5BPNLeYg1YPvO3Kcs79DHUtXpvf/QKspqVw0L
vaRiM21vx/wTAJxg/n1zgO5/wACMYOJGtWI4cna7+bO89J6VR+0uIRjJ4L3rUVFkEE586D+lrIgW
eXIAG8tLeKPJ6/xs+G14LmK4VFkkSmukvdDzuFRbB/44ktjoipmZY7XJA/ExDNUZnR8pK8k/tgHr
Q8vqbdXwL6dEJNmlq9D5k9pbyGUmg7eLiqJAeelKRrNKiTe9lcMoqSqUCOfm37mPM6eqNiHstBOc
eCc1yjF8OpUaE96thnXAjkUefTqFCM40nEZOZKWjkYlvRFx7reG2nC2qKJCbn834SqgiCzufTZZB
tWKlDY2Xuh/RxTI+r7RyDgsQGk/devcqeclCDiTB2W/p9l+nYbiUkoQ4msnnNXg7XhXurW6gsoE2
bQmb+uWj9zZdIvJMuNgqbM6mvPOPk21YV5ZPeUCBPNtIgtX/CYKJk+d9CQcfU+qO0RoePkspGfB/
tRhOB2tTFIAdYvsYQe1KsPHfCrv6Vf/WUp6kHDz3jJjLs0+F5xz6pFzhY3d5tf3ehEGL1pdPT8qk
RgASczcWqE6COnbnmHdV7loVnrKpakLtTx+SCpfm1Lffn0MfAuBNaKIKmQz73M9wjg3NyB9tH5Pd
Bv8JtHjY227JmrV8qs/uAct5OpV51BZ5k8REco76KggCnywZrJeH1Wb7YW3PM1DPNX2qDlBexDhZ
uTIeJURC55sKJFE9i8Gm0lcZi+zhN84cutqiLrMcDZny5NxYr00jvfJ1/HOSPqAUfwKA68nkcdXI
kQcgwLiscPbwMBCfc7cJhNrjv7vsE1L6ALalvruwg08rqm8xYfvHVpM5YGudG1X5fxZUnQQZBjXc
V1bAF2iSMe461WhczezdElPfEJ+KdlZpK6i9t3/5Z58SFHT+tE4rD3SmgKjnjCh7ary0/d1slUux
GEeLkjw9A0OJKAsRZBgPgTXCnaNzGZVZ8KWolCmcAQwNy5ZE/wxesl2AQDObuv6JlSzHw2BdH2Dh
rmzhQJ4zD9UJrpzqPt4Oy1wvPKyJBpqdasXZ7uwuBs0Lj5vF/aP3rMptVFuaYrgrquvOWsGd75gO
80qI5tgJilvJ9fVjNJrNYiPh4DvoF6jzOjRZSLVjqyMZhieM6my5zReMKcqGS08c+PI9jk9JlyPM
VvW7N8NYTsCpvFsR62kmT8CR9a70UhhMD9w6NeY0ULKEnqa00whScI2Tvl8HovWW9wUdBrVZlB9n
/SzmC4gUdhWhFuab0akh7V55WOPM0RNdIdWEmA2sFNrdm3BjTXlbAeEnxPYjsc4Ab94saFi5e+PU
qQvuzucDeux4jaDJneebe9U7A5ifhke5iiNGKKwAA3V/C+DiQzhvBcp826tTHUAeWpmerwCriYl8
7OxAYrZXdgLcu6SieAyCfANO89hBhheHEPJzwWycT+T3SedMARi5aWfT8EukgMvKOWFtkvDXdq4l
+pw4lDPDm7pBtm12+mWAEo07RBDaAZ6MxJ/ykZe1euIN7SaoVeoTF687iGYY6DrvsWRjZyI0OBJ7
T++uY4zhkskyrpBuBw29K8UhzgFrDWpReO23UEJXZj7bLlpwEo8dBozfKAQom6bFOfcu4ZQshs3J
7TP0itWA6sFKOjdKWbaroS5L2+vzyRAMEspv3+TPOI4Q3dufuni6U7+P30pMTsxU3zD8GjAQv0Ss
l7RKECZGy9Z9tgeqnm50BZflqeJDxHSzt4ICqDrf13fZyWC2AGDiPn898TOWndE58u+Zw6DH4WlM
rDLEi1ddF+wR9oY7J36HVPxEHGykkk2XgS/Hla4uaC1YiUGCZl8PggsnuMxsP2XGI/F0rY3i6c8N
qWztOkSTj7pWXJhH93MfK8BGsH2ZFmW+sMAh3jxk37N+FguIin9BCCvz1GEZt8ciA7X0N1iH4C67
lE0ibUD35MVUfDj75JjOrhPMxoTQKORphC6jBi4qatGN1KRnYnGr9pxDEVAU0p9LXfIRE6qnUM/Q
kGrpDDlBpdnS7omC9Wqh3aIOOOoXv80qJamYGcy4NkKG4Jny9oani+hLjQ5Mh7TpVOJlIuTxybow
EcfTVlGMEem9vUf03+TyVFGh4CiO4Nxc/c9Q+UICWIHCDrbG9RyJT6i9WNfj1icolLSvuEOQ+n9d
rszSTOY1xMX32yc+Z5rXPZSOOMy8agyTbkka9c0cL0aNBD0bOjTiuJbXx4gR5lGCDRCIhfleoSIo
hqcFJBdUQ2Us2KGPEZwLz0apq6X60TBPijb3JXhYoWPD3cUSwmqouaWggI4gg1fGfeE9gqrT/Sgg
EU+6aF4ccjM0FtytAphjzTK1Ud2UezjoTqO0Gzl6o4JZecfN/UtQeXwha+AcwfwGdK1sknumNCQ9
LLyiZ5H66kgKfEOa6UNvYnIWTOcurww+CExwIX0lzCudzEZWVAYzfjLucIzw5mQu1SK1CEISrkwA
l07Nhi+UmwkP+sy+xDCZF+4pPL67SZIofxEA5Ro9P+xVWI13DfVMYM4qC+RmqMh4Ym/OxE8j/55B
rm2ftKxqRDvhG7YQjIQU1S+g2ZuMBA2eD8ajBhMEBPsBgOKRlAWS6CP8URq5JCgtriVLt52ipApj
7Mc8rx2KGtqDU3qERvP5jRFjg3Wi4ipqA6A8MM3ERmNYpDRe2u1dUM3EpQRdN0N2/78YSIjBwHES
HsKCc/lUXvISI9u+mEbpb7gCaGugsv9x46J1S+VL2Ftt8g5LHUt5ynZUFvShbRPqGv3EiC07C+gN
RXj49vCsqaOMweF5/x6n5h8BSY8bMXgnkCAlglmc0dWLdy7C29xFEO1UhOd26r1oK8oSX/XlbDZx
LUHaPyu9gSUrc0dJI6rqaldk9/egkRXJqNuxs5LMkaFJcAxeUxpl6M5ssLd6VFylhPDlSajullQR
aGWYNnq/tTi9UplvQGNBZ8/qPErbFOnNSic0OD7LCc2FujMx2FgIlLZaFCOIRTgWuFKOMotY1Ddw
NXXO4Y+Wqvq4mhtwqOi61FVS9r8hD+9DE8tK4ysdl+rDdZ92jnjoC5Kl+27RfWwx+WYZGblfMvAt
Vdkvp6T0hwBlZ55CkXEGwEjtjYYfUGl6y6AJiE1deeezHG3mD8XwcqfukMMgvm/yMc+nwYdx0Id1
J8V65w1GVAv/ixI3oDHTC+gHYtnwuwuHXamV5F0hrfKd8BoSEy0Z5DqsK6iv/E6l8a+qiRs86Ypq
soTRqdrsPTNeDDLM6lT/DFw9XOVdbjFGqXHSAUjbzGU6ZpQJXhO0mzR1W2v1NkyidbaQsVRK3Qph
dIjLmh5dIFgQa0sICd4LxgL86AhtXTPVPAnONBCRf/lGCMImtyvZWRyR9gelOGusnev2BL9rCDdX
1bGIzS7K58cdDyl734dxoQPCcs6RwfLTwoHJFl0fHH3BIaHS1bqYEpFk2yGljFL4Af/o/UOWviLo
aitknySZj7LtVyLZzxExFSXUid3DLc6EmOrdr1TSdP85h9T+0lwPDw0G8CzjArQYRoKK//wGgdRA
maSZcnV3lHZkI//fguepqqEShfwWZ8wuoKdp5/fNV94WwLIe7epKJimiFIXR3/U2GiWtKuqn/2Px
ATCa2ibZoxqmcJb8r4aZBodd8iiS2MwJBCWI9Z0b/W6pV/Rnq+MiIhqhlxyYnhz6yjeS5iTx8Chb
ZJf2NC76UGggwFME5l/zGS7rjCXLikPYNTohJmn9C8xKglviSiOIGtDijtbIEFAsOuabUq7nI3OP
iiYK3Bz+VxOLvVEhZ6KmXRSqBrYS6wksny5BW9ps9XGZDyZ8SUj7DdYUrFyp1Il/QvlaiqlOS9AQ
r0DFsan2ip9jwcT4KWnrTdAnmafsRbF6EE8CY4OBf0IBzMVvFPd+7iRPkmMvxtd2RG1+HlNIEw2t
BjW8h0rAJB+vPixyzBW4pEgO5W2HUbCXKWDTZYN78ziKt9QOV0cPg30Pr649kn3/7MJxva/utqMg
jQsqZjc36RM4ScjmuviwvNU3A8LvKnuJL1032FZNH2oKAt4itBniFq9hElWKaR2y3AkejcbBkz3h
1En9/pn/6kXuEYBbFYCRRjixMqLeYqcf15MnsfvCcuXfjwDkTpC/6SUej4nSVTJ/7yVWsT2R3NuP
OVFNnoGmUxUUMxgbWQt8YMmcJnyAD1bbP04IPPghj8S9H35FYdzxWjDD23FACXAubA5D7HpE4O+R
WntasIaWUaQB1taY4jUSK/tXfDE2B5wFfMXi7b4QJ257lb6T4DZbeAHjx0+04EhNuow7PO5Xis53
P92Oh1XHH5M3u74GJjQwGVNKqDY562QSSWo9J0VogZ9a6uWBCVNUgPJH3a6OOnHis1QsejxB8Ok3
kZ/IdHhUjWkhrpcHKJpYdbGg9HUOb9qH2V2OACzYSDwPxy7m89YuB9qtXkxWhgToUVXoz4rLeOAr
j9IhLnYF6YmI8uq92+ZObzO6MYGtz+W/Ya0YCQmIUsIxepdzP6odnEflK30CR95VS+5TSDIFg+Tp
Vu1Orc/0BlCuusajd9QvWdft4A5nRcdRo+f/vBsk73H2nSGWP7SpGcgWnomINHgsMFduQGXaj97d
Ep4nPkhGaYb9vBYk//CYwcO4T0jdtjjegw7AEEUuFoChE7RPE7ZE1xevHeF0QmiqYXX0PHr9LpoP
h0TuqbCJg8NRsNxcOXnnhswkxmBDaLZwLeQ1xEc2Oj7dBflV9vlS4dKknN2XXeCWWOp+R+Nd3R9o
28/nXfrofbyziHWpJ6GXi8on5Mqml4rgWxRQmvrivat1ElTFEaIgLFQOp/9tPyt7Pi24EdcW6Nuq
KknqhIqrBRa1NOa3NfRE3LK8kGJDHeTMuqB6MGF3+Yby7q968Su6To545lcM4ot1+HeJ8vRw4zI4
ihoIt65AYFkSRkmqfmRT9pA1MU9jqw1Bsz8+iDs8kXQikA/OdkxdxQSuRvLWLM/CVqW5qMQScQDt
Lcq6q1AuyyVT/VFTCs+ddp0cad6wEifcImgh0Wl2akAB+xiXI5Pdc8RSKfdMuqgGCzPKCiX7nuxb
aqL5VFML9Iajqhq3E/GxtdHqURzukg6lfjHHEmFykyWWTEhmlk0wJHuTB8hO7Ey9Y0LnooODjFIh
kj9dXz78ayNlG3qWnxg9aIe6LQX8Nf+TdqDj7ijPFUddqOGrIX2bgJXulyRL/xQoVHONXCuKBrS8
UrFpNv5UgBLp730Is6ehQhZgpNOzt3tzeEae+cN3shslrKIvr3ZxrcoZs6mjZamIgAo/NhB+5u2v
UEE11mhCrCFr8vixva9HRoL+ACdnDYv5fwQQ24zsd14ueUrjCZYNZibTcC6ugsJHj1ISC+HXqbTy
CQlrj+N3yB4JrkgZdDCwPEP1wU6qReOTp45+sgxhFOQbWzE2mG0b4X1jWofxvglI2L3H8sG8ebQU
sH0bKFoT4iNGp+M5JLFLJe0Wmqyo85a/2tUiMWD0gcZ4/bGAOXu7YCrRz+cWm4V/mpNRrtGjhunl
fXoy49jrpYdF2mAPaWp3HzSxncNWvGbYW2Igbb1dTmiCiuxHXVlwZxzWPrURlVZa2hHlq5ss5SKe
4OVNb4uQl6UZ7MP5fo/KjwrV+SlV4kuWbXbWPpZZ9fvl2rdB4lJ48XBBFfEZjF0UyRjgnvXsCZwF
lSaNhFBRmsM4lWSVFynbJNKp7eUowgBO05wqs3QRfLltJXbtpuJB8Uore7YUtFrNMtHXzcGhH/Z4
O3stea7YVGAehiDmHykLQD2pjwTAF7q3dV4GtCmJ3ux5O6LOSU79x2pTnbvJJc9ZGpuWcrKPAche
JFPJHDE+dG31VwCLYPOtT4lGGUEppwBrE0wNQosTWkvAzthdrxoF0LR2vyvAPwMYoaSqp2z29VaI
CjVe60ETUc1cQ/rwNw4PWOVYAuHkn6c0rFizcnJWWZb5FG31rqJSqfkClDLL1LhmjrasdTu7niLA
djID9DzX3PJe2e1QKZm57pFLws2q7kKXr6t35XrBC8tzmudsewboQazCfYeDNifOgkg2V/2phiIT
MRr8FshOBVCCrReMulQKi6vV6eZiQsl1bMO3lixK5kaYckRuPgMEmtwbXi7FRdbZTHaVqBZANAwA
eNR/0LC5QjvIfS1LRskYQfXjnUKQikyygPRCsBJ+fAKB2bqSMEynqC5PlEpXQBSNl4bZV0Q0F4IB
p5etA5fXEv+OdQdEP9oChx5TNZ9kBBGpoTevlXv3L6vkv18+xGbNxNEgWrpEgT/dvEE/edgnUaNt
3Y5+k+lZ2zSP+nO0t4S+xloiQaBdqJI0IW29yCTzUYWBMHDilqx+qWWUL4n65DLtAo+hr7Knuu2O
/lQk1aqAWhNTkZd1buJzmHBxUBaoLFBjoWj7nQTshtGyKVvOTfsvASnkl6z1v41ufyXi7xvNC1+4
pqDYX3UenFXMHXvNNDmv9sqFVq1qqAzUEUxxxU4l7oIuSM69NIhK3WDrz/m0P82Msw3asL5QNKIx
dTQxlJKLpk2Gkd01iQf3IDjj07BwON/aXBk279ljnQXWXHBVdNHQy0TOFj91QJgsUaWeA/TV5I/a
ACmdmx+PiycePKSmdn0rlGsDzvZVcY0CasfnSoUoY/xOQfskJFiJp2GU/HNgP3gw17+ItXaDhNCe
5gefZS+PRl5XXnk8RcYlH/2i17peT7fcnsLukHneQn+p6SOAi5EgcFM2x9jWUt7Vk2FGjNWtHJUY
29TIIcyKeWuSQNZu0YROVq4Uj+GTNDlcdwZMz4AuNrZdOF5QHP8j3SpvByHCVyGCx5QR/7C7SosC
ZFks1KOqDgIaTgRQd+5+C2hyV+P4zYRMaiMHqphyXJHnJ+JafKovjXkPs7IeK1ttyDhNfziDTLUP
7azXbuELE24TW3Xfd0G/YretpGAtRPOMgo3TZcWbAaUUObufv3Oomuvfwi0rzbOQuvjgBaRbSpwn
qS0HoLfQ8l/4i96zPmnV0JX/ctm+rZ4rZLEEjBJGac/lzOsngpiynDeHICPPqU/2lVfDl9oB2C8E
TPHAsgL6OECZ7ngKhkmLraAWLbs2Xuxky5Jac8w0mdNyjmSVi1/6l7HQkzSHgzc6HoAieu2bauNE
NYh/pOBejrjMxQeh8023SmaYk7QGujX/Nv+JggCuV4ylcIOHK3sM7bUkcb9uPZGekXx5g/QH5If6
xzCgjBkbCAq2fHtFB56nI4mavUrVxXJPuQ6w8Sr00qNtVDlzpuinUmGRczolxFfTSYn8XGuZHGgo
GZseFFlbR3zgufPL6KKE+l8GxGP9dhEmIPEyzdmxwuar0Ci/VkhMmSzPFNmW0UU/6ZKNbEYWyJHL
+Kv0E0Pzp9NFthu5AHl2EYM/GcVmjnWitqP1qGRayKLAEMd/U6v6POnvXtUunBo4YPepgqyqb/0s
uNLcos9kXJWkZgVckFj0Ue1KPMBO/yg4FTfwLf5xFkWSoPmXMlahY+pi2jPy3Synzv+JqIJ/OZPE
BZWk3Vali3WvwouGv+zAMSAi3ELrAbkC0D3Gb4CXOn5oxewYZC8nfZuVWGy3cbVEA55h2mPnDCIT
UjjfiXhtrsXtHckvfIZPL7OpL0Es8hit/LnwSRAEowXITS7NBJejta9tRHgxa/4rTf9x3Pt7cFDx
uyP67Ut1uP5A69JW6FcdzxYEwUB77xHyKFxzi388LQyBoTh+bTPfu/eDVDCS6PnhWTjI5RDB17Rz
XdG3cSdnw69S2tXk39HT8nylDpuMhyeTqraQVLq6N8zvBPryLrsvtsEsEZb5wsQnHTNd0o98AKWD
ncR62JQLDGr9AG89E76tiiLUwC0AwO5yFHwtgyr8HCisKrhWDTR8q7nm9HWtTCY098liMpPoGQWT
A42uBcRfyKs5wwQNWGhOgOYngfKWMR6KRf1YBMFOCfb2/fquWLQQ9AEl+3os3ao3vlQeiwGZVLcu
1GD8JRoTTxgcy+zoaJGmst4QM58Hnkwy8PF7mE63rf4IycVD2z6d+gWBjJqSO9T8dWh0bAF+M4O4
Bml06sbzvf6YT/5W+praxRlGpesDNEYXtL5atZ44z/WZG8JfQN5u5alCa3psyv47os15VagQkZSn
WQD9WpLmNJS8u4fFSwUWNcq7kOevOV+EfI7/f9m/dMKDQnuC/jxLdfoHz9o7mJkDv7z17fRn335E
bYURJnpbangehWRalN42CKmUooktfE/YJvSvlM3Y4EpOwuKX1rhLG194BRpSMcwhE0y0i2N4ifVW
cVu0hpms92pnX49eg40fCWhArvViw+OxpBSVkAqfvMODUqzif1JdnGiS2dV/IbFGDlOX5iTksQCK
qol0pJZCu5v9JJn4Ecu+5a3WuxJ/2R9CTMgEX12V7rcbuIfcumXrBCyzoeI5n8rFqmG4CIzhvX+H
p7Y4OMUgEp+28Ux/jt4jlipddcfBR5v4ovYV/bbhxTx0SyUz4IGC7tURnJ6MsrU8T0qxvy0wYq3D
NoDEenaRup1Z3fF/rb43HecphU3tMp5+HfpsGzyYWG95P9J/29Aoq38Foqq9CIPGkvDWpBTSRXZk
DnFgBkFUNBuKp3UBpFk6UH8mf5sFgmJait4O6CX+bYImnyTiYtcuVAedgO56kSZMHmKcWuxhhPMN
Dt95h8N3j3ZvY1fg/pocpBCVMa/QZzAXIlVqbc4v7fjrlWo/CKLbaCvGbXY+L1qupP9dE3Wc/QXw
HITHMavMTZFhIWIDE5rTam55m1c3vLmrpD4f7ov9d6huFtSaB8uq/iVgbslvY88Ca/nxDrxoTMfZ
GaFL/98YCOKS7/s1I1Ikt5y7fJ3iO5YIi+mtMiijeX2g2zEo0gNG6UPY1/fmmb8nRUEdixrbVAwR
qsqFpy9WBiewGX5ZQ1uFx98AmcYmqToyOM/TXrlLtKI1JNIQk97nWX2Vwtxu8QXGsQvdU8tqV+V3
yZKRheA9qH6nvHHyO5yBsvj9QIsbbW3rUlMhLOsYpfJX/XgLmfwR6yaN6B+4vb62YY/IvS/4Pb/h
p207MFwNnUBy5loytVSghkoh0mw53IojR59D+1cLRAqdAB3Tq0ozXzzS/aJYawHuZRXRrOKKvpoy
E5FAFoO1ppGAT4qkRguICf0vFwyCc7ExTEsHkag0UR7wW6wggjGEHanCrJgZ/3NTQJGDKZU35kzd
FCO3DE7kXMJuxZzpbE0pezj8v89A/xiGPE2/nTaYptC1oSHSRdYORDF5CM1U42IHRPZvqhIDfoFV
jM8w2JRNi+TjsJJXxE2pUhmm334eqWMVh3LwYwni6GaKVXwHGVJCPHUwDSM7iMyV4NJe/1EAsMg3
ZCl/z3CZe7NBDLddFx69zHyzQ7LOr8Jxcw5+sbnHArg/hAZJ4ADQqeGfGZNN/0igJK3O3jPG9lbn
VEpqvPDjPXXJCgo6bkiEqJefPzIdDSXJbSBT+cVZ7kr3fSe9S03NplkBCMbhFKIUctwClgebsBsm
IMKjRbTHkjbPms9doUfG2XmgY9fY10oDi49a38xY1YLxnKRxK9uhoTcyYTUh2wqqkpXw5Sl0Ca97
VlCsT+57OhW3B+AuAIziLXxJ0lhC8UOx4/5IrDDWDFIz3jSPdLrCTDKnUkrYrBRgLR5mhQl1Gttv
eUnxgECqjTdVZYfu1XJ145G3wf4Y/UGDJ55dCUpUrBltN+dhQ1I1SaIAtEO2c8OVTpp+I0gnzOMX
eg7q/8S8X/HZFv09PD5x2AxBNqdUMsnj9ReQJfneBSqH8L2KgnLl0YOIr8jWJBF4BL7fr1eDtAEz
5/lSGoq33YxxpPd33k6UJpTgfavmTd/holVnz/2XosEbU5YgmNcm+z5u8OHl+Yffv+rRnLElxJ9m
HbbFKg4KIyorwLe5Wc/jHrUwBxtUEt90NjwelONU8vHnqAHmNoF4hAlA6LuWAvieSjqq30Bw3PqT
q2EcyilBqPrtc/0nhYWaQF1Lr48K/ouoRpPFKHuKlU412CyQ/2UEYouvjxAB4fyqMSloR4aa2vHi
n8dZtc0hZVVqx0phI5/YDxET3T1GyIMb6n82zS/QXjxMxyjEND5L5rHlI4fhnMXyG/+aoTVMw1+P
iQ/x9Fw+4RNIosHz7SJTGGqL9gWDgWH87ZM5QA/rD97vUMMZeadwEOtowEBJ6QLZ/KwBnbzSBpAv
5IeybrgWLJCqhJe8xtuR0DPnrQ+6WjyBsLOvqngRaLdiWpMtZnS/c64ghUFFJGelAITdymP6WjMH
bV7z6X7fY9SEquxSUtsj95xSdEPYSHavYIrSnLmvqcc8nn/vOl8NpWeLpc3M0UxDeTc4oYR1ZCJh
Vct7q+FpGA5nQmLFl1jGdn4WSNEFimweZhIbByLMEt3Cqk15QhztxncszvgaRay0f2FXopp2ahgc
MPc+2p3I/adsfw04YNXo9pn4A/oK0LJHgxBLH08XGeBVmjT4/GRC5dwMpOY/VLqprssShkXPIvU2
ic/8/pSXJP9+dVPToDLK1SWweLkFsB6GybG93NRUltjbV1S9UfoQZJMdzSog0JRAkWagDKOsKWPB
hB3kyA2lC7NqAp00mWq1QaHEVNXl2kNEN/hIv0Qz76rXZGcqz0vDtJMW86j02P219Sscboq3fB5J
msfs8rUAXXevm2peMhAGipbo0GztDJ3ylZ1S+pDHc772oi5Uiz18Rrc3kyH0j51vd6aV9mKq6OSA
BsfqfmJq/dz6c53P5cen3P3veh9dtcM3x9Lk8z0AACLQ7qonqJnzejD+fSY/EEHPzPfytgrVzslT
IE3B62RYRDnLt3HGT3/S0h8UXZNT0/DuWSFwZ6j/njiIwkXjmREdxLPUnLk5Q02T4RmBwmjkVXhg
wtal4UNgY2Ulbq1d/rr3c3qB2EIJy1/oHCMcsT+Jg8iTpKdPjmWZXI89A94lpLZrxLNx6Y2vdLZU
OCUKgMLoCORBc/TtcXllpnVlqvqIr5/ikaEHsFN9jeEz8MqKgpM6PFYMzI4Yl/dZGBVT1S8GcuLW
jyn01cblCWzY2F1tur3kHDegOWPR0kxxlkr7YTcY0ZZzaHIGXz79jMcXbql8LSCYXuhMI23eokJJ
raxMDLx0Z34fPinslGSve5H8DSoP+lAvIhDQyEhusXslzI67dT1rNjRrFpfd2menk2UapJyzhMAX
OMo8RveKM+rs4/nt64aILIDPIgEEm2Ae6otQO9zKtHQ3cLI6439KBjU1WDUnsP68H0vHZigaiLBi
XdhtZtmPZmmbRG0BpVpOoxmwQ1Fh+UQUpibuZuhS/KiONUJGx1EVWuJYp3rntLaLrRHEhJH+oLd9
ZmCItXYCBVz2eFMA7Mouwo3v0ld7H3KR+faVl3vktl1/PcktGZiBFGahCom1aui/9W1zKUP8UIkO
hVetOHbPzC1WVhG1Ho9CVGO05dgdxXAunQIqCwzAee205mDOOuFnLJH3IV+EEK4QPIrEtNv1ESgW
SOTHTKgukHQq+1AOGBFj5mN+ZR5V1T76IVRcCmvKO0hvyTpeOC2gU+Y4oRdLQ/uaN8tLDQeZkXBJ
CO5uY4Vj+yZrpc4nWbUrmMkMkLLusAM7e/DCFKYXjmNDu2eR+LHy5lxzKAGJMUtUyMeAEefab98Q
Ztm5IiOg9HQAj9yZqo4Bta8bAY0pFWqqgjAYlSeBG6xsvjdobkTZm/p5PZ8R8KO+IhlHqVHDdaC/
DG9SsQQpp/wgqSAqJlaN6QTSrADOmFzhnqSkyiuGCa1CB1mMytJ0PMJ946WVuX/5wzjAL6/FhhWR
WVzpdKVUlId9Hu5E8BKMG2KXX1S8VUfRhdYL7VPfBfFZmB4Ck1Xm54WLl99HSWEQjNt3cv1oe5j7
TSvfN7V4aabDCka3D0h9RQ8LsTPyjKgC2nMnljbpNAWren/JZfn2RUXOuW/XDx17UqwlPdnpHZXs
gdrOBQWQ2NriADyvEdDK2pYOQwebvasxdcyyt6sf+z4nFAFHhq7V/vlpc88C4L7FjSbdWmxecCyD
IXQr5alC7BEvuw/rIiSRFPWqoX2pO9XqOdkyItezosTb64u9+HgaX5vtFDPWubfz4AhM7Itg5+WZ
by3H5SwJP6L4DQax/Lpbha1jsh+C3YgfiHH19KcVEs2vKNUEB2tIO9MmGZYu0nzrKrNBn07jjcuh
3Xsp5cIpJ3RsV1M0sn/lBEHbCZ/S1gX8faq6RP1pPvg3pMPlJA9gyP/uUByOde0v2fiWKNfdIli5
AE9NINzVYexjPVxyp7eKPbRmtYjCrIyCvK0kQwJtM+qHcDbk+XpAIXRmIa1u3eUx2kejLF5Ce0wU
3W5XQF3AHLHCkuntDwuvYPa5K4RRD+AQzPn6Sr0Hpa/IDErimPwJ0JAtLof74xIqq3ynDCHEB8Jz
jPissabw1LPbRYBlEou+lQh96Ge0p0fbJZ/DSDINFJrzxX4axkzhoSdrDVqmkQY4jB1GOLjkYCcT
UPQ4yZkD4LGUq7Z4kbgju824TU2c/9T0zAEOKxZHE97DtjYjUAuVsR41ajUHEz6/FTROVIHUS4NK
6Pzk4cl7E955/qaLHlqPnYCDVB/QwGVmtruewaKx2t5+lN2ULBXXRr3wjIKbZxa8m9p4pvY6vCFO
gBKJCUiV9pFzdYQTsefF3h/1npvJplpq0rSXajuZeQJdk4Gk36tlhRJ3rJCuZ++JIKSZWncOZMMU
M6Vpg0T8bRZ0fBDV0X7+pGY4oUn6qt4F9+d9srvXL4GsGWq/Uj4RQF7OixwWaqba7Y8DTVOK2ge5
ibZzAZHIs5pNGZhkjV2f+YTYvbk1aJFTfP5PvHPvD5OUV9wddFUPNUQtVdsf4SoBxBkSp8C07R3t
2rFHoRnek7SOrFFfj7/LVqKE+gmIA4KkjxnvWOv7e53Kk1xof4qglGniL8sUtmrHNPVEI2Mf2pqS
/8LijuD+QJqsVAa/m6opLt/37NCm0eWTmTDGZ6qaSMcerzPMuAbUq7TjUtZU6l5SsZ1Ca4IJPAv3
4IRWTNSal8WtreXLijrYNW4TOhLHNhb0EWKEU5Ljk6AFQJk+wuGxNbMp/EX7O3inJuWVyygX9UPB
P1QeC7GqEi5CObYdms3eu/C1tVOWvpc5sO2F4d+LygPHdz7ZJVMQroYHwrkvTawdPgtRDrAhC70c
0DMXtpE7rN4DQPv/BVC2tafzMDrmp82/FsadOsRoQ7AsE5KHEZFEn0pBTBF956RFT71zESIeJe/f
pubgmn3SwCOrelMjew7UzCaR/V16y1f0MqhtpBrX/4EeWkvXAxd1rULd01r02Ge7doZ/RjdFktuS
K7LeXyxuZ502QwEtElqO0l2/OeemH5EKm6TqVs3u9jAJ+Ui4tsmwpl4RKPLXP/BFvkmfgQI+wINL
An2JFUU54OE6xjlgzsn6abXg++IhJtv1n07Ke0oVVEGb3gyTp9xztn9CYk9cNAvKhpQvY7AOXWUT
Ez4zfAUpRmMQshwp+hz8icqIs7x24EhDs431Rn1R24b+F2jyy1DQ+xce3OccxBw/o+/8s/IOeLja
RI3P4qYz0AYKbSa1rjyN/InpjglaqNJEw6qPNxUtDJh+8upruM2wCxylwI00XZuY1VZQKdA2NnUb
Uzwee31+El1iNxLKhuzz3xrPapWrll5JQMwI0quLXKxsaTFdFMCghplU/4Gc2cbMO82vF+2k89Di
ydfKADUwx+fgnwc7enbCI2OCG/ZD5nr/fr0lHlV+ShnfcIyKkSdQPjzK8SqL9+2HxEiJPlDXQpOO
r/YHkfMXxL5cL0gN0Ce/+goVUAqH4qvNZTpdP4g79Rrs/KQ/56rI9QVH6tg01rBWKaLI5Z3+RLpZ
95MRxuBPePrOzz34dzQ9UE7WuWs1uVa3VbKYu7spG2r5wWBmMsM86J/afcShLmQPH6VS7QrkfK0m
eT4e0scMlIvSGDKwzOCeSE/Ps7OsnclyiLnuYvKFhSDo+UgbyNOa8M3nVx8w/lqpvl6NWrgjZ2gf
yDYgoZ54aERKyI2YvIQQodsBYp1JqKsfSGHGkQqLoq4jJg7Y1hux7qJIkxUAHC6wkVrwLB+Mgulb
Tlbsza90MZRA4Df7N9LcEfmwZ+2DZZFAnN9URImzuoJsUorjo88/Yb7CHQ4YTXW05xvVhSIut7OU
xrE4yF7c8776WGp6KQ442ke8A+uw3eqsSEqelWUbbEXHqHPzuyh2ZnRzOfqO0KNSapxBaGv6Qo3p
KyYpUZ9Ey4oU/9TPLlu32FhGeJWJ9oIycalf7+86Hh9xIzjCYJ5MEB7VszgG7sUMi2a/4D/uMMQg
o5q5fstDXJulSIq5m/7uLYDtDISbpHw9VzF1d5JCGkpky+OR1KPuyhSEcTABi/YdhmfSa5giLbIS
RsZQLfBpjT6YylaIRjVvcR2d7wWotU0F9F7D8c/tAmsjGHmtkgu0rKOSGPHxGqKL2OhGYR2/daZe
p0YldMKHqsotwdifAwpv4vddVAtEvRzyYj6j4K4SNUhnpeNtEuFnmEykZMSqfqkUG7Omo5mH3zrr
WbqvbScxSDN1YWWfgcrvnbCJMxPJBGGsH16pYt2FqmjmfwAw/DZqCvzUL0JY9h/N0gfm8IGSlRu4
qEjYuyfuKgxAWrht7m5XMcAOYYbJRq/aZNY5NP93A1+L8EX/BZvE/4biwHya7kJ8ElpGAsP539ex
M6oiALzDeQpDMVkhTxtxrkA2H7vHtGkIiZNIkssp6J7RaEQf8pvAP3VmfEQCbLUX6ML/ZdShNLBz
2lBzIkAWB0jqt+G7vaGEI0GCbhBGDxMDaNIaFQFVuEQKBP8fFqRYSQEUAqF+4GbcMZv0j8wgzGuK
AYycDoAlU4xUIK9uEsLw4dpdx4yBW67BKrTWF/k60QaRupyKgM+26f6PeYdXtoOFWEaKTD3Le+EI
RczwTfCF//de3hJN41i27+i2m9ggzIulY3ZMIvpRMH0cHICGbXj9fE+FBFP+5ZdtdDXkZf/a6Zgl
u0ZvDZ495GxsBXbCd2sTGshaK5X+tmBrWe2xrNwGIfRkTzQ45mErITXiXLshC2aDWCiGyBnTRwix
UaKZykCjch9tBIuTsop1bx9APU9Rsd5DYFxnxu2s6LKpC1Kr+B4=
`protect end_protected
