../../../../../VHDL_Files/V3/regFile.vhd