../../../../../VHDL_Files/V3/DSP48E1.vhd