../../../../../RTL/FGPU.vhd