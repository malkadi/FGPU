../../../../../VHDL_Files/V3/lmem.vhd