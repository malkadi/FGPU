../../../../../RTL/gmem_atomics.vhd