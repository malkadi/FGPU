../../../../../VHDL_Files/V3/CV.vhd